module fake_netlist_6_1030_n_5453 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5453);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5453;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_3294;
wire n_2457;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_3517;
wire n_4045;
wire n_3893;
wire n_4598;
wire n_2945;
wire n_3061;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_740;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_5382;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_880;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_3141;
wire n_2755;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3501;
wire n_3475;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5387;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5425;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_3114;
wire n_2741;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_5369;
wire n_975;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4336;
wire n_4201;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_L g710 ( 
.A(n_388),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_150),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_202),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_35),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_242),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_160),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_261),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_685),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_47),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_136),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_259),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_348),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_627),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_667),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_506),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_520),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_351),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_487),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_27),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_280),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_429),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_557),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_258),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_529),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_182),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_695),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_138),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_301),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_708),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_137),
.Y(n_739)
);

CKINVDCx14_ASAP7_75t_R g740 ( 
.A(n_523),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_509),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_512),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_272),
.Y(n_743)
);

CKINVDCx14_ASAP7_75t_R g744 ( 
.A(n_291),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_381),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_296),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_385),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_664),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_223),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_669),
.Y(n_750)
);

INVxp33_ASAP7_75t_L g751 ( 
.A(n_500),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_682),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_292),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_678),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_633),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_644),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_497),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_603),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_506),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_91),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_331),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_518),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_503),
.Y(n_763)
);

CKINVDCx14_ASAP7_75t_R g764 ( 
.A(n_293),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_207),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_444),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_601),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_35),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_228),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_48),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_412),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_84),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_135),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_297),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_327),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_461),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_684),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_447),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_407),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_213),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_61),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_280),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_481),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_369),
.Y(n_784)
);

BUFx8_ASAP7_75t_SL g785 ( 
.A(n_48),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_441),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_394),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_184),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_233),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_534),
.Y(n_790)
);

CKINVDCx16_ASAP7_75t_R g791 ( 
.A(n_485),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_165),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_498),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_437),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_458),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_235),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_459),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_207),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_536),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_12),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_444),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_625),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_97),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_456),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_481),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_555),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_574),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_86),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_375),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_687),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_580),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_504),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_165),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_345),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_37),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_336),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_221),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_320),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_337),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_251),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_701),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_613),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_602),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_434),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_468),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_683),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_597),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_512),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_509),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_361),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_462),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_416),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_263),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_29),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_251),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_49),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_247),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_628),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_706),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_471),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_0),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_482),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_268),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_508),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_708),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_676),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_600),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_217),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_126),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_604),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_692),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_668),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_441),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_237),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_379),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_220),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_174),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_320),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_286),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_140),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_44),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_427),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_448),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_153),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_637),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_464),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_34),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_599),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_27),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_704),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_574),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_651),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_648),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_695),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_232),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_5),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_643),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_501),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_583),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_302),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_573),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_524),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_653),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_673),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_315),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_393),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_13),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_663),
.Y(n_888)
);

CKINVDCx14_ASAP7_75t_R g889 ( 
.A(n_215),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_461),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_371),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_681),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_426),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_543),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_282),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_214),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_75),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_425),
.Y(n_898)
);

BUFx10_ASAP7_75t_L g899 ( 
.A(n_107),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_492),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_206),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_105),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_570),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_145),
.Y(n_904)
);

CKINVDCx14_ASAP7_75t_R g905 ( 
.A(n_351),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_191),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_87),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_566),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_518),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_391),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_131),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_419),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_73),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_285),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_585),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_405),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_469),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_496),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_279),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_689),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_225),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_65),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_330),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_702),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_478),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_566),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_681),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_300),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_301),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_390),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_411),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_354),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_564),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_85),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_330),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_89),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_84),
.Y(n_937)
);

CKINVDCx14_ASAP7_75t_R g938 ( 
.A(n_175),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_287),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_69),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_29),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_108),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_644),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_166),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_28),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_367),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_691),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_121),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_261),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_448),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_15),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_122),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_237),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_357),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_437),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_358),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_39),
.Y(n_957)
);

BUFx10_ASAP7_75t_L g958 ( 
.A(n_134),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_637),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_93),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_543),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_534),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_365),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_95),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_105),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_88),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_396),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_640),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_153),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_510),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_667),
.Y(n_971)
);

CKINVDCx16_ASAP7_75t_R g972 ( 
.A(n_148),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_656),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_596),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_686),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_22),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_215),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_660),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_4),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_539),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_129),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_70),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_598),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_195),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_562),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_588),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_672),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_453),
.Y(n_988)
);

BUFx5_ASAP7_75t_L g989 ( 
.A(n_674),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_240),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_294),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_242),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_187),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_289),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_459),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_495),
.Y(n_996)
);

BUFx10_ASAP7_75t_L g997 ( 
.A(n_412),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_198),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_309),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_21),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_358),
.Y(n_1001)
);

BUFx10_ASAP7_75t_L g1002 ( 
.A(n_577),
.Y(n_1002)
);

BUFx5_ASAP7_75t_L g1003 ( 
.A(n_396),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_256),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_617),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_104),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_19),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_389),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_418),
.Y(n_1009)
);

CKINVDCx12_ASAP7_75t_R g1010 ( 
.A(n_84),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_184),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_547),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_435),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_648),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_552),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_633),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_420),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_411),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_130),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_263),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_19),
.Y(n_1021)
);

BUFx5_ASAP7_75t_L g1022 ( 
.A(n_100),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_6),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_668),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_106),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_523),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_345),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_189),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_705),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_522),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_86),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_199),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_281),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_90),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_228),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_572),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_319),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_488),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_229),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_346),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_551),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_599),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_308),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_689),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_540),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1022),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_1022),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_785),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1022),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_740),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_744),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1022),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1022),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_754),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1022),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_764),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1022),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_889),
.Y(n_1058)
);

XNOR2xp5_ASAP7_75t_L g1059 ( 
.A(n_781),
.B(n_0),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_794),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_849),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_905),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_938),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1022),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_791),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_989),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_989),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_989),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_989),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_738),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_718),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_989),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_794),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_989),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_989),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_989),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1003),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_1003),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_1003),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_875),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1003),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_972),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_775),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_747),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_1034),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1003),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1003),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_718),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_776),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_777),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_881),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1003),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1003),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_719),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_739),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_800),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_834),
.Y(n_1097)
);

CKINVDCx14_ASAP7_75t_R g1098 ( 
.A(n_899),
.Y(n_1098)
);

CKINVDCx14_ASAP7_75t_R g1099 ( 
.A(n_899),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_782),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_794),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_899),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_836),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_794),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_771),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_817),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_869),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_732),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_794),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_787),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_788),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_898),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_902),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_922),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_898),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_937),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_945),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_789),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_732),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_952),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_964),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_965),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_898),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_966),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1019),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_792),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1025),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_761),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_761),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_898),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_864),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_801),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_801),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_793),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_986),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_986),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_1018),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_898),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_797),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_904),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_904),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_798),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_904),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_904),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_799),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_904),
.Y(n_1146)
);

CKINVDCx16_ASAP7_75t_R g1147 ( 
.A(n_958),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_804),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_772),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_914),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_773),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_914),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_803),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1010),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_914),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_914),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_914),
.Y(n_1157)
);

CKINVDCx14_ASAP7_75t_R g1158 ( 
.A(n_958),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_974),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_974),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_808),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_974),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_974),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_774),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_974),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_805),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1020),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_806),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1020),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_807),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_812),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1020),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_813),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1020),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1020),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1029),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1029),
.Y(n_1177)
);

CKINVDCx16_ASAP7_75t_R g1178 ( 
.A(n_958),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1029),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_968),
.B(n_0),
.Y(n_1180)
);

CKINVDCx16_ASAP7_75t_R g1181 ( 
.A(n_982),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1029),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_814),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1029),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_779),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_710),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_816),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_815),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_714),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_841),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_860),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_715),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_751),
.B(n_888),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_734),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_786),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_861),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_982),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_716),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_722),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_795),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_734),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_725),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_728),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_867),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_762),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_762),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_729),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_818),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_730),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_802),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_735),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_745),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_819),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_810),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_809),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_748),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_830),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_750),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_755),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_821),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_823),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_756),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_766),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_769),
.Y(n_1224)
);

INVxp33_ASAP7_75t_L g1225 ( 
.A(n_778),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_780),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_825),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_784),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_790),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_796),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_826),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_820),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_713),
.B(n_2),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_828),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_822),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_827),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_810),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_829),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_831),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_838),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_840),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_844),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_982),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_832),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_833),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_837),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_850),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_852),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_835),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_859),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_853),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_728),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_839),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_854),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_842),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_843),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_855),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_846),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_811),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_847),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_863),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_848),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_811),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_874),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_851),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_868),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_877),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_856),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_858),
.Y(n_1269)
);

INVxp33_ASAP7_75t_SL g1270 ( 
.A(n_736),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_891),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_893),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_862),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_894),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_896),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_900),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_865),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_736),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_866),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_870),
.Y(n_1280)
);

INVxp67_ASAP7_75t_SL g1281 ( 
.A(n_845),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_908),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_924),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_929),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_845),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_933),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_939),
.Y(n_1287)
);

CKINVDCx14_ASAP7_75t_R g1288 ( 
.A(n_783),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_969),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_871),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_872),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_873),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_879),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_880),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_760),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_882),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_970),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_760),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_971),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_935),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_978),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_SL g1302 ( 
.A(n_783),
.Y(n_1302)
);

CKINVDCx16_ASAP7_75t_R g1303 ( 
.A(n_783),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_883),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_935),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_980),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_990),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_990),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_985),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_987),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_992),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_768),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_994),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_884),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_995),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_885),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_999),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_886),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1011),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1012),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_895),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1013),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1028),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1030),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_927),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1040),
.Y(n_1326)
);

XNOR2x1_ASAP7_75t_L g1327 ( 
.A(n_768),
.B(n_2),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1045),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1028),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_901),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_927),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_927),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_919),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_903),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_947),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_997),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_906),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_967),
.Y(n_1338)
);

CKINVDCx16_ASAP7_75t_R g1339 ( 
.A(n_997),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_909),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_997),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1002),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_888),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1002),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1002),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_770),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_993),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_993),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_912),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_916),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1032),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_917),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_920),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_921),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_876),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_923),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_925),
.Y(n_1357)
);

CKINVDCx14_ASAP7_75t_R g1358 ( 
.A(n_887),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_770),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_926),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_928),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_930),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1000),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_931),
.Y(n_1364)
);

CKINVDCx16_ASAP7_75t_R g1365 ( 
.A(n_1037),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1039),
.Y(n_1366)
);

BUFx8_ASAP7_75t_SL g1367 ( 
.A(n_1000),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_897),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_907),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_911),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_932),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_913),
.B(n_1),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_943),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1006),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_944),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_934),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_936),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_946),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_940),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_949),
.Y(n_1380)
);

CKINVDCx16_ASAP7_75t_R g1381 ( 
.A(n_711),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_950),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_953),
.B(n_1),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_955),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_941),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_956),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_959),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_961),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_962),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_942),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_963),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_973),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1006),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_975),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_977),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_983),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1007),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_948),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_951),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_957),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_960),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_976),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_979),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_981),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_712),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_712),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1007),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_717),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1021),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1070),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1140),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1109),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1138),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1141),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1367),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1109),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1050),
.B(n_1021),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1070),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1051),
.B(n_1376),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1149),
.Y(n_1421)
);

BUFx2_ASAP7_75t_SL g1422 ( 
.A(n_1377),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1144),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1146),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1151),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1156),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1203),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1157),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1159),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1153),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1160),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_1047),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1161),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1162),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1165),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1167),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1169),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1112),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1278),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1188),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1084),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1054),
.B(n_1056),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1190),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1084),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1105),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1172),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1047),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1054),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1353),
.B(n_1023),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1105),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1378),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1174),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1056),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1068),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1060),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1058),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1175),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1058),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1176),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1062),
.B(n_1023),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1068),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1062),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1177),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1063),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1179),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1060),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1112),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1115),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1354),
.B(n_1031),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1063),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1184),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1065),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1048),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1164),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1377),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1191),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1155),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1196),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1155),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1263),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1078),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1281),
.Y(n_1482)
);

NOR2xp67_ASAP7_75t_L g1483 ( 
.A(n_1204),
.B(n_1),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1046),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1164),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1356),
.B(n_1031),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1108),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1049),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1390),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1065),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1053),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1400),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1185),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1055),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1185),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1057),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1401),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1374),
.Y(n_1498)
);

NOR2xp67_ASAP7_75t_L g1499 ( 
.A(n_1346),
.B(n_2),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1083),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1064),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1358),
.B(n_1193),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1195),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1073),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1083),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1195),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1073),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1073),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1089),
.B(n_717),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1089),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1101),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1090),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1101),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1090),
.B(n_720),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1100),
.Y(n_1515)
);

INVxp33_ASAP7_75t_L g1516 ( 
.A(n_1393),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1101),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1123),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1123),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1071),
.Y(n_1520)
);

INVxp67_ASAP7_75t_SL g1521 ( 
.A(n_1078),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_1365),
.Y(n_1522)
);

CKINVDCx14_ASAP7_75t_R g1523 ( 
.A(n_1098),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1123),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1130),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1100),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1130),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1130),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1288),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1110),
.B(n_720),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1357),
.B(n_721),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1079),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1115),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1360),
.B(n_721),
.Y(n_1534)
);

BUFx10_ASAP7_75t_L g1535 ( 
.A(n_1302),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1110),
.B(n_723),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1088),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1111),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1163),
.Y(n_1539)
);

CKINVDCx16_ASAP7_75t_R g1540 ( 
.A(n_1099),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1163),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1111),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1182),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1182),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1186),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1189),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1200),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1192),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1200),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1198),
.Y(n_1550)
);

INVxp33_ASAP7_75t_SL g1551 ( 
.A(n_1080),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1210),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1079),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1118),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1199),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1210),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1202),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1207),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1209),
.Y(n_1559)
);

CKINVDCx16_ASAP7_75t_R g1560 ( 
.A(n_1158),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1118),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1249),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1215),
.Y(n_1563)
);

NOR2xp67_ASAP7_75t_L g1564 ( 
.A(n_1126),
.B(n_3),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1215),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1217),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1378),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1126),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1060),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1211),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1212),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1217),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1250),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1108),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1134),
.Y(n_1575)
);

CKINVDCx14_ASAP7_75t_R g1576 ( 
.A(n_1080),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1250),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1134),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1216),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1218),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1139),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1219),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1139),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1338),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1222),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1223),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1224),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1264),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1264),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1142),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1082),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1226),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1142),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1145),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1145),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1148),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1148),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1333),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1228),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1166),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1333),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1166),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1229),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1168),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1168),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1230),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1362),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1060),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1232),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1235),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1335),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1236),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1240),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1241),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1335),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1242),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1060),
.Y(n_1617)
);

NOR2xp67_ASAP7_75t_L g1618 ( 
.A(n_1170),
.B(n_3),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1247),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1351),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1248),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1251),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1170),
.B(n_723),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1171),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1171),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1254),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1257),
.Y(n_1627)
);

XNOR2xp5_ASAP7_75t_L g1628 ( 
.A(n_1351),
.B(n_1327),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1401),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1261),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1173),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1364),
.B(n_724),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1266),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1102),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1267),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1147),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1271),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1173),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1272),
.Y(n_1639)
);

INVxp33_ASAP7_75t_L g1640 ( 
.A(n_1295),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1366),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1298),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1183),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1274),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1183),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1275),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1373),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1276),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1282),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1187),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1283),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1284),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1178),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1181),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1187),
.B(n_724),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1286),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1208),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1287),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_L g1659 ( 
.A(n_1208),
.B(n_3),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1104),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1213),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1289),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1243),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1297),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1299),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1213),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1301),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1306),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1220),
.B(n_726),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1309),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1082),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1310),
.Y(n_1672)
);

CKINVDCx20_ASAP7_75t_R g1673 ( 
.A(n_1303),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1311),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_1331),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1375),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1313),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1315),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1220),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1221),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1221),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1339),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1317),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1131),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1319),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1320),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1312),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1227),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_R g1689 ( 
.A(n_1227),
.B(n_726),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_R g1690 ( 
.A(n_1231),
.B(n_731),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1231),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1234),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1322),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1359),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1104),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1381),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1234),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1238),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1324),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1326),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1328),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1104),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1128),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1129),
.Y(n_1704)
);

CKINVDCx16_ASAP7_75t_R g1705 ( 
.A(n_1302),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_1407),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1238),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1239),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1132),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1133),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1239),
.B(n_731),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1104),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1244),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1244),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1245),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1245),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1684),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1412),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1562),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1412),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1703),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1704),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1502),
.A2(n_1647),
.B1(n_1676),
.B2(n_1607),
.Y(n_1723)
);

INVx5_ASAP7_75t_L g1724 ( 
.A(n_1455),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1417),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1709),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1455),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1477),
.B(n_1368),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1710),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1417),
.Y(n_1730)
);

CKINVDCx6p67_ASAP7_75t_R g1731 ( 
.A(n_1540),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1545),
.Y(n_1732)
);

BUFx12f_ASAP7_75t_L g1733 ( 
.A(n_1416),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1432),
.B(n_1368),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1584),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_SL g1736 ( 
.A1(n_1628),
.A2(n_1059),
.B1(n_1270),
.B2(n_733),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1438),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1546),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1696),
.A2(n_1270),
.B1(n_733),
.B2(n_741),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1479),
.B(n_1369),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1438),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1487),
.B(n_1201),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1480),
.B(n_1369),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1467),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1467),
.Y(n_1745)
);

BUFx12f_ASAP7_75t_L g1746 ( 
.A(n_1416),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1468),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1487),
.B(n_1201),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1548),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1449),
.A2(n_1370),
.B1(n_1385),
.B2(n_1355),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1550),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1574),
.B(n_1451),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1455),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1422),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1555),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1574),
.B(n_1206),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1557),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1558),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1469),
.A2(n_1486),
.B1(n_1567),
.B2(n_1534),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1468),
.Y(n_1760)
);

INVx5_ASAP7_75t_L g1761 ( 
.A(n_1455),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1559),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1451),
.B(n_1206),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1570),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1539),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1447),
.B(n_1379),
.Y(n_1766)
);

OA21x2_ASAP7_75t_L g1767 ( 
.A1(n_1484),
.A2(n_1067),
.B(n_1066),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1641),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1696),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1413),
.A2(n_1052),
.B(n_1069),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1571),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1482),
.B(n_1379),
.Y(n_1772)
);

OAI22x1_ASAP7_75t_R g1773 ( 
.A1(n_1410),
.A2(n_737),
.B1(n_742),
.B2(n_741),
.Y(n_1773)
);

AND2x6_ASAP7_75t_L g1774 ( 
.A(n_1488),
.B(n_1398),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1454),
.B(n_1380),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1460),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1706),
.A2(n_737),
.B1(n_743),
.B2(n_742),
.Y(n_1778)
);

AND2x6_ASAP7_75t_L g1779 ( 
.A(n_1491),
.B(n_1399),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1494),
.A2(n_1074),
.B(n_1072),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1579),
.Y(n_1781)
);

AND2x6_ASAP7_75t_L g1782 ( 
.A(n_1496),
.B(n_1402),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1580),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1466),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1531),
.A2(n_1052),
.B(n_1069),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1466),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1582),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1466),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1585),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1461),
.B(n_1214),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1569),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1586),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1587),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1569),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1632),
.A2(n_1370),
.B1(n_1385),
.B2(n_1355),
.Y(n_1795)
);

INVx5_ASAP7_75t_L g1796 ( 
.A(n_1608),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1483),
.B(n_1246),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1539),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1481),
.A2(n_1076),
.B(n_1075),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1608),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1509),
.B(n_1246),
.Y(n_1801)
);

AOI22x1_ASAP7_75t_SL g1802 ( 
.A1(n_1410),
.A2(n_743),
.B1(n_749),
.B2(n_746),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1689),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1520),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1592),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1521),
.B(n_1384),
.Y(n_1806)
);

AND2x2_ASAP7_75t_SL g1807 ( 
.A(n_1514),
.B(n_1233),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1532),
.B(n_1214),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1617),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1541),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1427),
.A2(n_1409),
.B1(n_1407),
.B2(n_1106),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1553),
.B(n_1237),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1599),
.Y(n_1813)
);

OA21x2_ASAP7_75t_L g1814 ( 
.A1(n_1501),
.A2(n_1081),
.B(n_1077),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1617),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1660),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1603),
.B(n_1387),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1606),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1609),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1541),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1533),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1537),
.Y(n_1822)
);

AND2x2_ASAP7_75t_SL g1823 ( 
.A(n_1530),
.B(n_1372),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1536),
.B(n_1253),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1610),
.B(n_1388),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1504),
.B(n_1507),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1612),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1508),
.B(n_1391),
.Y(n_1828)
);

AND2x6_ASAP7_75t_L g1829 ( 
.A(n_1442),
.B(n_1403),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1642),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1543),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1511),
.B(n_1392),
.Y(n_1832)
);

INVx6_ASAP7_75t_L g1833 ( 
.A(n_1535),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1613),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1614),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1660),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1687),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_L g1838 ( 
.A1(n_1695),
.A2(n_1087),
.B(n_1086),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1616),
.B(n_1237),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1564),
.B(n_1180),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1694),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1544),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1695),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1619),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1623),
.B(n_1253),
.Y(n_1845)
);

OA21x2_ASAP7_75t_L g1846 ( 
.A1(n_1513),
.A2(n_1518),
.B(n_1517),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1621),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1702),
.Y(n_1848)
);

BUFx12f_ASAP7_75t_L g1849 ( 
.A(n_1535),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1622),
.B(n_1259),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1519),
.A2(n_1093),
.B(n_1092),
.Y(n_1851)
);

OA21x2_ASAP7_75t_L g1852 ( 
.A1(n_1524),
.A2(n_1300),
.B(n_1259),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1618),
.B(n_1255),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1655),
.A2(n_1255),
.B1(n_1258),
.B2(n_1256),
.Y(n_1854)
);

OAI21x1_ASAP7_75t_L g1855 ( 
.A1(n_1702),
.A2(n_1395),
.B(n_1394),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1525),
.B(n_1396),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1712),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1712),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1414),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1527),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1415),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1523),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1659),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1528),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1626),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1423),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1424),
.B(n_1404),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1627),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1426),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1428),
.B(n_1150),
.Y(n_1870)
);

OA21x2_ASAP7_75t_L g1871 ( 
.A1(n_1429),
.A2(n_1305),
.B(n_1300),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1669),
.A2(n_1256),
.B1(n_1260),
.B2(n_1258),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1431),
.Y(n_1873)
);

NAND2xp33_ASAP7_75t_L g1874 ( 
.A(n_1690),
.B(n_1260),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1439),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1630),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1633),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1635),
.B(n_1305),
.Y(n_1878)
);

INVx5_ASAP7_75t_L g1879 ( 
.A(n_1535),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1637),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1434),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1498),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1639),
.B(n_1308),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1435),
.B(n_1150),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1644),
.B(n_1308),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1711),
.B(n_1262),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1436),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1706),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1646),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1560),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1500),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1420),
.A2(n_1409),
.B1(n_1137),
.B2(n_1091),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1437),
.B(n_1104),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1419),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1446),
.Y(n_1895)
);

INVx5_ASAP7_75t_L g1896 ( 
.A(n_1705),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1648),
.B(n_1329),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1452),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1457),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1459),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1463),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1465),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1471),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1649),
.B(n_1143),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1651),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1652),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1529),
.B(n_1262),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1499),
.A2(n_1268),
.B1(n_1269),
.B2(n_1265),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1656),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1658),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1662),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1664),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1634),
.A2(n_1636),
.B1(n_1654),
.B2(n_1653),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1665),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1667),
.B(n_1329),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1668),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1670),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1672),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1419),
.Y(n_1919)
);

AND2x6_ASAP7_75t_L g1920 ( 
.A(n_1418),
.B(n_1405),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1674),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1677),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1505),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1678),
.Y(n_1924)
);

AND2x6_ASAP7_75t_L g1925 ( 
.A(n_1683),
.B(n_1406),
.Y(n_1925)
);

INVx5_ASAP7_75t_L g1926 ( 
.A(n_1522),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1685),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1576),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1686),
.B(n_1693),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1699),
.B(n_1700),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1701),
.B(n_1094),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1421),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1516),
.B(n_1408),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1640),
.B(n_1135),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1688),
.B(n_1095),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1713),
.B(n_1096),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1425),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1430),
.B(n_1143),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1715),
.Y(n_1939)
);

BUFx8_ASAP7_75t_L g1940 ( 
.A(n_1475),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1433),
.B(n_1143),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1472),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1440),
.B(n_1143),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1443),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1448),
.A2(n_1268),
.B1(n_1269),
.B2(n_1265),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1478),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1489),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1490),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1591),
.Y(n_1949)
);

BUFx8_ASAP7_75t_L g1950 ( 
.A(n_1497),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1671),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1492),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1510),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1476),
.B(n_1273),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1512),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1476),
.B(n_1097),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1515),
.B(n_1136),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1526),
.B(n_1273),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1538),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1526),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1624),
.B(n_1277),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1542),
.B(n_1119),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1554),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1561),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1568),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1575),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1578),
.B(n_1119),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1624),
.B(n_1277),
.Y(n_1968)
);

OA21x2_ASAP7_75t_L g1969 ( 
.A1(n_1716),
.A2(n_1348),
.B(n_1343),
.Y(n_1969)
);

OAI22x1_ASAP7_75t_L g1970 ( 
.A1(n_1625),
.A2(n_1061),
.B1(n_1197),
.B2(n_1325),
.Y(n_1970)
);

CKINVDCx6p67_ASAP7_75t_R g1971 ( 
.A(n_1634),
.Y(n_1971)
);

OA21x2_ASAP7_75t_L g1972 ( 
.A1(n_1625),
.A2(n_1348),
.B(n_1343),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1581),
.B(n_1103),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1583),
.Y(n_1974)
);

INVx5_ASAP7_75t_L g1975 ( 
.A(n_1551),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1590),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1593),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1594),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1595),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1596),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1597),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1600),
.B(n_1085),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1551),
.A2(n_1279),
.B1(n_1290),
.B2(n_1280),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1602),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1604),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1605),
.B(n_1107),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1650),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1657),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1679),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1680),
.B(n_1113),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1681),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1707),
.B(n_1143),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1708),
.Y(n_1993)
);

OAI21x1_ASAP7_75t_L g1994 ( 
.A1(n_1631),
.A2(n_1347),
.B(n_1116),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1631),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1638),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1638),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1643),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1643),
.B(n_1152),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1645),
.B(n_1114),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1645),
.B(n_1117),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1661),
.Y(n_2002)
);

BUFx3_ASAP7_75t_L g2003 ( 
.A(n_1661),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1666),
.A2(n_1121),
.B(n_1120),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_L g2005 ( 
.A1(n_1666),
.A2(n_1124),
.B(n_1122),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1691),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1823),
.A2(n_1692),
.B1(n_1697),
.B2(n_1691),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1823),
.A2(n_1807),
.B1(n_1759),
.B2(n_1920),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1807),
.A2(n_1920),
.B1(n_1829),
.B2(n_1723),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1920),
.A2(n_1697),
.B1(n_1698),
.B2(n_1692),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1717),
.B(n_1719),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1840),
.A2(n_1280),
.B1(n_1290),
.B2(n_1279),
.Y(n_2012)
);

INVx3_ASAP7_75t_SL g2013 ( 
.A(n_1862),
.Y(n_2013)
);

OA22x2_ASAP7_75t_L g2014 ( 
.A1(n_1778),
.A2(n_1970),
.B1(n_1983),
.B2(n_1872),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1718),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1718),
.Y(n_2016)
);

AO22x2_ASAP7_75t_L g2017 ( 
.A1(n_1892),
.A2(n_1327),
.B1(n_1811),
.B2(n_1802),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1920),
.A2(n_1714),
.B1(n_1716),
.B2(n_1698),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1720),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1776),
.B(n_1714),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1920),
.A2(n_1453),
.B1(n_1456),
.B2(n_1448),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1920),
.A2(n_1456),
.B1(n_1458),
.B2(n_1453),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1717),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1735),
.B(n_1291),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1871),
.Y(n_2025)
);

AO22x2_ASAP7_75t_L g2026 ( 
.A1(n_1750),
.A2(n_824),
.B1(n_857),
.B2(n_727),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1768),
.B(n_1291),
.Y(n_2027)
);

OAI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1734),
.A2(n_1766),
.B1(n_1806),
.B2(n_1775),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1829),
.A2(n_1462),
.B1(n_1464),
.B2(n_1458),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1829),
.A2(n_1464),
.B1(n_1470),
.B2(n_1462),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1934),
.B(n_1292),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1742),
.B(n_1125),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1720),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1934),
.B(n_1292),
.Y(n_2034)
);

XNOR2xp5_ASAP7_75t_L g2035 ( 
.A(n_1913),
.B(n_1441),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1933),
.B(n_1293),
.Y(n_2036)
);

AOI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1829),
.A2(n_1470),
.B1(n_1294),
.B2(n_1296),
.Y(n_2037)
);

OAI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_1840),
.A2(n_1294),
.B1(n_1296),
.B2(n_1293),
.Y(n_2038)
);

AOI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1790),
.A2(n_1383),
.B1(n_1314),
.B2(n_1316),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1871),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1725),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1725),
.Y(n_2042)
);

AO22x2_ASAP7_75t_L g2043 ( 
.A1(n_1795),
.A2(n_915),
.B1(n_918),
.B2(n_910),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1933),
.B(n_1304),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_SL g2045 ( 
.A(n_1928),
.B(n_1473),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_SL g2046 ( 
.A1(n_1736),
.A2(n_1629),
.B1(n_1444),
.B2(n_1445),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1829),
.A2(n_1304),
.B1(n_1316),
.B2(n_1314),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1871),
.Y(n_2048)
);

CKINVDCx6p67_ASAP7_75t_R g2049 ( 
.A(n_1926),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_SL g2050 ( 
.A1(n_1840),
.A2(n_1853),
.B1(n_1797),
.B2(n_1999),
.Y(n_2050)
);

OAI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1840),
.A2(n_1854),
.B1(n_1914),
.B2(n_1910),
.Y(n_2051)
);

OAI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1910),
.A2(n_1321),
.B1(n_1330),
.B2(n_1318),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1875),
.B(n_1363),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1829),
.A2(n_1318),
.B1(n_1330),
.B2(n_1321),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1852),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_1801),
.A2(n_1334),
.B1(n_1340),
.B2(n_1337),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1852),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1982),
.B(n_1334),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1730),
.Y(n_2059)
);

OAI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1910),
.A2(n_1340),
.B1(n_1352),
.B2(n_1337),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_1763),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_SL g2062 ( 
.A1(n_1894),
.A2(n_1629),
.B1(n_1444),
.B2(n_1445),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1730),
.Y(n_2063)
);

OAI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1914),
.A2(n_1361),
.B1(n_1371),
.B2(n_1352),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1824),
.A2(n_1361),
.B1(n_1386),
.B2(n_1371),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1737),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1982),
.B(n_1386),
.Y(n_2067)
);

INVx3_ASAP7_75t_L g2068 ( 
.A(n_1742),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1737),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1741),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1803),
.B(n_1389),
.Y(n_2071)
);

OR2x6_ASAP7_75t_L g2072 ( 
.A(n_1946),
.B(n_1332),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1803),
.B(n_1389),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1845),
.A2(n_1886),
.B1(n_1808),
.B2(n_1812),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1852),
.Y(n_2075)
);

OAI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1914),
.A2(n_1017),
.B1(n_1024),
.B2(n_954),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1875),
.B(n_1154),
.Y(n_2077)
);

AO22x2_ASAP7_75t_L g2078 ( 
.A1(n_1945),
.A2(n_1336),
.B1(n_1342),
.B2(n_1341),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1742),
.Y(n_2079)
);

AO22x2_ASAP7_75t_L g2080 ( 
.A1(n_1995),
.A2(n_1344),
.B1(n_1345),
.B2(n_1127),
.Y(n_2080)
);

AND2x2_ASAP7_75t_SL g2081 ( 
.A(n_1891),
.B(n_1441),
.Y(n_2081)
);

AO22x2_ASAP7_75t_L g2082 ( 
.A1(n_1995),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2082)
);

OR2x6_ASAP7_75t_L g2083 ( 
.A(n_1946),
.B(n_1450),
.Y(n_2083)
);

OAI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1863),
.A2(n_749),
.B1(n_752),
.B2(n_746),
.Y(n_2084)
);

OAI22xp33_ASAP7_75t_SL g2085 ( 
.A1(n_1853),
.A2(n_753),
.B1(n_757),
.B2(n_752),
.Y(n_2085)
);

NAND3x1_ASAP7_75t_L g2086 ( 
.A(n_1954),
.B(n_1653),
.C(n_1636),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1790),
.A2(n_1473),
.B1(n_1302),
.B2(n_1673),
.Y(n_2087)
);

NAND3x1_ASAP7_75t_L g2088 ( 
.A(n_1996),
.B(n_1663),
.C(n_1654),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1748),
.Y(n_2089)
);

AO22x2_ASAP7_75t_L g2090 ( 
.A1(n_2006),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1790),
.A2(n_1673),
.B1(n_1682),
.B2(n_1675),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1741),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1918),
.A2(n_757),
.B1(n_758),
.B2(n_753),
.Y(n_2093)
);

OA22x2_ASAP7_75t_L g2094 ( 
.A1(n_1970),
.A2(n_984),
.B1(n_1008),
.B2(n_758),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1808),
.A2(n_1675),
.B1(n_1682),
.B2(n_1663),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1962),
.B(n_1252),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1962),
.B(n_1252),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_SL g2098 ( 
.A1(n_1894),
.A2(n_1474),
.B1(n_1485),
.B2(n_1450),
.Y(n_2098)
);

AO22x2_ASAP7_75t_L g2099 ( 
.A1(n_2006),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2099)
);

OAI22xp33_ASAP7_75t_SL g2100 ( 
.A1(n_1797),
.A2(n_763),
.B1(n_765),
.B2(n_759),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1838),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1808),
.A2(n_1205),
.B1(n_1285),
.B2(n_1194),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1744),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1838),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_1812),
.A2(n_1205),
.B1(n_1285),
.B2(n_1194),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1744),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1745),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1748),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_1918),
.A2(n_763),
.B1(n_765),
.B2(n_759),
.Y(n_2109)
);

AOI22x1_ASAP7_75t_L g2110 ( 
.A1(n_1728),
.A2(n_878),
.B1(n_890),
.B2(n_767),
.Y(n_2110)
);

AOI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1812),
.A2(n_1957),
.B1(n_1956),
.B2(n_2000),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_1748),
.B(n_1756),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_1957),
.A2(n_1205),
.B1(n_1285),
.B2(n_1194),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_1956),
.A2(n_1205),
.B1(n_1285),
.B2(n_1194),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1745),
.Y(n_2115)
);

XNOR2xp5_ASAP7_75t_L g2116 ( 
.A(n_1919),
.B(n_1474),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1747),
.Y(n_2117)
);

OA22x2_ASAP7_75t_L g2118 ( 
.A1(n_1935),
.A2(n_998),
.B1(n_1016),
.B2(n_767),
.Y(n_2118)
);

AO22x2_ASAP7_75t_L g2119 ( 
.A1(n_1908),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1967),
.B(n_1252),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1967),
.B(n_1397),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1747),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1756),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1760),
.Y(n_2124)
);

OAI22xp5_ASAP7_75t_SL g2125 ( 
.A1(n_1919),
.A2(n_1493),
.B1(n_1495),
.B2(n_1485),
.Y(n_2125)
);

OAI22xp33_ASAP7_75t_SL g2126 ( 
.A1(n_1732),
.A2(n_890),
.B1(n_892),
.B2(n_878),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1756),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_1846),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1760),
.Y(n_2129)
);

AOI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1956),
.A2(n_1205),
.B1(n_1285),
.B2(n_1194),
.Y(n_2130)
);

INVx2_ASAP7_75t_SL g2131 ( 
.A(n_1763),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1763),
.B(n_1397),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1765),
.Y(n_2133)
);

OAI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1918),
.A2(n_1225),
.B1(n_984),
.B2(n_988),
.Y(n_2134)
);

OR2x6_ASAP7_75t_L g2135 ( 
.A(n_1946),
.B(n_1493),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_1973),
.Y(n_2136)
);

OAI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_1828),
.A2(n_988),
.B1(n_991),
.B2(n_892),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1765),
.Y(n_2138)
);

OAI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_1832),
.A2(n_996),
.B1(n_998),
.B2(n_991),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2000),
.B(n_1397),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1798),
.Y(n_2141)
);

AOI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2000),
.A2(n_2001),
.B1(n_1772),
.B2(n_1743),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2001),
.B(n_996),
.Y(n_2143)
);

OAI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_1856),
.A2(n_1004),
.B1(n_1005),
.B2(n_1001),
.Y(n_2144)
);

AND2x2_ASAP7_75t_SL g2145 ( 
.A(n_1891),
.B(n_1495),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1928),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2001),
.A2(n_1323),
.B1(n_1307),
.B2(n_1004),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1873),
.B(n_1887),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1969),
.A2(n_1005),
.B1(n_1008),
.B2(n_1001),
.Y(n_2149)
);

AOI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1743),
.A2(n_1323),
.B1(n_1307),
.B2(n_1014),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1873),
.B(n_1307),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1772),
.A2(n_1323),
.B1(n_1307),
.B2(n_1014),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_SL g2153 ( 
.A(n_1997),
.B(n_1009),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1798),
.Y(n_2154)
);

OAI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1929),
.A2(n_1930),
.B1(n_1905),
.B2(n_1909),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_1769),
.Y(n_2156)
);

CKINVDCx14_ASAP7_75t_R g2157 ( 
.A(n_1731),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1810),
.Y(n_2158)
);

OAI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_1905),
.A2(n_1015),
.B1(n_1016),
.B2(n_1009),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1973),
.B(n_1015),
.Y(n_2160)
);

NOR2x1p5_ASAP7_75t_L g2161 ( 
.A(n_1849),
.B(n_1026),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1973),
.A2(n_1323),
.B1(n_1307),
.B2(n_1027),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1810),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1986),
.B(n_1990),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1986),
.A2(n_1323),
.B1(n_1027),
.B2(n_1033),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1820),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1986),
.B(n_1026),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_1990),
.A2(n_1035),
.B1(n_1036),
.B2(n_1033),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1990),
.B(n_1035),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_1935),
.A2(n_1936),
.B1(n_1777),
.B2(n_1825),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1820),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1864),
.Y(n_2172)
);

OAI22xp5_ASAP7_75t_SL g2173 ( 
.A1(n_1739),
.A2(n_1506),
.B1(n_1547),
.B2(n_1503),
.Y(n_2173)
);

BUFx3_ASAP7_75t_L g2174 ( 
.A(n_1946),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1846),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1935),
.B(n_1036),
.Y(n_2176)
);

OAI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_1738),
.A2(n_1751),
.B1(n_1755),
.B2(n_1749),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1864),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1936),
.A2(n_1041),
.B1(n_1042),
.B2(n_1038),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1936),
.B(n_1038),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1821),
.Y(n_2181)
);

AOI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_1777),
.A2(n_1042),
.B1(n_1043),
.B2(n_1041),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1752),
.B(n_1043),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1846),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1752),
.B(n_1044),
.Y(n_2185)
);

AO22x2_ASAP7_75t_L g2186 ( 
.A1(n_1958),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2186)
);

OAI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_1906),
.A2(n_1044),
.B1(n_1506),
.B2(n_1503),
.Y(n_2187)
);

OA22x2_ASAP7_75t_L g2188 ( 
.A1(n_1939),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2188)
);

BUFx4f_ASAP7_75t_L g2189 ( 
.A(n_1946),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_1882),
.B(n_10),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_1939),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_1752),
.B(n_1547),
.Y(n_2192)
);

OAI22xp33_ASAP7_75t_SL g2193 ( 
.A1(n_1757),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1996),
.B(n_1563),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1821),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1831),
.Y(n_2196)
);

OAI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_1906),
.A2(n_1552),
.B1(n_1556),
.B2(n_1549),
.Y(n_2197)
);

CKINVDCx6p67_ASAP7_75t_R g2198 ( 
.A(n_1926),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_1817),
.A2(n_1152),
.B1(n_1150),
.B2(n_1549),
.Y(n_2199)
);

OA22x2_ASAP7_75t_L g2200 ( 
.A1(n_1942),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1831),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_1916),
.B(n_13),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_1839),
.Y(n_2203)
);

OAI22xp33_ASAP7_75t_L g2204 ( 
.A1(n_1909),
.A2(n_1556),
.B1(n_1563),
.B2(n_1552),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1996),
.B(n_1588),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_1839),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_SL g2207 ( 
.A1(n_1769),
.A2(n_1566),
.B1(n_1572),
.B2(n_1565),
.Y(n_2207)
);

AO22x2_ASAP7_75t_L g2208 ( 
.A1(n_1958),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_2208)
);

OAI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_1912),
.A2(n_1566),
.B1(n_1572),
.B2(n_1565),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_SL g2210 ( 
.A1(n_1888),
.A2(n_1577),
.B1(n_1588),
.B2(n_1573),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1842),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1817),
.A2(n_1825),
.B1(n_1925),
.B2(n_1740),
.Y(n_2212)
);

OAI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_1912),
.A2(n_1577),
.B1(n_1589),
.B2(n_1573),
.Y(n_2213)
);

AO22x2_ASAP7_75t_L g2214 ( 
.A1(n_1961),
.A2(n_1968),
.B1(n_1977),
.B2(n_1955),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_1925),
.A2(n_1152),
.B1(n_1150),
.B2(n_1589),
.Y(n_2215)
);

INVx2_ASAP7_75t_SL g2216 ( 
.A(n_1728),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1842),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1873),
.B(n_1150),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1916),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1881),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_1979),
.B(n_1598),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1843),
.Y(n_2222)
);

OAI22xp33_ASAP7_75t_SL g2223 ( 
.A1(n_1758),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_2223)
);

OR2x6_ASAP7_75t_L g2224 ( 
.A(n_1947),
.B(n_1598),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1979),
.B(n_1601),
.Y(n_2225)
);

AOI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_1925),
.A2(n_1152),
.B1(n_1611),
.B2(n_1601),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_1925),
.A2(n_1152),
.B1(n_1615),
.B2(n_1611),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_1804),
.B(n_16),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1881),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1925),
.A2(n_1620),
.B1(n_1615),
.B2(n_146),
.Y(n_2230)
);

AO22x2_ASAP7_75t_L g2231 ( 
.A1(n_1961),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1887),
.B(n_17),
.Y(n_2232)
);

OR2x6_ASAP7_75t_L g2233 ( 
.A(n_1947),
.B(n_1620),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1898),
.Y(n_2234)
);

OAI22xp33_ASAP7_75t_R g2235 ( 
.A1(n_1773),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1740),
.B(n_705),
.Y(n_2236)
);

AO22x2_ASAP7_75t_L g2237 ( 
.A1(n_1968),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_1822),
.B(n_20),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_1830),
.B(n_21),
.Y(n_2239)
);

OAI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_1917),
.A2(n_1921),
.B1(n_1924),
.B2(n_1922),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1843),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1857),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1964),
.B(n_145),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1964),
.B(n_692),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_1923),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_1925),
.A2(n_147),
.B1(n_148),
.B2(n_146),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_1901),
.A2(n_149),
.B1(n_150),
.B2(n_147),
.Y(n_2247)
);

AO22x2_ASAP7_75t_L g2248 ( 
.A1(n_1984),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1964),
.B(n_698),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1837),
.B(n_1841),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1762),
.A2(n_151),
.B1(n_152),
.B2(n_149),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_1764),
.A2(n_1781),
.B1(n_1783),
.B2(n_1771),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1857),
.Y(n_2253)
);

XOR2xp5_ASAP7_75t_L g2254 ( 
.A(n_1890),
.B(n_151),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1981),
.B(n_700),
.Y(n_2255)
);

OR2x6_ASAP7_75t_L g2256 ( 
.A(n_1947),
.B(n_22),
.Y(n_2256)
);

OAI22xp5_ASAP7_75t_SL g2257 ( 
.A1(n_1888),
.A2(n_31),
.B1(n_39),
.B2(n_23),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1858),
.Y(n_2258)
);

OAI22xp33_ASAP7_75t_SL g2259 ( 
.A1(n_1787),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2259)
);

AO22x2_ASAP7_75t_L g2260 ( 
.A1(n_1985),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2260)
);

OAI22xp33_ASAP7_75t_SL g2261 ( 
.A1(n_1789),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_1981),
.B(n_706),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_1948),
.B(n_26),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1981),
.B(n_709),
.Y(n_2264)
);

OR2x6_ASAP7_75t_L g2265 ( 
.A(n_1947),
.B(n_28),
.Y(n_2265)
);

OAI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_1917),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2266)
);

OAI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_1921),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2267)
);

AOI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_1792),
.A2(n_154),
.B1(n_155),
.B2(n_152),
.Y(n_2268)
);

OAI22xp33_ASAP7_75t_SL g2269 ( 
.A1(n_1793),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_1975),
.B(n_1923),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1858),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_1975),
.B(n_694),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_1949),
.B(n_32),
.Y(n_2273)
);

OAI22xp33_ASAP7_75t_SL g2274 ( 
.A1(n_1805),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1975),
.B(n_697),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1860),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_1813),
.A2(n_155),
.B1(n_156),
.B2(n_154),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_1818),
.A2(n_157),
.B1(n_158),
.B2(n_156),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1898),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_1819),
.A2(n_158),
.B1(n_159),
.B2(n_157),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1975),
.B(n_702),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1860),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1922),
.Y(n_2283)
);

OAI22xp33_ASAP7_75t_SL g2284 ( 
.A1(n_1827),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1860),
.Y(n_2285)
);

OAI22xp33_ASAP7_75t_SL g2286 ( 
.A1(n_1834),
.A2(n_37),
.B1(n_33),
.B2(n_36),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_1975),
.B(n_707),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_SL g2288 ( 
.A1(n_1960),
.A2(n_1976),
.B1(n_1993),
.B2(n_1754),
.Y(n_2288)
);

OR2x2_ASAP7_75t_L g2289 ( 
.A(n_1951),
.B(n_36),
.Y(n_2289)
);

OAI22xp5_ASAP7_75t_SL g2290 ( 
.A1(n_1976),
.A2(n_45),
.B1(n_53),
.B2(n_37),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1851),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1924),
.Y(n_2292)
);

AOI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_1835),
.A2(n_160),
.B1(n_161),
.B2(n_159),
.Y(n_2293)
);

OAI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_1867),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1839),
.Y(n_2295)
);

OAI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_1844),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_1847),
.A2(n_1868),
.B1(n_1876),
.B2(n_1865),
.Y(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_1877),
.A2(n_1889),
.B1(n_1880),
.B2(n_1722),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_1874),
.A2(n_162),
.B1(n_163),
.B2(n_161),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_1879),
.B(n_38),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_1993),
.B(n_694),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1887),
.B(n_40),
.Y(n_2302)
);

OR2x6_ASAP7_75t_L g2303 ( 
.A(n_1947),
.B(n_41),
.Y(n_2303)
);

OAI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_1969),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2304)
);

AOI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_1874),
.A2(n_163),
.B1(n_164),
.B2(n_162),
.Y(n_2305)
);

OAI22xp33_ASAP7_75t_SL g2306 ( 
.A1(n_1992),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2306)
);

AO22x2_ASAP7_75t_L g2307 ( 
.A1(n_1989),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2307)
);

XNOR2x2_ASAP7_75t_SL g2308 ( 
.A(n_1971),
.B(n_46),
.Y(n_2308)
);

OAI22xp33_ASAP7_75t_SL g2309 ( 
.A1(n_1721),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_1959),
.B(n_704),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_1959),
.B(n_707),
.Y(n_2311)
);

AOI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_1903),
.A2(n_1726),
.B1(n_1729),
.B2(n_1774),
.Y(n_2312)
);

AO22x2_ASAP7_75t_L g2313 ( 
.A1(n_1963),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2313)
);

AO22x2_ASAP7_75t_L g2314 ( 
.A1(n_1963),
.A2(n_1978),
.B1(n_1980),
.B2(n_1966),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_1903),
.A2(n_166),
.B1(n_167),
.B2(n_164),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1851),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1895),
.B(n_48),
.Y(n_2317)
);

AOI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_1903),
.A2(n_168),
.B1(n_169),
.B2(n_167),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_L g2319 ( 
.A(n_1938),
.B(n_49),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1851),
.Y(n_2320)
);

OAI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_1944),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2321)
);

OAI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_1944),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_SL g2323 ( 
.A1(n_1754),
.A2(n_58),
.B1(n_66),
.B2(n_50),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_1969),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1850),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1850),
.Y(n_2326)
);

AOI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_1774),
.A2(n_169),
.B1(n_170),
.B2(n_168),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2295),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2008),
.B(n_1997),
.Y(n_2329)
);

AOI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2186),
.A2(n_1972),
.B1(n_1780),
.B2(n_1814),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2074),
.B(n_1972),
.Y(n_2331)
);

INVx1_ASAP7_75t_SL g2332 ( 
.A(n_2011),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2053),
.B(n_1974),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2020),
.B(n_2036),
.Y(n_2334)
);

BUFx10_ASAP7_75t_L g2335 ( 
.A(n_2146),
.Y(n_2335)
);

XNOR2xp5_ASAP7_75t_L g2336 ( 
.A(n_2116),
.B(n_1890),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2044),
.B(n_1932),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2107),
.Y(n_2338)
);

OR2x2_ASAP7_75t_L g2339 ( 
.A(n_2023),
.B(n_2003),
.Y(n_2339)
);

INVx2_ASAP7_75t_SL g2340 ( 
.A(n_2192),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_2191),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2031),
.B(n_2034),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2028),
.B(n_1972),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2325),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2009),
.B(n_1997),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2326),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2089),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2276),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2107),
.Y(n_2349)
);

BUFx3_ASAP7_75t_L g2350 ( 
.A(n_2174),
.Y(n_2350)
);

BUFx4f_ASAP7_75t_L g2351 ( 
.A(n_2049),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_2089),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2050),
.B(n_1997),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2276),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2089),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2282),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2282),
.Y(n_2357)
);

AND3x2_ASAP7_75t_L g2358 ( 
.A(n_2045),
.B(n_1978),
.C(n_1966),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2117),
.Y(n_2359)
);

NAND2xp33_ASAP7_75t_SL g2360 ( 
.A(n_2164),
.B(n_2002),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2285),
.Y(n_2361)
);

BUFx3_ASAP7_75t_L g2362 ( 
.A(n_2189),
.Y(n_2362)
);

INVxp67_ASAP7_75t_SL g2363 ( 
.A(n_2108),
.Y(n_2363)
);

INVx5_ASAP7_75t_L g2364 ( 
.A(n_2128),
.Y(n_2364)
);

AOI22xp33_ASAP7_75t_L g2365 ( 
.A1(n_2186),
.A2(n_1780),
.B1(n_1814),
.B2(n_1767),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2216),
.B(n_1941),
.Y(n_2366)
);

AND2x6_ASAP7_75t_L g2367 ( 
.A(n_2175),
.B(n_1997),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2285),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2117),
.Y(n_2369)
);

BUFx6f_ASAP7_75t_L g2370 ( 
.A(n_2108),
.Y(n_2370)
);

AND2x4_ASAP7_75t_L g2371 ( 
.A(n_2112),
.B(n_2004),
.Y(n_2371)
);

NAND2xp33_ASAP7_75t_L g2372 ( 
.A(n_2212),
.B(n_1774),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2068),
.Y(n_2373)
);

INVx6_ASAP7_75t_L g2374 ( 
.A(n_2108),
.Y(n_2374)
);

OR2x2_ASAP7_75t_L g2375 ( 
.A(n_2077),
.B(n_2003),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2189),
.B(n_1998),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2155),
.B(n_1943),
.Y(n_2377)
);

AOI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_2208),
.A2(n_2231),
.B1(n_2237),
.B2(n_2188),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2129),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2129),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_2024),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2068),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2123),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2154),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2154),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2245),
.Y(n_2386)
);

INVxp67_ASAP7_75t_SL g2387 ( 
.A(n_2127),
.Y(n_2387)
);

NAND2xp33_ASAP7_75t_SL g2388 ( 
.A(n_2270),
.B(n_1998),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2051),
.B(n_2111),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2123),
.Y(n_2390)
);

INVxp67_ASAP7_75t_SL g2391 ( 
.A(n_2127),
.Y(n_2391)
);

INVx3_ASAP7_75t_L g2392 ( 
.A(n_2127),
.Y(n_2392)
);

NAND2xp33_ASAP7_75t_L g2393 ( 
.A(n_2272),
.B(n_1774),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2157),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2061),
.B(n_1927),
.Y(n_2395)
);

INVxp33_ASAP7_75t_L g2396 ( 
.A(n_2027),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2163),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2163),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2131),
.B(n_1927),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_2112),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2203),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2203),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2206),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2171),
.Y(n_2404)
);

INVx4_ASAP7_75t_L g2405 ( 
.A(n_2219),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2171),
.Y(n_2406)
);

CKINVDCx16_ASAP7_75t_R g2407 ( 
.A(n_2098),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2058),
.B(n_1998),
.Y(n_2408)
);

OR2x6_ASAP7_75t_L g2409 ( 
.A(n_2083),
.B(n_1733),
.Y(n_2409)
);

BUFx10_ASAP7_75t_L g2410 ( 
.A(n_2238),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2206),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_2067),
.B(n_1932),
.Y(n_2412)
);

AOI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_2208),
.A2(n_1780),
.B1(n_1814),
.B2(n_1767),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2195),
.Y(n_2414)
);

INVx5_ASAP7_75t_L g2415 ( 
.A(n_2128),
.Y(n_2415)
);

INVx4_ASAP7_75t_L g2416 ( 
.A(n_2219),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2142),
.B(n_1927),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_SL g2418 ( 
.A(n_2170),
.B(n_1998),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2195),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2025),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2025),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2196),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2040),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2040),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2196),
.Y(n_2425)
);

NOR2x1p5_ASAP7_75t_L g2426 ( 
.A(n_2198),
.B(n_1731),
.Y(n_2426)
);

INVx4_ASAP7_75t_L g2427 ( 
.A(n_2219),
.Y(n_2427)
);

CKINVDCx20_ASAP7_75t_R g2428 ( 
.A(n_2062),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_2079),
.Y(n_2429)
);

AOI22xp33_ASAP7_75t_L g2430 ( 
.A1(n_2231),
.A2(n_1767),
.B1(n_1779),
.B2(n_1774),
.Y(n_2430)
);

OAI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2256),
.A2(n_1998),
.B1(n_2002),
.B2(n_1988),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2048),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2211),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2214),
.A2(n_1774),
.B1(n_1782),
.B2(n_1779),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2211),
.Y(n_2435)
);

NOR2x1p5_ASAP7_75t_L g2436 ( 
.A(n_2140),
.B(n_1849),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_2013),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2217),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2217),
.Y(n_2439)
);

AND2x6_ASAP7_75t_L g2440 ( 
.A(n_2175),
.B(n_2002),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2096),
.B(n_2002),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2222),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2222),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2236),
.B(n_2220),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2229),
.B(n_1927),
.Y(n_2445)
);

CKINVDCx6p67_ASAP7_75t_R g2446 ( 
.A(n_2083),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2048),
.Y(n_2447)
);

NAND2xp33_ASAP7_75t_R g2448 ( 
.A(n_2156),
.B(n_1862),
.Y(n_2448)
);

AOI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2214),
.A2(n_1779),
.B1(n_1782),
.B2(n_1980),
.Y(n_2449)
);

INVx1_ASAP7_75t_SL g2450 ( 
.A(n_2221),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_2234),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2055),
.Y(n_2452)
);

OR2x6_ASAP7_75t_L g2453 ( 
.A(n_2135),
.B(n_2224),
.Y(n_2453)
);

INVx4_ASAP7_75t_L g2454 ( 
.A(n_2202),
.Y(n_2454)
);

INVx11_ASAP7_75t_L g2455 ( 
.A(n_2135),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2241),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2279),
.B(n_1927),
.Y(n_2457)
);

AND2x6_ASAP7_75t_L g2458 ( 
.A(n_2291),
.B(n_2002),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2071),
.B(n_1932),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2283),
.B(n_2292),
.Y(n_2460)
);

OR2x6_ASAP7_75t_L g2461 ( 
.A(n_2224),
.B(n_1733),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2202),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2055),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2241),
.Y(n_2464)
);

AND2x6_ASAP7_75t_L g2465 ( 
.A(n_2291),
.B(n_1988),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2225),
.Y(n_2466)
);

INVx5_ASAP7_75t_L g2467 ( 
.A(n_2184),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2242),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2125),
.Y(n_2469)
);

INVxp33_ASAP7_75t_L g2470 ( 
.A(n_2250),
.Y(n_2470)
);

NAND3xp33_ASAP7_75t_L g2471 ( 
.A(n_2056),
.B(n_1987),
.C(n_1965),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2181),
.Y(n_2472)
);

AND2x2_ASAP7_75t_SL g2473 ( 
.A(n_2081),
.B(n_1988),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2057),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2242),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2253),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2253),
.Y(n_2477)
);

AOI22xp33_ASAP7_75t_L g2478 ( 
.A1(n_2237),
.A2(n_1779),
.B1(n_1782),
.B2(n_1897),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2097),
.B(n_1988),
.Y(n_2479)
);

OR2x6_ASAP7_75t_L g2480 ( 
.A(n_2233),
.B(n_1746),
.Y(n_2480)
);

INVx5_ASAP7_75t_L g2481 ( 
.A(n_2184),
.Y(n_2481)
);

INVx5_ASAP7_75t_L g2482 ( 
.A(n_2275),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2032),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2073),
.B(n_2120),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2258),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2201),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2319),
.B(n_1895),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2057),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2258),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2271),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2271),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2148),
.B(n_1895),
.Y(n_2492)
);

BUFx10_ASAP7_75t_L g2493 ( 
.A(n_2239),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2172),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2178),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2032),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2015),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2121),
.B(n_1988),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2075),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2240),
.B(n_1911),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2065),
.B(n_1987),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_2310),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2243),
.B(n_1911),
.Y(n_2503)
);

AOI22xp33_ASAP7_75t_L g2504 ( 
.A1(n_2200),
.A2(n_1779),
.B1(n_1782),
.B2(n_1897),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2016),
.Y(n_2505)
);

INVx4_ASAP7_75t_L g2506 ( 
.A(n_2072),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2244),
.B(n_2249),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2019),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_2233),
.Y(n_2509)
);

XNOR2xp5_ASAP7_75t_L g2510 ( 
.A(n_2086),
.B(n_1907),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2075),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2033),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2101),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2041),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2281),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2132),
.B(n_1953),
.Y(n_2516)
);

INVx4_ASAP7_75t_L g2517 ( 
.A(n_2072),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2042),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2136),
.B(n_1953),
.Y(n_2519)
);

BUFx10_ASAP7_75t_L g2520 ( 
.A(n_2145),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2101),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2104),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2104),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2059),
.Y(n_2524)
);

NAND2xp33_ASAP7_75t_SL g2525 ( 
.A(n_2255),
.B(n_1953),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2313),
.A2(n_1779),
.B1(n_1782),
.B2(n_1931),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_2063),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2066),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2069),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2070),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2092),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2007),
.B(n_1952),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2103),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2106),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2115),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2122),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2124),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2085),
.B(n_1952),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2133),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_2287),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2138),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2262),
.B(n_1911),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2141),
.Y(n_2543)
);

INVx4_ASAP7_75t_L g2544 ( 
.A(n_2314),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2158),
.Y(n_2545)
);

OR2x6_ASAP7_75t_L g2546 ( 
.A(n_2256),
.B(n_1746),
.Y(n_2546)
);

INVx6_ASAP7_75t_L g2547 ( 
.A(n_2194),
.Y(n_2547)
);

AND2x4_ASAP7_75t_L g2548 ( 
.A(n_2252),
.B(n_2004),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2166),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2316),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2312),
.B(n_1953),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2232),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2314),
.Y(n_2553)
);

CKINVDCx16_ASAP7_75t_R g2554 ( 
.A(n_2207),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2264),
.B(n_1911),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2302),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2316),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2311),
.B(n_2005),
.Y(n_2558)
);

OAI22xp33_ASAP7_75t_L g2559 ( 
.A1(n_2265),
.A2(n_1965),
.B1(n_1991),
.B2(n_1937),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_2317),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2151),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2183),
.B(n_2005),
.Y(n_2562)
);

INVx2_ASAP7_75t_SL g2563 ( 
.A(n_2263),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2320),
.Y(n_2564)
);

OR2x6_ASAP7_75t_L g2565 ( 
.A(n_2265),
.B(n_1965),
.Y(n_2565)
);

INVx4_ASAP7_75t_L g2566 ( 
.A(n_2303),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2177),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2320),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_L g2569 ( 
.A(n_2218),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2082),
.Y(n_2570)
);

NAND2xp33_ASAP7_75t_SL g2571 ( 
.A(n_2301),
.B(n_1965),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2100),
.B(n_1991),
.Y(n_2572)
);

BUFx6f_ASAP7_75t_L g2573 ( 
.A(n_2300),
.Y(n_2573)
);

OA22x2_ASAP7_75t_L g2574 ( 
.A1(n_2290),
.A2(n_1994),
.B1(n_1907),
.B2(n_1931),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2297),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2298),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2205),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2210),
.Y(n_2578)
);

INVxp67_ASAP7_75t_SL g2579 ( 
.A(n_2102),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2313),
.A2(n_1782),
.B1(n_1931),
.B2(n_1878),
.Y(n_2580)
);

INVx1_ASAP7_75t_SL g2581 ( 
.A(n_2228),
.Y(n_2581)
);

BUFx3_ASAP7_75t_L g2582 ( 
.A(n_2185),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2010),
.B(n_1991),
.Y(n_2583)
);

AOI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2014),
.A2(n_1861),
.B1(n_1866),
.B2(n_1859),
.Y(n_2584)
);

BUFx6f_ASAP7_75t_L g2585 ( 
.A(n_2303),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2190),
.B(n_1937),
.Y(n_2586)
);

NAND3xp33_ASAP7_75t_L g2587 ( 
.A(n_2039),
.B(n_1991),
.C(n_1926),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2105),
.Y(n_2588)
);

OR2x2_ASAP7_75t_L g2589 ( 
.A(n_2197),
.B(n_1971),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2082),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_2018),
.B(n_1926),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2150),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_SL g2593 ( 
.A(n_2029),
.B(n_1926),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2030),
.B(n_1896),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2149),
.B(n_1994),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2187),
.B(n_1896),
.Y(n_2596)
);

BUFx6f_ASAP7_75t_L g2597 ( 
.A(n_2273),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2090),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2152),
.Y(n_2599)
);

AND2x2_ASAP7_75t_SL g2600 ( 
.A(n_2327),
.B(n_1859),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2176),
.B(n_1896),
.Y(n_2601)
);

OR2x2_ASAP7_75t_L g2602 ( 
.A(n_2204),
.B(n_1896),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2080),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2090),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2099),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2209),
.B(n_1896),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2099),
.Y(n_2607)
);

BUFx3_ASAP7_75t_L g2608 ( 
.A(n_2226),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2080),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2149),
.B(n_1826),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_2052),
.B(n_1833),
.Y(n_2611)
);

INVxp33_ASAP7_75t_L g2612 ( 
.A(n_2143),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2021),
.B(n_2022),
.Y(n_2613)
);

BUFx8_ASAP7_75t_SL g2614 ( 
.A(n_2046),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2289),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2180),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2304),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2324),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2227),
.Y(n_2619)
);

AOI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2321),
.A2(n_1850),
.B1(n_1883),
.B2(n_1878),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2037),
.B(n_1859),
.Y(n_2621)
);

AOI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2047),
.A2(n_1861),
.B1(n_1866),
.B2(n_1859),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2160),
.Y(n_2623)
);

NOR3xp33_ASAP7_75t_L g2624 ( 
.A(n_2213),
.B(n_1885),
.C(n_1883),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2118),
.Y(n_2625)
);

INVx2_ASAP7_75t_SL g2626 ( 
.A(n_2167),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2199),
.B(n_1859),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2113),
.Y(n_2628)
);

NAND2xp33_ASAP7_75t_L g2629 ( 
.A(n_2215),
.B(n_1879),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2248),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2060),
.B(n_1833),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2078),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2054),
.B(n_1861),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2230),
.B(n_1861),
.Y(n_2634)
);

BUFx10_ASAP7_75t_L g2635 ( 
.A(n_2161),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_2173),
.Y(n_2636)
);

INVx4_ASAP7_75t_L g2637 ( 
.A(n_2078),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2064),
.B(n_1861),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2035),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2038),
.B(n_1833),
.Y(n_2640)
);

AND3x2_ASAP7_75t_L g2641 ( 
.A(n_2308),
.B(n_2235),
.C(n_2248),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2169),
.B(n_1833),
.Y(n_2642)
);

AND2x6_ASAP7_75t_L g2643 ( 
.A(n_2246),
.B(n_1800),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2147),
.Y(n_2644)
);

NOR2x1p5_ASAP7_75t_L g2645 ( 
.A(n_2088),
.B(n_1950),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2153),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2039),
.B(n_1866),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2322),
.A2(n_1883),
.B1(n_1885),
.B2(n_1878),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2114),
.Y(n_2649)
);

BUFx10_ASAP7_75t_L g2650 ( 
.A(n_2161),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2168),
.B(n_1899),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2260),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2162),
.B(n_2165),
.Y(n_2653)
);

BUFx10_ASAP7_75t_L g2654 ( 
.A(n_2012),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2091),
.B(n_1915),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2130),
.B(n_1866),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2179),
.B(n_1899),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2260),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2306),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2134),
.B(n_1866),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2110),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2288),
.A2(n_1869),
.B1(n_1900),
.B2(n_1899),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2087),
.B(n_1869),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2076),
.B(n_1869),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2307),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2110),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2095),
.Y(n_2667)
);

INVx3_ASAP7_75t_L g2668 ( 
.A(n_2119),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2126),
.B(n_1869),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2182),
.B(n_2026),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2299),
.A2(n_2305),
.B1(n_2318),
.B2(n_2315),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2119),
.Y(n_2672)
);

INVx4_ASAP7_75t_L g2673 ( 
.A(n_2307),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2137),
.B(n_1869),
.Y(n_2674)
);

AND2x2_ASAP7_75t_SL g2675 ( 
.A(n_2247),
.B(n_1899),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2094),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2139),
.B(n_1899),
.Y(n_2677)
);

NAND2xp33_ASAP7_75t_SL g2678 ( 
.A(n_2323),
.B(n_1800),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2251),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2144),
.B(n_1900),
.Y(n_2680)
);

INVx4_ASAP7_75t_L g2681 ( 
.A(n_2026),
.Y(n_2681)
);

BUFx10_ASAP7_75t_L g2682 ( 
.A(n_2043),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2342),
.B(n_2043),
.Y(n_2683)
);

NAND2xp33_ASAP7_75t_L g2684 ( 
.A(n_2465),
.B(n_1879),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2437),
.Y(n_2685)
);

AND2x4_ASAP7_75t_L g2686 ( 
.A(n_2454),
.B(n_1879),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2338),
.Y(n_2687)
);

NAND3xp33_ASAP7_75t_L g2688 ( 
.A(n_2334),
.B(n_2277),
.C(n_2268),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2338),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2454),
.B(n_1879),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2349),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2516),
.B(n_2582),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2349),
.Y(n_2693)
);

INVx3_ASAP7_75t_L g2694 ( 
.A(n_2352),
.Y(n_2694)
);

AND2x6_ASAP7_75t_L g2695 ( 
.A(n_2434),
.B(n_2278),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2359),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2408),
.B(n_2159),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2362),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2335),
.Y(n_2699)
);

OAI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2378),
.A2(n_2293),
.B1(n_2280),
.B2(n_2257),
.Y(n_2700)
);

INVx5_ASAP7_75t_L g2701 ( 
.A(n_2465),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2552),
.B(n_2556),
.Y(n_2702)
);

BUFx6f_ASAP7_75t_L g2703 ( 
.A(n_2362),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2359),
.Y(n_2704)
);

BUFx6f_ASAP7_75t_L g2705 ( 
.A(n_2352),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2369),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2369),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2379),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2379),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2380),
.Y(n_2710)
);

AND2x4_ASAP7_75t_L g2711 ( 
.A(n_2582),
.B(n_1885),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2380),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2470),
.B(n_2084),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_2412),
.B(n_1940),
.Y(n_2714)
);

BUFx6f_ASAP7_75t_L g2715 ( 
.A(n_2352),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2352),
.Y(n_2716)
);

AND2x4_ASAP7_75t_L g2717 ( 
.A(n_2441),
.B(n_1915),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2384),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2384),
.Y(n_2719)
);

OR2x2_ASAP7_75t_SL g2720 ( 
.A(n_2554),
.B(n_2017),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2334),
.B(n_1794),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_L g2722 ( 
.A(n_2470),
.B(n_2093),
.Y(n_2722)
);

NAND2x1p5_ASAP7_75t_L g2723 ( 
.A(n_2355),
.B(n_1855),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2385),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_2355),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2479),
.B(n_1915),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2385),
.Y(n_2727)
);

OAI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2378),
.A2(n_2478),
.B1(n_2430),
.B2(n_2526),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2397),
.Y(n_2729)
);

INVx2_ASAP7_75t_SL g2730 ( 
.A(n_2339),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2397),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2398),
.Y(n_2732)
);

NAND2xp33_ASAP7_75t_L g2733 ( 
.A(n_2465),
.B(n_1900),
.Y(n_2733)
);

INVx4_ASAP7_75t_SL g2734 ( 
.A(n_2367),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2553),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2420),
.B(n_1794),
.Y(n_2736)
);

INVx5_ASAP7_75t_L g2737 ( 
.A(n_2465),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2478),
.A2(n_2296),
.B1(n_2266),
.B2(n_2267),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2398),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2355),
.Y(n_2740)
);

NAND2x1p5_ASAP7_75t_L g2741 ( 
.A(n_2355),
.B(n_1855),
.Y(n_2741)
);

AO21x2_ASAP7_75t_L g2742 ( 
.A1(n_2343),
.A2(n_2353),
.B(n_2329),
.Y(n_2742)
);

NAND2x1p5_ASAP7_75t_L g2743 ( 
.A(n_2370),
.B(n_1799),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2553),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2420),
.B(n_1794),
.Y(n_2745)
);

AND2x4_ASAP7_75t_L g2746 ( 
.A(n_2498),
.B(n_1770),
.Y(n_2746)
);

NAND3xp33_ASAP7_75t_L g2747 ( 
.A(n_2484),
.B(n_2109),
.C(n_2294),
.Y(n_2747)
);

AND2x4_ASAP7_75t_L g2748 ( 
.A(n_2429),
.B(n_1770),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_L g2749 ( 
.A(n_2396),
.B(n_2254),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2404),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2332),
.B(n_2017),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2333),
.B(n_1904),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2462),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_2335),
.Y(n_2754)
);

AND2x6_ASAP7_75t_L g2755 ( 
.A(n_2550),
.B(n_1800),
.Y(n_2755)
);

NAND2x1p5_ASAP7_75t_L g2756 ( 
.A(n_2370),
.B(n_1799),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2404),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2421),
.B(n_1800),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2406),
.Y(n_2759)
);

INVx1_ASAP7_75t_SL g2760 ( 
.A(n_2386),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2484),
.B(n_1785),
.Y(n_2761)
);

INVx4_ASAP7_75t_L g2762 ( 
.A(n_2370),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2406),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2524),
.Y(n_2764)
);

AND2x4_ASAP7_75t_L g2765 ( 
.A(n_2429),
.B(n_1785),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2524),
.Y(n_2766)
);

NAND3xp33_ASAP7_75t_L g2767 ( 
.A(n_2412),
.B(n_2337),
.C(n_2501),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2421),
.B(n_1800),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2348),
.Y(n_2769)
);

AOI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2389),
.A2(n_2223),
.B1(n_2259),
.B2(n_2193),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2354),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2423),
.B(n_1809),
.Y(n_2772)
);

NAND2x1p5_ASAP7_75t_L g2773 ( 
.A(n_2370),
.B(n_1727),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2356),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2357),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2396),
.B(n_1900),
.Y(n_2776)
);

INVx2_ASAP7_75t_SL g2777 ( 
.A(n_2375),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2361),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2448),
.Y(n_2779)
);

BUFx3_ASAP7_75t_L g2780 ( 
.A(n_2547),
.Y(n_2780)
);

AND2x4_ASAP7_75t_L g2781 ( 
.A(n_2616),
.B(n_1900),
.Y(n_2781)
);

BUFx3_ASAP7_75t_L g2782 ( 
.A(n_2547),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2626),
.B(n_1902),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2368),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2442),
.Y(n_2785)
);

INVx4_ASAP7_75t_L g2786 ( 
.A(n_2374),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2443),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2456),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2350),
.Y(n_2789)
);

INVx6_ASAP7_75t_L g2790 ( 
.A(n_2426),
.Y(n_2790)
);

CKINVDCx16_ASAP7_75t_R g2791 ( 
.A(n_2448),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2544),
.Y(n_2792)
);

BUFx3_ASAP7_75t_L g2793 ( 
.A(n_2547),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_2612),
.B(n_2261),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2529),
.Y(n_2795)
);

BUFx2_ASAP7_75t_L g2796 ( 
.A(n_2577),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2496),
.B(n_1902),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2423),
.B(n_1809),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2464),
.Y(n_2799)
);

AND2x4_ASAP7_75t_L g2800 ( 
.A(n_2483),
.B(n_1902),
.Y(n_2800)
);

AND2x6_ASAP7_75t_L g2801 ( 
.A(n_2550),
.B(n_1809),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2468),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2601),
.B(n_1902),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2424),
.B(n_1809),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_L g2805 ( 
.A(n_2350),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_2394),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2371),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2475),
.Y(n_2808)
);

AO22x2_ASAP7_75t_L g2809 ( 
.A1(n_2673),
.A2(n_2274),
.B1(n_2284),
.B2(n_2269),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2337),
.B(n_1940),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2476),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2477),
.Y(n_2812)
);

AOI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2389),
.A2(n_2286),
.B1(n_2309),
.B2(n_1902),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2374),
.Y(n_2814)
);

OR2x2_ASAP7_75t_SL g2815 ( 
.A(n_2407),
.B(n_1940),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2485),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2529),
.Y(n_2817)
);

AND2x6_ASAP7_75t_L g2818 ( 
.A(n_2557),
.B(n_1809),
.Y(n_2818)
);

INVx4_ASAP7_75t_L g2819 ( 
.A(n_2374),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2381),
.B(n_1870),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2340),
.Y(n_2821)
);

INVx3_ASAP7_75t_L g2822 ( 
.A(n_2400),
.Y(n_2822)
);

INVx2_ASAP7_75t_SL g2823 ( 
.A(n_2597),
.Y(n_2823)
);

BUFx3_ASAP7_75t_L g2824 ( 
.A(n_2446),
.Y(n_2824)
);

INVxp67_ASAP7_75t_SL g2825 ( 
.A(n_2424),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2405),
.B(n_1727),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2615),
.B(n_1884),
.Y(n_2827)
);

INVx2_ASAP7_75t_SL g2828 ( 
.A(n_2597),
.Y(n_2828)
);

NOR2xp33_ASAP7_75t_L g2829 ( 
.A(n_2612),
.B(n_1950),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2489),
.Y(n_2830)
);

OAI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2574),
.A2(n_1893),
.B1(n_1815),
.B2(n_1816),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2371),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2450),
.B(n_2466),
.Y(n_2833)
);

AND2x4_ASAP7_75t_L g2834 ( 
.A(n_2405),
.B(n_1727),
.Y(n_2834)
);

AOI22xp5_ASAP7_75t_L g2835 ( 
.A1(n_2671),
.A2(n_1815),
.B1(n_1816),
.B2(n_1791),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2597),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2490),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2491),
.Y(n_2838)
);

INVx2_ASAP7_75t_SL g2839 ( 
.A(n_2597),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2414),
.Y(n_2840)
);

AO22x1_ASAP7_75t_L g2841 ( 
.A1(n_2636),
.A2(n_1950),
.B1(n_54),
.B2(n_52),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2530),
.Y(n_2842)
);

AO22x2_ASAP7_75t_L g2843 ( 
.A1(n_2673),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2530),
.Y(n_2844)
);

OAI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2430),
.A2(n_1848),
.B1(n_1815),
.B2(n_1816),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2409),
.Y(n_2846)
);

INVxp67_ASAP7_75t_L g2847 ( 
.A(n_2623),
.Y(n_2847)
);

INVx4_ASAP7_75t_L g2848 ( 
.A(n_2416),
.Y(n_2848)
);

OR2x2_ASAP7_75t_L g2849 ( 
.A(n_2581),
.B(n_1791),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2432),
.B(n_1848),
.Y(n_2850)
);

INVx4_ASAP7_75t_L g2851 ( 
.A(n_2416),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_L g2852 ( 
.A(n_2532),
.B(n_1791),
.Y(n_2852)
);

INVx3_ASAP7_75t_R g2853 ( 
.A(n_2586),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2427),
.B(n_1791),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2409),
.Y(n_2855)
);

AO22x2_ASAP7_75t_L g2856 ( 
.A1(n_2630),
.A2(n_2658),
.B1(n_2665),
.B2(n_2652),
.Y(n_2856)
);

INVx2_ASAP7_75t_SL g2857 ( 
.A(n_2563),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2419),
.Y(n_2858)
);

OAI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2526),
.A2(n_2431),
.B1(n_2580),
.B2(n_2570),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2422),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2371),
.Y(n_2861)
);

INVx4_ASAP7_75t_L g2862 ( 
.A(n_2427),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2425),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2506),
.B(n_1815),
.Y(n_2864)
);

BUFx2_ASAP7_75t_L g2865 ( 
.A(n_2565),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2341),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_2585),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2433),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2532),
.B(n_1816),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2506),
.B(n_1836),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2435),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2438),
.Y(n_2872)
);

BUFx6f_ASAP7_75t_L g2873 ( 
.A(n_2573),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2573),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2459),
.B(n_1836),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2533),
.Y(n_2876)
);

CKINVDCx20_ASAP7_75t_R g2877 ( 
.A(n_2336),
.Y(n_2877)
);

BUFx6f_ASAP7_75t_L g2878 ( 
.A(n_2573),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2544),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2439),
.Y(n_2880)
);

AND2x4_ASAP7_75t_L g2881 ( 
.A(n_2517),
.B(n_1836),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2432),
.B(n_1848),
.Y(n_2882)
);

NAND2x1p5_ASAP7_75t_L g2883 ( 
.A(n_2347),
.B(n_1836),
.Y(n_2883)
);

BUFx4f_ASAP7_75t_L g2884 ( 
.A(n_2409),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2517),
.B(n_2502),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2533),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2534),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2501),
.B(n_1848),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2455),
.Y(n_2889)
);

CKINVDCx20_ASAP7_75t_R g2890 ( 
.A(n_2639),
.Y(n_2890)
);

BUFx3_ASAP7_75t_L g2891 ( 
.A(n_2461),
.Y(n_2891)
);

NAND3xp33_ASAP7_75t_L g2892 ( 
.A(n_2459),
.B(n_1848),
.C(n_1786),
.Y(n_2892)
);

AO22x2_ASAP7_75t_L g2893 ( 
.A1(n_2630),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2400),
.B(n_1784),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2328),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2344),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2346),
.Y(n_2897)
);

INVx4_ASAP7_75t_L g2898 ( 
.A(n_2347),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2447),
.Y(n_2899)
);

INVx4_ASAP7_75t_L g2900 ( 
.A(n_2392),
.Y(n_2900)
);

BUFx3_ASAP7_75t_L g2901 ( 
.A(n_2461),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2681),
.B(n_1784),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2567),
.B(n_1784),
.Y(n_2903)
);

INVx4_ASAP7_75t_L g2904 ( 
.A(n_2392),
.Y(n_2904)
);

AND2x4_ASAP7_75t_L g2905 ( 
.A(n_2625),
.B(n_1784),
.Y(n_2905)
);

CKINVDCx14_ASAP7_75t_R g2906 ( 
.A(n_2461),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2447),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2473),
.B(n_703),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2534),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2452),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2452),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2463),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2463),
.B(n_1784),
.Y(n_2913)
);

INVx1_ASAP7_75t_SL g2914 ( 
.A(n_2655),
.Y(n_2914)
);

HB1xp67_ASAP7_75t_L g2915 ( 
.A(n_2604),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2474),
.Y(n_2916)
);

AOI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2329),
.A2(n_1788),
.B1(n_1786),
.B2(n_1753),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2536),
.Y(n_2918)
);

INVx4_ASAP7_75t_L g2919 ( 
.A(n_2351),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2474),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_2625),
.B(n_1786),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2536),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2585),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2488),
.Y(n_2924)
);

INVx1_ASAP7_75t_SL g2925 ( 
.A(n_2678),
.Y(n_2925)
);

AOI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2345),
.A2(n_1788),
.B1(n_1786),
.B2(n_1753),
.Y(n_2926)
);

BUFx3_ASAP7_75t_L g2927 ( 
.A(n_2480),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2537),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2436),
.B(n_1786),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2537),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2488),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2499),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2499),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2511),
.Y(n_2934)
);

NOR2xp33_ASAP7_75t_L g2935 ( 
.A(n_2538),
.B(n_1788),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2539),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2511),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_SL g2938 ( 
.A(n_2559),
.B(n_2431),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2539),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2480),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2473),
.B(n_703),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2543),
.Y(n_2942)
);

AND2x2_ASAP7_75t_SL g2943 ( 
.A(n_2675),
.B(n_2351),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2543),
.Y(n_2944)
);

AND2x4_ASAP7_75t_L g2945 ( 
.A(n_2363),
.B(n_1788),
.Y(n_2945)
);

INVxp67_ASAP7_75t_L g2946 ( 
.A(n_2575),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2681),
.B(n_1788),
.Y(n_2947)
);

BUFx3_ASAP7_75t_L g2948 ( 
.A(n_2480),
.Y(n_2948)
);

BUFx3_ASAP7_75t_L g2949 ( 
.A(n_2453),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_2520),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2545),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2545),
.Y(n_2952)
);

AO22x2_ASAP7_75t_L g2953 ( 
.A1(n_2652),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2549),
.Y(n_2954)
);

CKINVDCx5p33_ASAP7_75t_R g2955 ( 
.A(n_2520),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2667),
.B(n_170),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_L g2957 ( 
.A(n_2573),
.Y(n_2957)
);

BUFx3_ASAP7_75t_L g2958 ( 
.A(n_2453),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2576),
.B(n_1753),
.Y(n_2959)
);

AND2x6_ASAP7_75t_L g2960 ( 
.A(n_2557),
.B(n_1753),
.Y(n_2960)
);

OR2x6_ASAP7_75t_L g2961 ( 
.A(n_2565),
.B(n_1753),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2549),
.Y(n_2962)
);

BUFx12f_ASAP7_75t_L g2963 ( 
.A(n_2635),
.Y(n_2963)
);

INVx3_ASAP7_75t_L g2964 ( 
.A(n_2515),
.Y(n_2964)
);

BUFx10_ASAP7_75t_L g2965 ( 
.A(n_2572),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2515),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2387),
.B(n_1796),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2460),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2564),
.Y(n_2969)
);

AND2x4_ASAP7_75t_L g2970 ( 
.A(n_2391),
.B(n_1796),
.Y(n_2970)
);

INVx3_ASAP7_75t_L g2971 ( 
.A(n_2515),
.Y(n_2971)
);

INVx4_ASAP7_75t_L g2972 ( 
.A(n_2367),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2667),
.B(n_56),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2527),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2527),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_2914),
.B(n_2559),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2753),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2702),
.B(n_2679),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2914),
.B(n_2670),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2687),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2713),
.B(n_2572),
.Y(n_2981)
);

HB1xp67_ASAP7_75t_L g2982 ( 
.A(n_2753),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2702),
.B(n_2366),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2946),
.B(n_2925),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2946),
.B(n_2538),
.Y(n_2985)
);

NOR3xp33_ASAP7_75t_L g2986 ( 
.A(n_2688),
.B(n_2747),
.C(n_2471),
.Y(n_2986)
);

OAI22xp33_ASAP7_75t_SL g2987 ( 
.A1(n_2938),
.A2(n_2700),
.B1(n_2613),
.B2(n_2973),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2704),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2925),
.B(n_2659),
.Y(n_2989)
);

INVxp67_ASAP7_75t_L g2990 ( 
.A(n_2833),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2856),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2856),
.Y(n_2992)
);

INVx3_ASAP7_75t_L g2993 ( 
.A(n_2966),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2968),
.B(n_2659),
.Y(n_2994)
);

OR2x6_ASAP7_75t_L g2995 ( 
.A(n_2961),
.B(n_2453),
.Y(n_2995)
);

AND2x6_ASAP7_75t_SL g2996 ( 
.A(n_2749),
.B(n_2546),
.Y(n_2996)
);

AOI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2733),
.A2(n_2372),
.B(n_2507),
.Y(n_2997)
);

INVxp67_ASAP7_75t_L g2998 ( 
.A(n_2796),
.Y(n_2998)
);

NOR2xp33_ASAP7_75t_L g2999 ( 
.A(n_2713),
.B(n_2589),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_2791),
.B(n_2585),
.Y(n_3000)
);

INVxp67_ASAP7_75t_L g3001 ( 
.A(n_2760),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2827),
.B(n_2825),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2760),
.B(n_2722),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2709),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2825),
.B(n_2659),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2779),
.B(n_2585),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2767),
.B(n_2659),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2722),
.B(n_2410),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2683),
.B(n_2676),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2688),
.A2(n_2574),
.B1(n_2613),
.B2(n_2608),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2712),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2915),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2767),
.B(n_2642),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2915),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_2747),
.A2(n_2608),
.B1(n_2619),
.B2(n_2653),
.Y(n_3015)
);

OR2x2_ASAP7_75t_L g3016 ( 
.A(n_2777),
.B(n_2602),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2776),
.B(n_2642),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2794),
.B(n_2640),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2794),
.B(n_2640),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2692),
.B(n_2358),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2735),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2735),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2692),
.B(n_2570),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2718),
.Y(n_3024)
);

NAND2x1p5_ASAP7_75t_L g3025 ( 
.A(n_2701),
.B(n_2737),
.Y(n_3025)
);

AOI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2749),
.A2(n_2571),
.B1(n_2631),
.B2(n_2611),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2698),
.B(n_2566),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2726),
.B(n_2590),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2847),
.B(n_2410),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2684),
.A2(n_2372),
.B(n_2393),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2744),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2726),
.B(n_2590),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2820),
.B(n_2598),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2744),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_SL g3035 ( 
.A(n_2698),
.B(n_2703),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2724),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2847),
.B(n_2493),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2770),
.B(n_2598),
.Y(n_3038)
);

INVx4_ASAP7_75t_L g3039 ( 
.A(n_2698),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2785),
.Y(n_3040)
);

O2A1O1Ixp33_ASAP7_75t_L g3041 ( 
.A1(n_2700),
.A2(n_2353),
.B(n_2345),
.C(n_2583),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2770),
.B(n_2605),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2810),
.B(n_2493),
.Y(n_3043)
);

INVx3_ASAP7_75t_L g3044 ( 
.A(n_2966),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2738),
.A2(n_2619),
.B1(n_2617),
.B2(n_2618),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2717),
.B(n_2852),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2717),
.B(n_2605),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2852),
.B(n_2607),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2869),
.B(n_2607),
.Y(n_3049)
);

NAND2x1p5_ASAP7_75t_L g3050 ( 
.A(n_2701),
.B(n_2364),
.Y(n_3050)
);

AOI221xp5_ASAP7_75t_L g3051 ( 
.A1(n_2973),
.A2(n_2672),
.B1(n_2678),
.B2(n_2510),
.C(n_2603),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2966),
.Y(n_3052)
);

OAI22xp5_ASAP7_75t_L g3053 ( 
.A1(n_2943),
.A2(n_2482),
.B1(n_2631),
.B2(n_2611),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2729),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2703),
.B(n_2566),
.Y(n_3055)
);

AO22x1_ASAP7_75t_L g3056 ( 
.A1(n_2950),
.A2(n_2578),
.B1(n_2469),
.B2(n_2596),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2787),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2788),
.Y(n_3058)
);

AND2x6_ASAP7_75t_SL g3059 ( 
.A(n_2829),
.B(n_2546),
.Y(n_3059)
);

OR2x2_ASAP7_75t_L g3060 ( 
.A(n_2752),
.B(n_2730),
.Y(n_3060)
);

A2O1A1Ixp33_ASAP7_75t_SL g3061 ( 
.A1(n_2935),
.A2(n_2596),
.B(n_2651),
.C(n_2657),
.Y(n_3061)
);

BUFx8_ASAP7_75t_L g3062 ( 
.A(n_2963),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2869),
.B(n_2609),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_2738),
.A2(n_2617),
.B1(n_2618),
.B2(n_2675),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2689),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2799),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2888),
.B(n_2609),
.Y(n_3067)
);

NOR3xp33_ASAP7_75t_L g3068 ( 
.A(n_2714),
.B(n_2587),
.C(n_2571),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2691),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2693),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_2853),
.B(n_2606),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2802),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2965),
.B(n_2646),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2965),
.B(n_2637),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2703),
.B(n_2515),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2888),
.B(n_2604),
.Y(n_3076)
);

NAND3xp33_ASAP7_75t_SL g3077 ( 
.A(n_2813),
.B(n_2624),
.C(n_2449),
.Y(n_3077)
);

OAI22xp5_ASAP7_75t_L g3078 ( 
.A1(n_2859),
.A2(n_2728),
.B1(n_2482),
.B2(n_2651),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2829),
.A2(n_2583),
.B1(n_2565),
.B2(n_2418),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2823),
.B(n_2644),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2828),
.B(n_2836),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2808),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2839),
.B(n_2665),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2789),
.B(n_2540),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2696),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_2695),
.A2(n_2658),
.B1(n_2600),
.B2(n_2668),
.Y(n_3086)
);

INVxp67_ASAP7_75t_SL g3087 ( 
.A(n_2845),
.Y(n_3087)
);

AND3x1_ASAP7_75t_L g3088 ( 
.A(n_2751),
.B(n_2668),
.C(n_2632),
.Y(n_3088)
);

O2A1O1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_2697),
.A2(n_2418),
.B(n_2562),
.C(n_2661),
.Y(n_3089)
);

CKINVDCx5p33_ASAP7_75t_R g3090 ( 
.A(n_2806),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2956),
.B(n_2676),
.Y(n_3091)
);

O2A1O1Ixp33_ASAP7_75t_L g3092 ( 
.A1(n_2859),
.A2(n_2666),
.B(n_2610),
.C(n_2669),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2789),
.B(n_2540),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2809),
.B(n_2657),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2809),
.B(n_2811),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2792),
.B(n_2637),
.Y(n_3096)
);

AND3x2_ASAP7_75t_L g3097 ( 
.A(n_2908),
.B(n_2548),
.C(n_2558),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2812),
.B(n_2444),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2706),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_2890),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2707),
.Y(n_3101)
);

AO22x1_ASAP7_75t_L g3102 ( 
.A1(n_2955),
.A2(n_2509),
.B1(n_2548),
.B2(n_2632),
.Y(n_3102)
);

INVxp67_ASAP7_75t_L g3103 ( 
.A(n_2849),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2816),
.B(n_2540),
.Y(n_3104)
);

HB1xp67_ASAP7_75t_L g3105 ( 
.A(n_2792),
.Y(n_3105)
);

INVx1_ASAP7_75t_SL g3106 ( 
.A(n_2821),
.Y(n_3106)
);

NAND2xp33_ASAP7_75t_L g3107 ( 
.A(n_2873),
.B(n_2367),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2789),
.B(n_2540),
.Y(n_3108)
);

OAI21xp33_ASAP7_75t_L g3109 ( 
.A1(n_2813),
.A2(n_2664),
.B(n_2504),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2830),
.B(n_2837),
.Y(n_3110)
);

INVxp67_ASAP7_75t_SL g3111 ( 
.A(n_2845),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2805),
.B(n_2482),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2708),
.Y(n_3113)
);

INVx2_ASAP7_75t_SL g3114 ( 
.A(n_2805),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2838),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_2877),
.B(n_2857),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2805),
.B(n_2482),
.Y(n_3117)
);

AND2x2_ASAP7_75t_SL g3118 ( 
.A(n_2941),
.B(n_2600),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2867),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2710),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2840),
.B(n_2519),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2858),
.B(n_2519),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2860),
.B(n_2487),
.Y(n_3123)
);

NOR2x2_ASAP7_75t_L g3124 ( 
.A(n_2961),
.B(n_2546),
.Y(n_3124)
);

INVx2_ASAP7_75t_SL g3125 ( 
.A(n_2923),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2863),
.B(n_2504),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2719),
.Y(n_3127)
);

OR2x6_ASAP7_75t_L g3128 ( 
.A(n_2961),
.B(n_2645),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2868),
.B(n_2871),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2872),
.B(n_2592),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2711),
.B(n_2558),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2879),
.Y(n_3132)
);

INVx2_ASAP7_75t_SL g3133 ( 
.A(n_2846),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_2780),
.B(n_2428),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2880),
.B(n_2599),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2695),
.B(n_2548),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2727),
.Y(n_3137)
);

OR2x2_ASAP7_75t_L g3138 ( 
.A(n_2782),
.B(n_2494),
.Y(n_3138)
);

BUFx8_ASAP7_75t_L g3139 ( 
.A(n_2865),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_L g3140 ( 
.A(n_2793),
.B(n_2428),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2695),
.B(n_2560),
.Y(n_3141)
);

NAND2x1p5_ASAP7_75t_L g3142 ( 
.A(n_2701),
.B(n_2364),
.Y(n_3142)
);

INVx2_ASAP7_75t_SL g3143 ( 
.A(n_2855),
.Y(n_3143)
);

INVx2_ASAP7_75t_SL g3144 ( 
.A(n_2891),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2731),
.Y(n_3145)
);

AOI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2695),
.A2(n_2360),
.B1(n_2551),
.B2(n_2525),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2711),
.A2(n_2360),
.B1(n_2551),
.B2(n_2525),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2721),
.B(n_2560),
.Y(n_3148)
);

AND2x4_ASAP7_75t_L g3149 ( 
.A(n_2885),
.B(n_2401),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2721),
.B(n_2560),
.Y(n_3150)
);

INVx4_ASAP7_75t_L g3151 ( 
.A(n_2705),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2895),
.B(n_2560),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2896),
.B(n_2620),
.Y(n_3153)
);

BUFx3_ASAP7_75t_L g3154 ( 
.A(n_2699),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2897),
.B(n_2620),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2964),
.B(n_2648),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2964),
.B(n_2648),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2732),
.Y(n_3158)
);

INVxp67_ASAP7_75t_L g3159 ( 
.A(n_2879),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2949),
.B(n_2682),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2971),
.B(n_2377),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_SL g3162 ( 
.A(n_2885),
.B(n_2558),
.Y(n_3162)
);

OR2x6_ASAP7_75t_L g3163 ( 
.A(n_2754),
.B(n_2376),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2739),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_2866),
.B(n_2682),
.Y(n_3165)
);

BUFx3_ASAP7_75t_L g3166 ( 
.A(n_2685),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2769),
.Y(n_3167)
);

INVx2_ASAP7_75t_SL g3168 ( 
.A(n_2901),
.Y(n_3168)
);

NOR2x1_ASAP7_75t_L g3169 ( 
.A(n_2848),
.B(n_2376),
.Y(n_3169)
);

BUFx6f_ASAP7_75t_L g3170 ( 
.A(n_2705),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2750),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_2843),
.A2(n_2682),
.B1(n_2634),
.B2(n_2677),
.Y(n_3172)
);

NAND2x1_ASAP7_75t_L g3173 ( 
.A(n_2972),
.B(n_2367),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2971),
.B(n_2781),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2781),
.B(n_2579),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2783),
.B(n_2873),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2783),
.B(n_2580),
.Y(n_3177)
);

AOI221xp5_ASAP7_75t_L g3178 ( 
.A1(n_2843),
.A2(n_2680),
.B1(n_2677),
.B2(n_2674),
.C(n_2638),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_SL g3179 ( 
.A(n_2873),
.B(n_2662),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2874),
.B(n_2402),
.Y(n_3180)
);

AOI21x1_ASAP7_75t_L g3181 ( 
.A1(n_2875),
.A2(n_2331),
.B(n_2621),
.Y(n_3181)
);

AOI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_2803),
.A2(n_2388),
.B1(n_2663),
.B2(n_2797),
.Y(n_3182)
);

AND2x6_ASAP7_75t_SL g3183 ( 
.A(n_2929),
.B(n_2614),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_2958),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2874),
.B(n_2654),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_SL g3186 ( 
.A(n_2874),
.B(n_2654),
.Y(n_3186)
);

AOI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2803),
.A2(n_2388),
.B1(n_2663),
.B2(n_2634),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_SL g3188 ( 
.A(n_2878),
.B(n_2584),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2878),
.B(n_2403),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2771),
.Y(n_3190)
);

AOI22xp33_ASAP7_75t_L g3191 ( 
.A1(n_2893),
.A2(n_2674),
.B1(n_2680),
.B2(n_2595),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2878),
.B(n_2957),
.Y(n_3192)
);

OAI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_2728),
.A2(n_2737),
.B1(n_2503),
.B2(n_2555),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2757),
.Y(n_3194)
);

AND2x4_ASAP7_75t_L g3195 ( 
.A(n_2929),
.B(n_2411),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2774),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2957),
.B(n_2775),
.Y(n_3197)
);

BUFx8_ASAP7_75t_L g3198 ( 
.A(n_2824),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2778),
.Y(n_3199)
);

NOR2x1p5_ASAP7_75t_L g3200 ( 
.A(n_3018),
.B(n_2919),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_3025),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_3003),
.B(n_2884),
.Y(n_3202)
);

AO21x2_ASAP7_75t_L g3203 ( 
.A1(n_2986),
.A2(n_2831),
.B(n_2892),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_2995),
.B(n_2957),
.Y(n_3204)
);

INVx3_ASAP7_75t_L g3205 ( 
.A(n_3025),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_3008),
.B(n_2987),
.Y(n_3206)
);

INVx2_ASAP7_75t_SL g3207 ( 
.A(n_3166),
.Y(n_3207)
);

INVx6_ASAP7_75t_L g3208 ( 
.A(n_3139),
.Y(n_3208)
);

INVxp67_ASAP7_75t_L g3209 ( 
.A(n_3060),
.Y(n_3209)
);

AND2x6_ASAP7_75t_L g3210 ( 
.A(n_3146),
.B(n_2807),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_3100),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2983),
.B(n_2641),
.Y(n_3212)
);

AND2x6_ASAP7_75t_L g3213 ( 
.A(n_3147),
.B(n_2807),
.Y(n_3213)
);

BUFx2_ASAP7_75t_L g3214 ( 
.A(n_3001),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3064),
.B(n_2742),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_3039),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3110),
.Y(n_3217)
);

AO22x1_ASAP7_75t_L g3218 ( 
.A1(n_2999),
.A2(n_2919),
.B1(n_2940),
.B2(n_2927),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3129),
.Y(n_3219)
);

BUFx6f_ASAP7_75t_L g3220 ( 
.A(n_3170),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3040),
.Y(n_3221)
);

BUFx2_ASAP7_75t_L g3222 ( 
.A(n_3001),
.Y(n_3222)
);

OR2x2_ASAP7_75t_L g3223 ( 
.A(n_3019),
.B(n_2990),
.Y(n_3223)
);

INVx3_ASAP7_75t_L g3224 ( 
.A(n_3039),
.Y(n_3224)
);

INVxp67_ASAP7_75t_L g3225 ( 
.A(n_2977),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3057),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3058),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3066),
.Y(n_3228)
);

NOR2xp67_ASAP7_75t_L g3229 ( 
.A(n_2978),
.B(n_2985),
.Y(n_3229)
);

BUFx4f_ASAP7_75t_L g3230 ( 
.A(n_3128),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3002),
.B(n_2981),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3170),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2990),
.B(n_2984),
.Y(n_3233)
);

INVx2_ASAP7_75t_SL g3234 ( 
.A(n_3154),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_3139),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_3043),
.B(n_2614),
.Y(n_3236)
);

CKINVDCx11_ASAP7_75t_R g3237 ( 
.A(n_3183),
.Y(n_3237)
);

INVx2_ASAP7_75t_SL g3238 ( 
.A(n_3090),
.Y(n_3238)
);

AOI22xp5_ASAP7_75t_L g3239 ( 
.A1(n_2976),
.A2(n_2669),
.B1(n_2953),
.B2(n_2893),
.Y(n_3239)
);

BUFx6f_ASAP7_75t_L g3240 ( 
.A(n_3170),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3026),
.B(n_2720),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3072),
.Y(n_3242)
);

INVx2_ASAP7_75t_SL g3243 ( 
.A(n_3114),
.Y(n_3243)
);

AOI221xp5_ASAP7_75t_L g3244 ( 
.A1(n_2986),
.A2(n_2841),
.B1(n_2953),
.B2(n_2831),
.C(n_2638),
.Y(n_3244)
);

INVxp67_ASAP7_75t_L g3245 ( 
.A(n_2977),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_3073),
.B(n_2884),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2980),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_2995),
.B(n_2948),
.Y(n_3248)
);

BUFx6f_ASAP7_75t_L g3249 ( 
.A(n_2995),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2988),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3082),
.Y(n_3251)
);

AOI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_3118),
.A2(n_2647),
.B1(n_2903),
.B2(n_2660),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_2982),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3115),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2994),
.B(n_2737),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3167),
.Y(n_3256)
);

INVx6_ASAP7_75t_L g3257 ( 
.A(n_3198),
.Y(n_3257)
);

HB1xp67_ASAP7_75t_L g3258 ( 
.A(n_2982),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2989),
.B(n_2784),
.Y(n_3259)
);

HB1xp67_ASAP7_75t_L g3260 ( 
.A(n_2998),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3190),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3004),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_3195),
.B(n_2814),
.Y(n_3263)
);

NAND2x1p5_ASAP7_75t_L g3264 ( 
.A(n_3035),
.B(n_2848),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_SL g3265 ( 
.A(n_3071),
.B(n_2800),
.Y(n_3265)
);

INVxp67_ASAP7_75t_L g3266 ( 
.A(n_3029),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3011),
.Y(n_3267)
);

BUFx3_ASAP7_75t_L g3268 ( 
.A(n_3198),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3015),
.B(n_2759),
.Y(n_3269)
);

INVxp67_ASAP7_75t_L g3270 ( 
.A(n_3037),
.Y(n_3270)
);

INVx2_ASAP7_75t_SL g3271 ( 
.A(n_3106),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_3015),
.B(n_2763),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_3024),
.Y(n_3273)
);

A2O1A1Ixp33_ASAP7_75t_L g3274 ( 
.A1(n_3041),
.A2(n_2629),
.B(n_2902),
.C(n_2947),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3038),
.B(n_2974),
.Y(n_3275)
);

INVx2_ASAP7_75t_L g3276 ( 
.A(n_3036),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3064),
.B(n_2742),
.Y(n_3277)
);

BUFx2_ASAP7_75t_L g3278 ( 
.A(n_2998),
.Y(n_3278)
);

OAI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_3086),
.A2(n_2972),
.B1(n_2815),
.B2(n_2907),
.Y(n_3279)
);

OR2x6_ASAP7_75t_L g3280 ( 
.A(n_3030),
.B(n_2807),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3196),
.Y(n_3281)
);

INVx5_ASAP7_75t_L g3282 ( 
.A(n_3151),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3045),
.B(n_2899),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3045),
.B(n_2910),
.Y(n_3284)
);

INVx1_ASAP7_75t_SL g3285 ( 
.A(n_2979),
.Y(n_3285)
);

INVxp67_ASAP7_75t_L g3286 ( 
.A(n_3116),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3048),
.B(n_2911),
.Y(n_3287)
);

INVx4_ASAP7_75t_L g3288 ( 
.A(n_3151),
.Y(n_3288)
);

OR2x2_ASAP7_75t_L g3289 ( 
.A(n_3023),
.B(n_3016),
.Y(n_3289)
);

NOR2xp67_ASAP7_75t_L g3290 ( 
.A(n_3007),
.B(n_2822),
.Y(n_3290)
);

NOR2xp67_ASAP7_75t_L g3291 ( 
.A(n_3013),
.B(n_2822),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3049),
.B(n_2912),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_3050),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3118),
.A2(n_2647),
.B1(n_2903),
.B2(n_2591),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_L g3295 ( 
.A(n_3020),
.B(n_2889),
.Y(n_3295)
);

INVx3_ASAP7_75t_L g3296 ( 
.A(n_3050),
.Y(n_3296)
);

INVx4_ASAP7_75t_L g3297 ( 
.A(n_2993),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3042),
.B(n_2975),
.Y(n_3298)
);

BUFx2_ASAP7_75t_L g3299 ( 
.A(n_3091),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_3134),
.B(n_2814),
.Y(n_3300)
);

OR2x2_ASAP7_75t_L g3301 ( 
.A(n_3103),
.B(n_2939),
.Y(n_3301)
);

BUFx6f_ASAP7_75t_L g3302 ( 
.A(n_2993),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3098),
.B(n_2764),
.Y(n_3303)
);

OAI22xp5_ASAP7_75t_SL g3304 ( 
.A1(n_3172),
.A2(n_2906),
.B1(n_2947),
.B2(n_2902),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_SL g3305 ( 
.A(n_3046),
.B(n_2800),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3009),
.B(n_2905),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3199),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3017),
.B(n_2766),
.Y(n_3308)
);

INVxp67_ASAP7_75t_L g3309 ( 
.A(n_3140),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3065),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3130),
.B(n_2795),
.Y(n_3311)
);

AND2x4_ASAP7_75t_L g3312 ( 
.A(n_3195),
.B(n_2864),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3135),
.B(n_3033),
.Y(n_3313)
);

HB1xp67_ASAP7_75t_L g3314 ( 
.A(n_3105),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_3044),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_3079),
.B(n_2797),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3069),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3054),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3070),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3085),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_3133),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_3143),
.Y(n_3322)
);

CKINVDCx5p33_ASAP7_75t_R g3323 ( 
.A(n_3062),
.Y(n_3323)
);

OR2x2_ASAP7_75t_L g3324 ( 
.A(n_3103),
.B(n_2942),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3067),
.B(n_2916),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3051),
.B(n_2817),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_3051),
.B(n_2905),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_3144),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3099),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3123),
.B(n_3005),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_3080),
.B(n_2832),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3101),
.Y(n_3332)
);

AND3x2_ASAP7_75t_SL g3333 ( 
.A(n_3124),
.B(n_2844),
.C(n_2842),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_3077),
.A2(n_2591),
.B1(n_2593),
.B2(n_2594),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3113),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3063),
.B(n_2920),
.Y(n_3336)
);

INVx2_ASAP7_75t_SL g3337 ( 
.A(n_3168),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3076),
.B(n_2924),
.Y(n_3338)
);

BUFx5_ASAP7_75t_L g3339 ( 
.A(n_2991),
.Y(n_3339)
);

AO22x1_ASAP7_75t_L g3340 ( 
.A1(n_3074),
.A2(n_2870),
.B1(n_2881),
.B2(n_2864),
.Y(n_3340)
);

HB1xp67_ASAP7_75t_L g3341 ( 
.A(n_3105),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3120),
.Y(n_3342)
);

INVx1_ASAP7_75t_SL g3343 ( 
.A(n_3132),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3127),
.Y(n_3344)
);

BUFx3_ASAP7_75t_L g3345 ( 
.A(n_3062),
.Y(n_3345)
);

BUFx6f_ASAP7_75t_L g3346 ( 
.A(n_3044),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3028),
.B(n_2876),
.Y(n_3347)
);

INVx4_ASAP7_75t_L g3348 ( 
.A(n_3052),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3032),
.B(n_2886),
.Y(n_3349)
);

AOI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3010),
.A2(n_2417),
.B1(n_2593),
.B2(n_2594),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3137),
.Y(n_3351)
);

AND2x4_ASAP7_75t_L g3352 ( 
.A(n_3160),
.B(n_2870),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3145),
.Y(n_3353)
);

BUFx2_ASAP7_75t_L g3354 ( 
.A(n_3192),
.Y(n_3354)
);

BUFx3_ASAP7_75t_L g3355 ( 
.A(n_3184),
.Y(n_3355)
);

OR2x2_ASAP7_75t_L g3356 ( 
.A(n_3047),
.B(n_2944),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3158),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3164),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3175),
.B(n_2887),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3088),
.B(n_2921),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3138),
.B(n_2921),
.Y(n_3361)
);

BUFx4f_ASAP7_75t_L g3362 ( 
.A(n_3128),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3171),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3194),
.Y(n_3364)
);

A2O1A1Ixp33_ASAP7_75t_L g3365 ( 
.A1(n_3041),
.A2(n_2629),
.B(n_2393),
.C(n_2633),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3152),
.Y(n_3366)
);

INVx3_ASAP7_75t_L g3367 ( 
.A(n_3142),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3010),
.B(n_2931),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3000),
.B(n_2832),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_3053),
.B(n_2832),
.Y(n_3370)
);

AOI22xp33_ASAP7_75t_L g3371 ( 
.A1(n_3077),
.A2(n_2643),
.B1(n_2633),
.B2(n_2621),
.Y(n_3371)
);

INVx2_ASAP7_75t_SL g3372 ( 
.A(n_3119),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3012),
.Y(n_3373)
);

BUFx2_ASAP7_75t_L g3374 ( 
.A(n_3132),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_3056),
.B(n_2861),
.Y(n_3375)
);

INVx5_ASAP7_75t_L g3376 ( 
.A(n_3163),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3086),
.B(n_2932),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3014),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3021),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3022),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_3052),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_3125),
.Y(n_3382)
);

AND2x4_ASAP7_75t_L g3383 ( 
.A(n_3149),
.B(n_3027),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_SL g3384 ( 
.A(n_3078),
.B(n_2367),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_3031),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3094),
.B(n_2909),
.Y(n_3386)
);

AOI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_3178),
.A2(n_2495),
.B1(n_2761),
.B2(n_2627),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3034),
.Y(n_3388)
);

BUFx3_ASAP7_75t_L g3389 ( 
.A(n_3165),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_2992),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3109),
.B(n_2933),
.Y(n_3391)
);

INVxp67_ASAP7_75t_SL g3392 ( 
.A(n_3104),
.Y(n_3392)
);

INVx5_ASAP7_75t_L g3393 ( 
.A(n_3163),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3148),
.B(n_2934),
.Y(n_3394)
);

INVx2_ASAP7_75t_SL g3395 ( 
.A(n_3055),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3095),
.B(n_2881),
.Y(n_3396)
);

INVx2_ASAP7_75t_SL g3397 ( 
.A(n_3006),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3083),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3150),
.B(n_2937),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3197),
.Y(n_3400)
);

INVx3_ASAP7_75t_L g3401 ( 
.A(n_3142),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3161),
.B(n_2918),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3121),
.Y(n_3403)
);

NOR2x1p5_ASAP7_75t_L g3404 ( 
.A(n_3141),
.B(n_2786),
.Y(n_3404)
);

AOI22xp5_ASAP7_75t_L g3405 ( 
.A1(n_3178),
.A2(n_2643),
.B1(n_2382),
.B2(n_2383),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3122),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_3149),
.Y(n_3407)
);

HB1xp67_ASAP7_75t_L g3408 ( 
.A(n_3159),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3087),
.B(n_2969),
.Y(n_3409)
);

BUFx3_ASAP7_75t_L g3410 ( 
.A(n_3176),
.Y(n_3410)
);

BUFx3_ASAP7_75t_L g3411 ( 
.A(n_3163),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3180),
.Y(n_3412)
);

BUFx6f_ASAP7_75t_L g3413 ( 
.A(n_3128),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3390),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3231),
.B(n_3153),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3239),
.A2(n_3172),
.B1(n_3087),
.B2(n_3111),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_3239),
.A2(n_3111),
.B1(n_3191),
.B2(n_3155),
.Y(n_3417)
);

CKINVDCx5p33_ASAP7_75t_R g3418 ( 
.A(n_3211),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_3365),
.A2(n_3030),
.B(n_3061),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_3229),
.B(n_3068),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3330),
.B(n_3185),
.Y(n_3421)
);

OAI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3244),
.A2(n_3191),
.B1(n_3096),
.B2(n_3159),
.Y(n_3422)
);

OAI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_3405),
.A2(n_3096),
.B1(n_3136),
.B2(n_3177),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3204),
.B(n_3186),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3285),
.B(n_3084),
.Y(n_3425)
);

AOI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3274),
.A2(n_2997),
.B(n_3107),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_3371),
.A2(n_2997),
.B(n_3179),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_3229),
.B(n_3068),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3285),
.B(n_3093),
.Y(n_3429)
);

OAI22xp5_ASAP7_75t_L g3430 ( 
.A1(n_3405),
.A2(n_3126),
.B1(n_3157),
.B2(n_3156),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3313),
.B(n_3223),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3233),
.B(n_3102),
.Y(n_3432)
);

AOI21x1_ASAP7_75t_L g3433 ( 
.A1(n_3206),
.A2(n_3181),
.B(n_3188),
.Y(n_3433)
);

NAND2x1p5_ASAP7_75t_L g3434 ( 
.A(n_3376),
.B(n_3169),
.Y(n_3434)
);

O2A1O1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_3202),
.A2(n_3092),
.B(n_3162),
.C(n_3193),
.Y(n_3435)
);

AOI21x1_ASAP7_75t_L g3436 ( 
.A1(n_3218),
.A2(n_2959),
.B(n_3173),
.Y(n_3436)
);

AOI22x1_ASAP7_75t_L g3437 ( 
.A1(n_3200),
.A2(n_2862),
.B1(n_2851),
.B2(n_2786),
.Y(n_3437)
);

OAI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3334),
.A2(n_3350),
.B(n_3387),
.Y(n_3438)
);

AOI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3384),
.A2(n_3092),
.B(n_3089),
.Y(n_3439)
);

OAI21x1_ASAP7_75t_L g3440 ( 
.A1(n_3391),
.A2(n_3089),
.B(n_2741),
.Y(n_3440)
);

AOI21x1_ASAP7_75t_L g3441 ( 
.A1(n_3291),
.A2(n_2959),
.B(n_2892),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3221),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3217),
.B(n_3108),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3384),
.A2(n_2542),
.B(n_3187),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3219),
.B(n_3131),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3400),
.B(n_3075),
.Y(n_3446)
);

HB1xp67_ASAP7_75t_L g3447 ( 
.A(n_3374),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3286),
.B(n_2996),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3203),
.A2(n_2500),
.B(n_3182),
.Y(n_3449)
);

A2O1A1Ixp33_ASAP7_75t_L g3450 ( 
.A1(n_3241),
.A2(n_2622),
.B(n_3117),
.C(n_3112),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3329),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_L g3452 ( 
.A(n_3309),
.B(n_3059),
.Y(n_3452)
);

NOR2x1_ASAP7_75t_L g3453 ( 
.A(n_3389),
.B(n_3189),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3366),
.B(n_3081),
.Y(n_3454)
);

OR2x6_ASAP7_75t_SL g3455 ( 
.A(n_3323),
.B(n_3174),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3392),
.B(n_2952),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3289),
.B(n_2954),
.Y(n_3457)
);

OAI22xp5_ASAP7_75t_L g3458 ( 
.A1(n_3212),
.A2(n_2835),
.B1(n_2330),
.B2(n_2962),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3351),
.Y(n_3459)
);

BUFx3_ASAP7_75t_L g3460 ( 
.A(n_3355),
.Y(n_3460)
);

AOI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3246),
.A2(n_2635),
.B1(n_2650),
.B2(n_2790),
.Y(n_3461)
);

INVx1_ASAP7_75t_SL g3462 ( 
.A(n_3343),
.Y(n_3462)
);

OR2x6_ASAP7_75t_L g3463 ( 
.A(n_3280),
.B(n_2861),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_L g3464 ( 
.A(n_3266),
.B(n_2635),
.Y(n_3464)
);

NOR2x1_ASAP7_75t_L g3465 ( 
.A(n_3291),
.B(n_2762),
.Y(n_3465)
);

OR2x6_ASAP7_75t_L g3466 ( 
.A(n_3280),
.B(n_2861),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3226),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3203),
.A2(n_2835),
.B(n_2746),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3358),
.Y(n_3469)
);

AOI22xp5_ASAP7_75t_L g3470 ( 
.A1(n_3265),
.A2(n_2650),
.B1(n_2790),
.B2(n_3097),
.Y(n_3470)
);

AOI22xp5_ASAP7_75t_SL g3471 ( 
.A1(n_3375),
.A2(n_2465),
.B1(n_2440),
.B2(n_2458),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3398),
.B(n_3097),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3227),
.Y(n_3473)
);

O2A1O1Ixp33_ASAP7_75t_SL g3474 ( 
.A1(n_3255),
.A2(n_2649),
.B(n_2588),
.C(n_2399),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3316),
.A2(n_2746),
.B(n_2743),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3228),
.Y(n_3476)
);

BUFx3_ASAP7_75t_L g3477 ( 
.A(n_3207),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3209),
.B(n_3403),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_3397),
.B(n_2851),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3406),
.B(n_2922),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_SL g3481 ( 
.A(n_3230),
.B(n_2440),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_3280),
.A2(n_2756),
.B(n_2743),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3294),
.A2(n_2756),
.B(n_2656),
.Y(n_3483)
);

BUFx2_ASAP7_75t_L g3484 ( 
.A(n_3214),
.Y(n_3484)
);

AOI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3300),
.A2(n_3279),
.B1(n_3304),
.B2(n_3295),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3412),
.B(n_2928),
.Y(n_3486)
);

BUFx12f_ASAP7_75t_L g3487 ( 
.A(n_3237),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3242),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3376),
.B(n_2862),
.Y(n_3489)
);

BUFx3_ASAP7_75t_L g3490 ( 
.A(n_3234),
.Y(n_3490)
);

CKINVDCx5p33_ASAP7_75t_R g3491 ( 
.A(n_3238),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3283),
.A2(n_2395),
.B(n_2492),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3259),
.B(n_2930),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3308),
.B(n_2936),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3222),
.B(n_2951),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3283),
.A2(n_2415),
.B(n_2364),
.Y(n_3496)
);

AOI33xp33_ASAP7_75t_L g3497 ( 
.A1(n_3343),
.A2(n_3380),
.A3(n_3388),
.B1(n_3378),
.B2(n_3251),
.B3(n_3256),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3363),
.Y(n_3498)
);

NOR2x1_ASAP7_75t_L g3499 ( 
.A(n_3404),
.B(n_2762),
.Y(n_3499)
);

AND2x4_ASAP7_75t_SL g3500 ( 
.A(n_3306),
.B(n_2819),
.Y(n_3500)
);

A2O1A1Ixp33_ASAP7_75t_L g3501 ( 
.A1(n_3230),
.A2(n_2628),
.B(n_2690),
.C(n_2686),
.Y(n_3501)
);

O2A1O1Ixp33_ASAP7_75t_L g3502 ( 
.A1(n_3279),
.A2(n_2628),
.B(n_2373),
.C(n_2390),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3254),
.Y(n_3503)
);

INVx1_ASAP7_75t_SL g3504 ( 
.A(n_3253),
.Y(n_3504)
);

BUFx3_ASAP7_75t_L g3505 ( 
.A(n_3322),
.Y(n_3505)
);

BUFx12f_ASAP7_75t_L g3506 ( 
.A(n_3257),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3376),
.B(n_2686),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3410),
.B(n_2564),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3284),
.A2(n_2415),
.B(n_2364),
.Y(n_3509)
);

AND2x2_ASAP7_75t_SL g3510 ( 
.A(n_3362),
.B(n_2690),
.Y(n_3510)
);

NAND3xp33_ASAP7_75t_L g3511 ( 
.A(n_3305),
.B(n_2505),
.C(n_2497),
.Y(n_3511)
);

CKINVDCx14_ASAP7_75t_R g3512 ( 
.A(n_3257),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3311),
.B(n_2568),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3284),
.A2(n_2467),
.B(n_2415),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3261),
.Y(n_3515)
);

INVx4_ASAP7_75t_L g3516 ( 
.A(n_3282),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3215),
.A2(n_2467),
.B(n_2415),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3303),
.B(n_2568),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3281),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3359),
.B(n_2508),
.Y(n_3520)
);

AND2x6_ASAP7_75t_L g3521 ( 
.A(n_3252),
.B(n_2513),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3270),
.B(n_2819),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3275),
.B(n_2512),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_3299),
.B(n_2898),
.Y(n_3524)
);

CKINVDCx20_ASAP7_75t_R g3525 ( 
.A(n_3345),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3361),
.B(n_2694),
.Y(n_3526)
);

NAND2x1p5_ASAP7_75t_L g3527 ( 
.A(n_3393),
.B(n_3362),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_R g3528 ( 
.A(n_3407),
.B(n_2705),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_R g3529 ( 
.A(n_3407),
.B(n_2715),
.Y(n_3529)
);

INVx1_ASAP7_75t_SL g3530 ( 
.A(n_3258),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_SL g3531 ( 
.A(n_3393),
.B(n_2898),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3298),
.B(n_2514),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_3354),
.B(n_2694),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3247),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3250),
.Y(n_3535)
);

NOR3xp33_ASAP7_75t_L g3536 ( 
.A(n_3340),
.B(n_2472),
.C(n_2451),
.Y(n_3536)
);

O2A1O1Ixp33_ASAP7_75t_SL g3537 ( 
.A1(n_3331),
.A2(n_2740),
.B(n_2913),
.C(n_2745),
.Y(n_3537)
);

O2A1O1Ixp5_ASAP7_75t_L g3538 ( 
.A1(n_3370),
.A2(n_2748),
.B(n_2765),
.C(n_2900),
.Y(n_3538)
);

AOI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3215),
.A2(n_3277),
.B(n_3391),
.Y(n_3539)
);

AOI22xp33_ASAP7_75t_L g3540 ( 
.A1(n_3304),
.A2(n_2643),
.B1(n_2894),
.B2(n_2458),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3307),
.Y(n_3541)
);

O2A1O1Ixp33_ASAP7_75t_L g3542 ( 
.A1(n_3326),
.A2(n_2528),
.B(n_2531),
.C(n_2518),
.Y(n_3542)
);

BUFx2_ASAP7_75t_L g3543 ( 
.A(n_3248),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_3314),
.B(n_3341),
.Y(n_3544)
);

BUFx2_ASAP7_75t_L g3545 ( 
.A(n_3248),
.Y(n_3545)
);

O2A1O1Ixp5_ASAP7_75t_L g3546 ( 
.A1(n_3277),
.A2(n_2748),
.B(n_2765),
.C(n_2900),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3252),
.A2(n_2481),
.B(n_2467),
.Y(n_3547)
);

OAI22xp5_ASAP7_75t_L g3548 ( 
.A1(n_3350),
.A2(n_2330),
.B1(n_2413),
.B2(n_2365),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3387),
.A2(n_2481),
.B(n_2467),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3347),
.B(n_3349),
.Y(n_3550)
);

OAI21x1_ASAP7_75t_L g3551 ( 
.A1(n_3409),
.A2(n_2741),
.B(n_2723),
.Y(n_3551)
);

AND2x4_ASAP7_75t_L g3552 ( 
.A(n_3204),
.B(n_2740),
.Y(n_3552)
);

OAI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3409),
.A2(n_2723),
.B(n_2521),
.Y(n_3553)
);

AO21x1_ASAP7_75t_L g3554 ( 
.A1(n_3368),
.A2(n_2904),
.B(n_2521),
.Y(n_3554)
);

A2O1A1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_3369),
.A2(n_2451),
.B(n_2486),
.C(n_2472),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3373),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3262),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3271),
.B(n_2904),
.Y(n_3558)
);

A2O1A1Ixp33_ASAP7_75t_SL g3559 ( 
.A1(n_3201),
.A2(n_2486),
.B(n_2541),
.C(n_2535),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3236),
.B(n_2715),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3393),
.B(n_2715),
.Y(n_3561)
);

OAI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3225),
.A2(n_2413),
.B1(n_2365),
.B2(n_2513),
.Y(n_3562)
);

AOI21xp5_ASAP7_75t_L g3563 ( 
.A1(n_3325),
.A2(n_2481),
.B(n_2758),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3386),
.B(n_2522),
.Y(n_3564)
);

INVx2_ASAP7_75t_SL g3565 ( 
.A(n_3208),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_R g3566 ( 
.A(n_3208),
.B(n_2716),
.Y(n_3566)
);

O2A1O1Ixp5_ASAP7_75t_L g3567 ( 
.A1(n_3368),
.A2(n_2768),
.B(n_2772),
.C(n_2758),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3379),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3267),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3260),
.B(n_2522),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3273),
.Y(n_3571)
);

AO21x1_ASAP7_75t_L g3572 ( 
.A1(n_3325),
.A2(n_2523),
.B(n_2883),
.Y(n_3572)
);

INVx4_ASAP7_75t_L g3573 ( 
.A(n_3282),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3356),
.B(n_2523),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3276),
.Y(n_3575)
);

NOR3xp33_ASAP7_75t_L g3576 ( 
.A(n_3269),
.B(n_2457),
.C(n_2445),
.Y(n_3576)
);

AOI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_3413),
.A2(n_2643),
.B1(n_2440),
.B2(n_2458),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3318),
.Y(n_3578)
);

O2A1O1Ixp33_ASAP7_75t_L g3579 ( 
.A1(n_3272),
.A2(n_2894),
.B(n_2883),
.C(n_2745),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3396),
.B(n_2716),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3394),
.A2(n_2481),
.B(n_2804),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3394),
.A2(n_2850),
.B(n_2804),
.Y(n_3582)
);

AO22x1_ASAP7_75t_L g3583 ( 
.A1(n_3268),
.A2(n_2440),
.B1(n_2458),
.B2(n_2643),
.Y(n_3583)
);

OAI22x1_ASAP7_75t_L g3584 ( 
.A1(n_3245),
.A2(n_2917),
.B1(n_2926),
.B2(n_2826),
.Y(n_3584)
);

AO21x2_ASAP7_75t_L g3585 ( 
.A1(n_3290),
.A2(n_2917),
.B(n_2926),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3310),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3327),
.A2(n_2768),
.B1(n_2798),
.B2(n_2772),
.Y(n_3587)
);

AOI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3413),
.A2(n_2440),
.B1(n_2458),
.B2(n_2826),
.Y(n_3588)
);

OAI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_3377),
.A2(n_2798),
.B1(n_2882),
.B2(n_2850),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3385),
.Y(n_3590)
);

AOI21xp33_ASAP7_75t_L g3591 ( 
.A1(n_3377),
.A2(n_2882),
.B(n_2736),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3399),
.A2(n_2913),
.B(n_2736),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3399),
.A2(n_2945),
.B(n_2854),
.Y(n_3593)
);

OAI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3301),
.A2(n_3324),
.B1(n_3287),
.B2(n_3292),
.Y(n_3594)
);

AOI22x1_ASAP7_75t_L g3595 ( 
.A1(n_3395),
.A2(n_2725),
.B1(n_2716),
.B2(n_2834),
.Y(n_3595)
);

AOI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3413),
.A2(n_2834),
.B1(n_2854),
.B2(n_2945),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3317),
.Y(n_3597)
);

OAI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3287),
.A2(n_3292),
.B1(n_3336),
.B2(n_3408),
.Y(n_3598)
);

BUFx3_ASAP7_75t_L g3599 ( 
.A(n_3328),
.Y(n_3599)
);

AOI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3290),
.A2(n_3336),
.B(n_3338),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3319),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3278),
.B(n_2725),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3320),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3332),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3263),
.B(n_2725),
.Y(n_3605)
);

INVx2_ASAP7_75t_SL g3606 ( 
.A(n_3321),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3402),
.B(n_2561),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3338),
.A2(n_2734),
.B(n_2967),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_3383),
.B(n_2734),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3383),
.B(n_2734),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3335),
.B(n_2561),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3342),
.B(n_2561),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3352),
.B(n_2773),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_SL g3614 ( 
.A(n_3249),
.B(n_3352),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3201),
.A2(n_2970),
.B(n_2967),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_3205),
.A2(n_2970),
.B(n_2561),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_3249),
.B(n_2569),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3344),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3353),
.B(n_2569),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3205),
.A2(n_2569),
.B(n_2773),
.Y(n_3620)
);

A2O1A1Ixp33_ASAP7_75t_L g3621 ( 
.A1(n_3411),
.A2(n_2569),
.B(n_2960),
.C(n_2801),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3357),
.Y(n_3622)
);

AO22x1_ASAP7_75t_L g3623 ( 
.A1(n_3235),
.A2(n_2960),
.B1(n_2801),
.B2(n_2818),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3249),
.B(n_1796),
.Y(n_3624)
);

BUFx6f_ASAP7_75t_L g3625 ( 
.A(n_3220),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3364),
.B(n_171),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3312),
.B(n_3360),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_L g3628 ( 
.A(n_3263),
.B(n_171),
.Y(n_3628)
);

NOR2x1p5_ASAP7_75t_L g3629 ( 
.A(n_3401),
.B(n_2960),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_3312),
.A2(n_2960),
.B1(n_2801),
.B2(n_2818),
.Y(n_3630)
);

CKINVDCx10_ASAP7_75t_R g3631 ( 
.A(n_3333),
.Y(n_3631)
);

O2A1O1Ixp5_ASAP7_75t_L g3632 ( 
.A1(n_3293),
.A2(n_2801),
.B(n_2818),
.C(n_2755),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3586),
.Y(n_3633)
);

BUFx6f_ASAP7_75t_L g3634 ( 
.A(n_3505),
.Y(n_3634)
);

OAI21x1_ASAP7_75t_L g3635 ( 
.A1(n_3517),
.A2(n_3296),
.B(n_3293),
.Y(n_3635)
);

BUFx6f_ASAP7_75t_L g3636 ( 
.A(n_3599),
.Y(n_3636)
);

OAI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3419),
.A2(n_3367),
.B(n_3296),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_3504),
.B(n_3367),
.Y(n_3638)
);

A2O1A1Ixp33_ASAP7_75t_L g3639 ( 
.A1(n_3438),
.A2(n_3337),
.B(n_3382),
.C(n_3372),
.Y(n_3639)
);

NAND3xp33_ASAP7_75t_L g3640 ( 
.A(n_3485),
.B(n_3315),
.C(n_3302),
.Y(n_3640)
);

A2O1A1Ixp33_ASAP7_75t_L g3641 ( 
.A1(n_3438),
.A2(n_3401),
.B(n_3224),
.C(n_3216),
.Y(n_3641)
);

OR2x2_ASAP7_75t_L g3642 ( 
.A(n_3544),
.B(n_3339),
.Y(n_3642)
);

OAI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3420),
.A2(n_3213),
.B(n_3210),
.Y(n_3643)
);

AO31x2_ASAP7_75t_L g3644 ( 
.A1(n_3572),
.A2(n_3348),
.A3(n_3297),
.B(n_3339),
.Y(n_3644)
);

OAI21x1_ASAP7_75t_L g3645 ( 
.A1(n_3496),
.A2(n_3264),
.B(n_3224),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3431),
.B(n_3339),
.Y(n_3646)
);

BUFx3_ASAP7_75t_L g3647 ( 
.A(n_3460),
.Y(n_3647)
);

AOI21x1_ASAP7_75t_L g3648 ( 
.A1(n_3428),
.A2(n_3243),
.B(n_3339),
.Y(n_3648)
);

AOI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3439),
.A2(n_3426),
.B(n_3549),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3414),
.Y(n_3650)
);

NOR2xp67_ASAP7_75t_SL g3651 ( 
.A(n_3506),
.B(n_3282),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3442),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3415),
.B(n_3339),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3462),
.B(n_3210),
.Y(n_3654)
);

NAND3xp33_ASAP7_75t_L g3655 ( 
.A(n_3422),
.B(n_3315),
.C(n_3302),
.Y(n_3655)
);

BUFx6f_ASAP7_75t_L g3656 ( 
.A(n_3625),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3467),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3603),
.Y(n_3658)
);

AOI211x1_ASAP7_75t_L g3659 ( 
.A1(n_3432),
.A2(n_173),
.B(n_190),
.C(n_181),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3540),
.A2(n_3216),
.B1(n_3288),
.B2(n_3297),
.Y(n_3660)
);

A2O1A1Ixp33_ASAP7_75t_L g3661 ( 
.A1(n_3435),
.A2(n_3315),
.B(n_3346),
.C(n_3302),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3604),
.Y(n_3662)
);

NAND2x1p5_ASAP7_75t_L g3663 ( 
.A(n_3453),
.B(n_3489),
.Y(n_3663)
);

OAI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_3449),
.A2(n_3213),
.B(n_3210),
.Y(n_3664)
);

OAI21x1_ASAP7_75t_SL g3665 ( 
.A1(n_3608),
.A2(n_3288),
.B(n_3348),
.Y(n_3665)
);

AOI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3501),
.A2(n_3210),
.B(n_3213),
.Y(n_3666)
);

BUFx6f_ASAP7_75t_L g3667 ( 
.A(n_3625),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3427),
.A2(n_3213),
.B(n_3220),
.Y(n_3668)
);

AO21x1_ASAP7_75t_L g3669 ( 
.A1(n_3422),
.A2(n_57),
.B(n_58),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3444),
.A2(n_3232),
.B(n_3220),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3538),
.A2(n_3240),
.B(n_3232),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3470),
.B(n_3346),
.Y(n_3672)
);

OA21x2_ASAP7_75t_L g3673 ( 
.A1(n_3509),
.A2(n_2818),
.B(n_2755),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3462),
.B(n_3346),
.Y(n_3674)
);

AO21x1_ASAP7_75t_L g3675 ( 
.A1(n_3598),
.A2(n_57),
.B(n_58),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3473),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3476),
.Y(n_3677)
);

INVx3_ASAP7_75t_L g3678 ( 
.A(n_3424),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3550),
.B(n_3381),
.Y(n_3679)
);

AND2x4_ASAP7_75t_L g3680 ( 
.A(n_3504),
.B(n_3381),
.Y(n_3680)
);

OAI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3579),
.A2(n_2755),
.B(n_1796),
.Y(n_3681)
);

AOI21x1_ASAP7_75t_SL g3682 ( 
.A1(n_3421),
.A2(n_173),
.B(n_172),
.Y(n_3682)
);

AOI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3475),
.A2(n_3240),
.B(n_3232),
.Y(n_3683)
);

OAI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3514),
.A2(n_2755),
.B(n_1796),
.Y(n_3684)
);

O2A1O1Ixp5_ASAP7_75t_L g3685 ( 
.A1(n_3547),
.A2(n_3381),
.B(n_61),
.C(n_59),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3581),
.A2(n_3240),
.B(n_1761),
.Y(n_3686)
);

OAI21x1_ASAP7_75t_L g3687 ( 
.A1(n_3553),
.A2(n_1761),
.B(n_1724),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3543),
.B(n_690),
.Y(n_3688)
);

HB1xp67_ASAP7_75t_L g3689 ( 
.A(n_3447),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3618),
.Y(n_3690)
);

AOI21xp33_ASAP7_75t_L g3691 ( 
.A1(n_3584),
.A2(n_59),
.B(n_60),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3545),
.B(n_690),
.Y(n_3692)
);

BUFx2_ASAP7_75t_L g3693 ( 
.A(n_3484),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3548),
.A2(n_3468),
.B(n_3481),
.Y(n_3694)
);

AND2x4_ASAP7_75t_L g3695 ( 
.A(n_3530),
.B(n_59),
.Y(n_3695)
);

INVxp67_ASAP7_75t_L g3696 ( 
.A(n_3478),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3448),
.B(n_172),
.Y(n_3697)
);

OAI21x1_ASAP7_75t_L g3698 ( 
.A1(n_3563),
.A2(n_1761),
.B(n_1724),
.Y(n_3698)
);

NAND3xp33_ASAP7_75t_L g3699 ( 
.A(n_3497),
.B(n_60),
.C(n_61),
.Y(n_3699)
);

OA21x2_ASAP7_75t_L g3700 ( 
.A1(n_3440),
.A2(n_69),
.B(n_60),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3530),
.B(n_174),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3433),
.A2(n_1761),
.B(n_1724),
.Y(n_3702)
);

HB1xp67_ASAP7_75t_L g3703 ( 
.A(n_3594),
.Y(n_3703)
);

NOR2xp33_ASAP7_75t_L g3704 ( 
.A(n_3418),
.B(n_3452),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3556),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3594),
.B(n_175),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3598),
.B(n_3425),
.Y(n_3707)
);

A2O1A1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3416),
.A2(n_3450),
.B(n_3417),
.C(n_3464),
.Y(n_3708)
);

OR2x2_ASAP7_75t_L g3709 ( 
.A(n_3488),
.B(n_3503),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3429),
.B(n_176),
.Y(n_3710)
);

BUFx3_ASAP7_75t_L g3711 ( 
.A(n_3477),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3515),
.Y(n_3712)
);

AOI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3416),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3713)
);

AOI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3548),
.A2(n_3481),
.B(n_3593),
.Y(n_3714)
);

AO21x1_ASAP7_75t_L g3715 ( 
.A1(n_3472),
.A2(n_3417),
.B(n_3443),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3568),
.B(n_176),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3519),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_3546),
.A2(n_1761),
.B(n_1724),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3474),
.A2(n_1724),
.B(n_62),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3492),
.A2(n_62),
.B(n_63),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3541),
.Y(n_3721)
);

OA22x2_ASAP7_75t_L g3722 ( 
.A1(n_3424),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3537),
.A2(n_64),
.B(n_65),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_L g3724 ( 
.A(n_3631),
.B(n_177),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3597),
.Y(n_3725)
);

OAI21x1_ASAP7_75t_L g3726 ( 
.A1(n_3436),
.A2(n_66),
.B(n_67),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3590),
.B(n_177),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3457),
.B(n_178),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3601),
.B(n_178),
.Y(n_3729)
);

CKINVDCx11_ASAP7_75t_R g3730 ( 
.A(n_3487),
.Y(n_3730)
);

A2O1A1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3539),
.A2(n_180),
.B(n_181),
.C(n_179),
.Y(n_3731)
);

AO31x2_ASAP7_75t_L g3732 ( 
.A1(n_3554),
.A2(n_68),
.A3(n_66),
.B(n_67),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3482),
.A2(n_67),
.B(n_68),
.Y(n_3733)
);

BUFx3_ASAP7_75t_L g3734 ( 
.A(n_3490),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3441),
.A2(n_68),
.B(n_69),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3622),
.B(n_179),
.Y(n_3736)
);

OR2x2_ASAP7_75t_L g3737 ( 
.A(n_3627),
.B(n_180),
.Y(n_3737)
);

INVx3_ASAP7_75t_L g3738 ( 
.A(n_3527),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_3507),
.A2(n_70),
.B(n_71),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3526),
.B(n_698),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3551),
.A2(n_70),
.B(n_71),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3542),
.A2(n_71),
.B(n_72),
.Y(n_3742)
);

AOI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3621),
.A2(n_72),
.B(n_73),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3454),
.B(n_182),
.Y(n_3744)
);

BUFx6f_ASAP7_75t_L g3745 ( 
.A(n_3625),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3483),
.A2(n_72),
.B(n_73),
.Y(n_3746)
);

OA21x2_ASAP7_75t_L g3747 ( 
.A1(n_3567),
.A2(n_82),
.B(n_74),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3456),
.B(n_183),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3451),
.B(n_3459),
.Y(n_3749)
);

AOI211x1_ASAP7_75t_L g3750 ( 
.A1(n_3626),
.A2(n_194),
.B(n_202),
.C(n_186),
.Y(n_3750)
);

NAND3x1_ASAP7_75t_L g3751 ( 
.A(n_3461),
.B(n_74),
.C(n_75),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3469),
.B(n_183),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3600),
.A2(n_74),
.B(n_75),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_3582),
.A2(n_76),
.B(n_77),
.Y(n_3754)
);

NAND3x1_ASAP7_75t_L g3755 ( 
.A(n_3602),
.B(n_76),
.C(n_77),
.Y(n_3755)
);

OAI22xp5_ASAP7_75t_L g3756 ( 
.A1(n_3455),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_3756)
);

INVx2_ASAP7_75t_SL g3757 ( 
.A(n_3606),
.Y(n_3757)
);

A2O1A1Ixp33_ASAP7_75t_L g3758 ( 
.A1(n_3502),
.A2(n_186),
.B(n_187),
.C(n_185),
.Y(n_3758)
);

BUFx10_ASAP7_75t_L g3759 ( 
.A(n_3558),
.Y(n_3759)
);

AOI21xp33_ASAP7_75t_L g3760 ( 
.A1(n_3430),
.A2(n_78),
.B(n_79),
.Y(n_3760)
);

CKINVDCx5p33_ASAP7_75t_R g3761 ( 
.A(n_3491),
.Y(n_3761)
);

AOI21x1_ASAP7_75t_L g3762 ( 
.A1(n_3531),
.A2(n_78),
.B(n_79),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3498),
.B(n_185),
.Y(n_3763)
);

CKINVDCx20_ASAP7_75t_R g3764 ( 
.A(n_3525),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3592),
.A2(n_79),
.B(n_80),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3534),
.B(n_188),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3535),
.Y(n_3767)
);

CKINVDCx5p33_ASAP7_75t_R g3768 ( 
.A(n_3512),
.Y(n_3768)
);

AOI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3561),
.A2(n_80),
.B(n_81),
.Y(n_3769)
);

OAI21x1_ASAP7_75t_L g3770 ( 
.A1(n_3632),
.A2(n_80),
.B(n_81),
.Y(n_3770)
);

OAI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3434),
.A2(n_81),
.B(n_82),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3434),
.A2(n_82),
.B(n_83),
.Y(n_3772)
);

AOI21x1_ASAP7_75t_L g3773 ( 
.A1(n_3624),
.A2(n_83),
.B(n_85),
.Y(n_3773)
);

INVx3_ASAP7_75t_L g3774 ( 
.A(n_3527),
.Y(n_3774)
);

A2O1A1Ixp33_ASAP7_75t_L g3775 ( 
.A1(n_3471),
.A2(n_189),
.B(n_190),
.C(n_188),
.Y(n_3775)
);

OAI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3511),
.A2(n_92),
.B(n_83),
.Y(n_3776)
);

BUFx2_ASAP7_75t_L g3777 ( 
.A(n_3566),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3557),
.B(n_191),
.Y(n_3778)
);

INVx3_ASAP7_75t_L g3779 ( 
.A(n_3569),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3620),
.A2(n_85),
.B(n_86),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3533),
.B(n_688),
.Y(n_3781)
);

O2A1O1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_3559),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_3782)
);

OAI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3522),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3783)
);

OR2x6_ASAP7_75t_L g3784 ( 
.A(n_3463),
.B(n_192),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3571),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3580),
.B(n_3560),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3628),
.B(n_693),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_SL g3788 ( 
.A1(n_3577),
.A2(n_193),
.B(n_192),
.Y(n_3788)
);

OAI21x1_ASAP7_75t_L g3789 ( 
.A1(n_3589),
.A2(n_90),
.B(n_91),
.Y(n_3789)
);

BUFx3_ASAP7_75t_L g3790 ( 
.A(n_3565),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3575),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3589),
.A2(n_90),
.B(n_91),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3578),
.B(n_193),
.Y(n_3793)
);

CKINVDCx20_ASAP7_75t_R g3794 ( 
.A(n_3500),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3583),
.A2(n_92),
.B(n_93),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3510),
.A2(n_92),
.B(n_93),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3495),
.B(n_194),
.Y(n_3797)
);

OAI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3430),
.A2(n_102),
.B(n_94),
.Y(n_3798)
);

NOR2xp33_ASAP7_75t_L g3799 ( 
.A(n_3605),
.B(n_195),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3445),
.B(n_196),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3423),
.B(n_3570),
.Y(n_3801)
);

BUFx8_ASAP7_75t_L g3802 ( 
.A(n_3552),
.Y(n_3802)
);

BUFx2_ASAP7_75t_L g3803 ( 
.A(n_3528),
.Y(n_3803)
);

OAI21x1_ASAP7_75t_L g3804 ( 
.A1(n_3587),
.A2(n_94),
.B(n_95),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3536),
.A2(n_94),
.B(n_95),
.Y(n_3805)
);

OAI21x1_ASAP7_75t_L g3806 ( 
.A1(n_3587),
.A2(n_96),
.B(n_97),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3623),
.A2(n_96),
.B(n_97),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3446),
.Y(n_3808)
);

AOI221xp5_ASAP7_75t_SL g3809 ( 
.A1(n_3423),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.C(n_100),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3585),
.A2(n_98),
.B(n_99),
.Y(n_3810)
);

NAND2x1_ASAP7_75t_L g3811 ( 
.A(n_3516),
.B(n_196),
.Y(n_3811)
);

NOR2xp67_ASAP7_75t_L g3812 ( 
.A(n_3516),
.B(n_197),
.Y(n_3812)
);

AND2x4_ASAP7_75t_L g3813 ( 
.A(n_3614),
.B(n_98),
.Y(n_3813)
);

AOI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3617),
.A2(n_99),
.B(n_100),
.Y(n_3814)
);

CKINVDCx11_ASAP7_75t_R g3815 ( 
.A(n_3552),
.Y(n_3815)
);

OAI21x1_ASAP7_75t_L g3816 ( 
.A1(n_3458),
.A2(n_101),
.B(n_102),
.Y(n_3816)
);

OA21x2_ASAP7_75t_L g3817 ( 
.A1(n_3591),
.A2(n_101),
.B(n_102),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_L g3818 ( 
.A(n_3524),
.B(n_197),
.Y(n_3818)
);

OR2x2_ASAP7_75t_L g3819 ( 
.A(n_3607),
.B(n_3574),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3458),
.A2(n_101),
.B(n_103),
.Y(n_3820)
);

AO31x2_ASAP7_75t_L g3821 ( 
.A1(n_3630),
.A2(n_105),
.A3(n_103),
.B(n_104),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3480),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3585),
.A2(n_103),
.B(n_104),
.Y(n_3823)
);

AOI221x1_ASAP7_75t_L g3824 ( 
.A1(n_3591),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_3824)
);

BUFx4f_ASAP7_75t_SL g3825 ( 
.A(n_3609),
.Y(n_3825)
);

AND3x1_ASAP7_75t_L g3826 ( 
.A(n_3499),
.B(n_106),
.C(n_107),
.Y(n_3826)
);

OAI21x1_ASAP7_75t_L g3827 ( 
.A1(n_3630),
.A2(n_108),
.B(n_109),
.Y(n_3827)
);

OAI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3615),
.A2(n_109),
.B(n_110),
.Y(n_3828)
);

OAI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3588),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_3829)
);

OAI21x1_ASAP7_75t_L g3830 ( 
.A1(n_3562),
.A2(n_3564),
.B(n_3611),
.Y(n_3830)
);

OAI21x1_ASAP7_75t_L g3831 ( 
.A1(n_3562),
.A2(n_110),
.B(n_111),
.Y(n_3831)
);

NOR2xp67_ASAP7_75t_SL g3832 ( 
.A(n_3573),
.B(n_111),
.Y(n_3832)
);

OAI21x1_ASAP7_75t_L g3833 ( 
.A1(n_3612),
.A2(n_112),
.B(n_113),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_3619),
.Y(n_3834)
);

AND2x4_ASAP7_75t_L g3835 ( 
.A(n_3463),
.B(n_3466),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3493),
.B(n_198),
.Y(n_3836)
);

AOI21xp5_ASAP7_75t_L g3837 ( 
.A1(n_3616),
.A2(n_3520),
.B(n_3523),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3521),
.Y(n_3838)
);

CKINVDCx8_ASAP7_75t_R g3839 ( 
.A(n_3521),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3532),
.A2(n_112),
.B(n_113),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3521),
.Y(n_3841)
);

BUFx2_ASAP7_75t_L g3842 ( 
.A(n_3529),
.Y(n_3842)
);

OAI21x1_ASAP7_75t_L g3843 ( 
.A1(n_3465),
.A2(n_113),
.B(n_114),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3463),
.B(n_114),
.Y(n_3844)
);

NAND3xp33_ASAP7_75t_L g3845 ( 
.A(n_3508),
.B(n_114),
.C(n_115),
.Y(n_3845)
);

OAI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3596),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3846)
);

OAI21x1_ASAP7_75t_L g3847 ( 
.A1(n_3595),
.A2(n_3513),
.B(n_3494),
.Y(n_3847)
);

OA22x2_ASAP7_75t_L g3848 ( 
.A1(n_3610),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3848)
);

AO31x2_ASAP7_75t_L g3849 ( 
.A1(n_3573),
.A2(n_118),
.A3(n_116),
.B(n_117),
.Y(n_3849)
);

NAND3xp33_ASAP7_75t_L g3850 ( 
.A(n_3479),
.B(n_3486),
.C(n_3555),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3518),
.B(n_199),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3466),
.Y(n_3852)
);

OAI22xp5_ASAP7_75t_L g3853 ( 
.A1(n_3466),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_3853)
);

O2A1O1Ixp5_ASAP7_75t_L g3854 ( 
.A1(n_3613),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_3854)
);

NOR2xp67_ASAP7_75t_L g3855 ( 
.A(n_3521),
.B(n_200),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3576),
.Y(n_3856)
);

NOR2x1_ASAP7_75t_SL g3857 ( 
.A(n_3629),
.B(n_200),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3437),
.B(n_201),
.Y(n_3858)
);

OA21x2_ASAP7_75t_L g3859 ( 
.A1(n_3517),
.A2(n_119),
.B(n_120),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3414),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_3439),
.A2(n_121),
.B(n_122),
.Y(n_3861)
);

OAI21x1_ASAP7_75t_L g3862 ( 
.A1(n_3698),
.A2(n_121),
.B(n_122),
.Y(n_3862)
);

A2O1A1Ixp33_ASAP7_75t_L g3863 ( 
.A1(n_3699),
.A2(n_203),
.B(n_204),
.C(n_201),
.Y(n_3863)
);

AO31x2_ASAP7_75t_L g3864 ( 
.A1(n_3649),
.A2(n_125),
.A3(n_123),
.B(n_124),
.Y(n_3864)
);

AND2x6_ASAP7_75t_SL g3865 ( 
.A(n_3724),
.B(n_123),
.Y(n_3865)
);

O2A1O1Ixp5_ASAP7_75t_SL g3866 ( 
.A1(n_3856),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_3866)
);

A2O1A1Ixp33_ASAP7_75t_L g3867 ( 
.A1(n_3699),
.A2(n_204),
.B(n_205),
.C(n_203),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3664),
.A2(n_124),
.B(n_125),
.Y(n_3868)
);

NOR4xp25_ASAP7_75t_L g3869 ( 
.A(n_3755),
.B(n_128),
.C(n_126),
.D(n_127),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3639),
.B(n_3715),
.Y(n_3870)
);

NAND2x1_ASAP7_75t_L g3871 ( 
.A(n_3738),
.B(n_205),
.Y(n_3871)
);

O2A1O1Ixp33_ASAP7_75t_L g3872 ( 
.A1(n_3731),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_SL g3873 ( 
.A1(n_3664),
.A2(n_127),
.B(n_128),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3861),
.A2(n_129),
.B(n_130),
.Y(n_3874)
);

AOI221x1_ASAP7_75t_L g3875 ( 
.A1(n_3798),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.C(n_132),
.Y(n_3875)
);

AO21x2_ASAP7_75t_L g3876 ( 
.A1(n_3810),
.A2(n_131),
.B(n_132),
.Y(n_3876)
);

AOI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_3713),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_3877)
);

O2A1O1Ixp33_ASAP7_75t_L g3878 ( 
.A1(n_3798),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_3878)
);

CKINVDCx5p33_ASAP7_75t_R g3879 ( 
.A(n_3730),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3696),
.B(n_206),
.Y(n_3880)
);

AND2x4_ASAP7_75t_L g3881 ( 
.A(n_3852),
.B(n_208),
.Y(n_3881)
);

BUFx2_ASAP7_75t_R g3882 ( 
.A(n_3768),
.Y(n_3882)
);

AO21x1_ASAP7_75t_L g3883 ( 
.A1(n_3706),
.A2(n_133),
.B(n_135),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3646),
.B(n_208),
.Y(n_3884)
);

NAND3x1_ASAP7_75t_L g3885 ( 
.A(n_3713),
.B(n_136),
.C(n_137),
.Y(n_3885)
);

INVx3_ASAP7_75t_SL g3886 ( 
.A(n_3761),
.Y(n_3886)
);

INVx4_ASAP7_75t_L g3887 ( 
.A(n_3634),
.Y(n_3887)
);

AOI21xp5_ASAP7_75t_L g3888 ( 
.A1(n_3681),
.A2(n_3714),
.B(n_3666),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3650),
.Y(n_3889)
);

OAI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_3746),
.A2(n_136),
.B(n_137),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3681),
.A2(n_3708),
.B(n_3694),
.Y(n_3891)
);

OAI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3826),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_3892)
);

OA21x2_ASAP7_75t_L g3893 ( 
.A1(n_3823),
.A2(n_138),
.B(n_139),
.Y(n_3893)
);

NAND3x1_ASAP7_75t_L g3894 ( 
.A(n_3697),
.B(n_139),
.C(n_140),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3837),
.A2(n_141),
.B(n_142),
.Y(n_3895)
);

OAI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3720),
.A2(n_141),
.B(n_142),
.Y(n_3896)
);

CKINVDCx5p33_ASAP7_75t_R g3897 ( 
.A(n_3764),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3652),
.Y(n_3898)
);

OAI22x1_ASAP7_75t_L g3899 ( 
.A1(n_3693),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3657),
.Y(n_3900)
);

INVx3_ASAP7_75t_SL g3901 ( 
.A(n_3634),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3709),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3641),
.A2(n_143),
.B(n_144),
.Y(n_3903)
);

AOI221x1_ASAP7_75t_L g3904 ( 
.A1(n_3756),
.A2(n_143),
.B1(n_144),
.B2(n_209),
.C(n_210),
.Y(n_3904)
);

OR2x2_ASAP7_75t_L g3905 ( 
.A(n_3707),
.B(n_209),
.Y(n_3905)
);

OAI21x1_ASAP7_75t_L g3906 ( 
.A1(n_3702),
.A2(n_144),
.B(n_210),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3719),
.A2(n_211),
.B(n_212),
.Y(n_3907)
);

OAI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3826),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3676),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3677),
.Y(n_3910)
);

CKINVDCx6p67_ASAP7_75t_R g3911 ( 
.A(n_3647),
.Y(n_3911)
);

AO32x2_ASAP7_75t_L g3912 ( 
.A1(n_3783),
.A2(n_217),
.A3(n_214),
.B1(n_216),
.B2(n_218),
.Y(n_3912)
);

OAI21x1_ASAP7_75t_L g3913 ( 
.A1(n_3687),
.A2(n_216),
.B(n_218),
.Y(n_3913)
);

AOI221xp5_ASAP7_75t_L g3914 ( 
.A1(n_3659),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.C(n_222),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3705),
.Y(n_3915)
);

AO31x2_ASAP7_75t_L g3916 ( 
.A1(n_3824),
.A2(n_3669),
.A3(n_3675),
.B(n_3723),
.Y(n_3916)
);

OAI221xp5_ASAP7_75t_L g3917 ( 
.A1(n_3828),
.A2(n_223),
.B1(n_219),
.B2(n_222),
.C(n_224),
.Y(n_3917)
);

OAI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3754),
.A2(n_224),
.B(n_225),
.Y(n_3918)
);

AO31x2_ASAP7_75t_L g3919 ( 
.A1(n_3758),
.A2(n_3838),
.A3(n_3841),
.B(n_3742),
.Y(n_3919)
);

OAI21x1_ASAP7_75t_L g3920 ( 
.A1(n_3686),
.A2(n_226),
.B(n_227),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3653),
.B(n_226),
.Y(n_3921)
);

AO31x2_ASAP7_75t_L g3922 ( 
.A1(n_3718),
.A2(n_230),
.A3(n_227),
.B(n_229),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3643),
.A2(n_230),
.B(n_231),
.Y(n_3923)
);

OAI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3648),
.A2(n_231),
.B(n_232),
.Y(n_3924)
);

AO31x2_ASAP7_75t_L g3925 ( 
.A1(n_3668),
.A2(n_235),
.A3(n_233),
.B(n_234),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3712),
.Y(n_3926)
);

OAI21x1_ASAP7_75t_L g3927 ( 
.A1(n_3684),
.A2(n_234),
.B(n_236),
.Y(n_3927)
);

A2O1A1Ixp33_ASAP7_75t_L g3928 ( 
.A1(n_3776),
.A2(n_239),
.B(n_236),
.C(n_238),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3717),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3704),
.B(n_238),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3684),
.A2(n_239),
.B(n_240),
.Y(n_3931)
);

OAI21x1_ASAP7_75t_L g3932 ( 
.A1(n_3637),
.A2(n_241),
.B(n_243),
.Y(n_3932)
);

AND2x4_ASAP7_75t_L g3933 ( 
.A(n_3689),
.B(n_3642),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3721),
.Y(n_3934)
);

OA21x2_ASAP7_75t_L g3935 ( 
.A1(n_3741),
.A2(n_241),
.B(n_243),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3655),
.A2(n_244),
.B(n_245),
.Y(n_3936)
);

OAI21x1_ASAP7_75t_L g3937 ( 
.A1(n_3635),
.A2(n_244),
.B(n_245),
.Y(n_3937)
);

OAI21x1_ASAP7_75t_L g3938 ( 
.A1(n_3645),
.A2(n_246),
.B(n_247),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3819),
.B(n_246),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3786),
.B(n_248),
.Y(n_3940)
);

INVx3_ASAP7_75t_L g3941 ( 
.A(n_3634),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3678),
.B(n_248),
.Y(n_3942)
);

BUFx2_ASAP7_75t_R g3943 ( 
.A(n_3839),
.Y(n_3943)
);

AO31x2_ASAP7_75t_L g3944 ( 
.A1(n_3671),
.A2(n_252),
.A3(n_249),
.B(n_250),
.Y(n_3944)
);

O2A1O1Ixp33_ASAP7_75t_L g3945 ( 
.A1(n_3775),
.A2(n_252),
.B(n_249),
.C(n_250),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3703),
.B(n_253),
.Y(n_3946)
);

NOR2xp67_ASAP7_75t_L g3947 ( 
.A(n_3757),
.B(n_253),
.Y(n_3947)
);

BUFx6f_ASAP7_75t_L g3948 ( 
.A(n_3636),
.Y(n_3948)
);

OAI21x1_ASAP7_75t_L g3949 ( 
.A1(n_3847),
.A2(n_254),
.B(n_255),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3801),
.B(n_254),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3860),
.Y(n_3951)
);

O2A1O1Ixp33_ASAP7_75t_SL g3952 ( 
.A1(n_3661),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_3952)
);

AOI21xp5_ASAP7_75t_L g3953 ( 
.A1(n_3655),
.A2(n_3776),
.B(n_3788),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3808),
.B(n_257),
.Y(n_3954)
);

AOI22xp5_ASAP7_75t_SL g3955 ( 
.A1(n_3722),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3725),
.Y(n_3956)
);

OAI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3765),
.A2(n_260),
.B(n_262),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3633),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3678),
.B(n_262),
.Y(n_3959)
);

BUFx3_ASAP7_75t_L g3960 ( 
.A(n_3636),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3658),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3662),
.Y(n_3962)
);

NOR3xp33_ASAP7_75t_L g3963 ( 
.A(n_3760),
.B(n_264),
.C(n_265),
.Y(n_3963)
);

AND2x6_ASAP7_75t_L g3964 ( 
.A(n_3844),
.B(n_264),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3759),
.B(n_3640),
.Y(n_3965)
);

A2O1A1Ixp33_ASAP7_75t_L g3966 ( 
.A1(n_3685),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_3966)
);

AOI21xp5_ASAP7_75t_L g3967 ( 
.A1(n_3782),
.A2(n_266),
.B(n_267),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3670),
.A2(n_268),
.B(n_269),
.Y(n_3968)
);

INVx3_ASAP7_75t_SL g3969 ( 
.A(n_3636),
.Y(n_3969)
);

INVxp67_ASAP7_75t_SL g3970 ( 
.A(n_3779),
.Y(n_3970)
);

AO22x2_ASAP7_75t_L g3971 ( 
.A1(n_3659),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3690),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3767),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_SL g3974 ( 
.A(n_3759),
.B(n_3640),
.Y(n_3974)
);

OAI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3733),
.A2(n_270),
.B(n_271),
.Y(n_3975)
);

OAI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3840),
.A2(n_272),
.B(n_273),
.Y(n_3976)
);

AO32x2_ASAP7_75t_L g3977 ( 
.A1(n_3853),
.A2(n_3829),
.A3(n_3846),
.B1(n_3660),
.B2(n_3809),
.Y(n_3977)
);

AND2x4_ASAP7_75t_L g3978 ( 
.A(n_3638),
.B(n_273),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3822),
.B(n_274),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_SL g3980 ( 
.A(n_3651),
.B(n_3794),
.Y(n_3980)
);

AOI21xp5_ASAP7_75t_L g3981 ( 
.A1(n_3845),
.A2(n_274),
.B(n_275),
.Y(n_3981)
);

CKINVDCx5p33_ASAP7_75t_R g3982 ( 
.A(n_3815),
.Y(n_3982)
);

AOI221xp5_ASAP7_75t_SL g3983 ( 
.A1(n_3796),
.A2(n_3739),
.B1(n_3743),
.B2(n_3805),
.C(n_3795),
.Y(n_3983)
);

AOI21xp5_ASAP7_75t_L g3984 ( 
.A1(n_3845),
.A2(n_3683),
.B(n_3850),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3638),
.B(n_275),
.Y(n_3985)
);

OAI21x1_ASAP7_75t_L g3986 ( 
.A1(n_3726),
.A2(n_276),
.B(n_277),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_SL g3987 ( 
.A(n_3777),
.B(n_276),
.Y(n_3987)
);

BUFx3_ASAP7_75t_L g3988 ( 
.A(n_3711),
.Y(n_3988)
);

HB1xp67_ASAP7_75t_L g3989 ( 
.A(n_3779),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3738),
.B(n_277),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_SL g3991 ( 
.A(n_3734),
.B(n_278),
.Y(n_3991)
);

A2O1A1Ixp33_ASAP7_75t_L g3992 ( 
.A1(n_3809),
.A2(n_281),
.B(n_278),
.C(n_279),
.Y(n_3992)
);

BUFx3_ASAP7_75t_L g3993 ( 
.A(n_3790),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3834),
.B(n_282),
.Y(n_3994)
);

NAND3xp33_ASAP7_75t_SL g3995 ( 
.A(n_3854),
.B(n_283),
.C(n_284),
.Y(n_3995)
);

AO31x2_ASAP7_75t_L g3996 ( 
.A1(n_3654),
.A2(n_285),
.A3(n_283),
.B(n_284),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3680),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3850),
.A2(n_286),
.B(n_287),
.Y(n_3998)
);

AOI22xp33_ASAP7_75t_L g3999 ( 
.A1(n_3691),
.A2(n_3784),
.B1(n_3832),
.B2(n_3848),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3785),
.Y(n_4000)
);

OAI21x1_ASAP7_75t_L g4001 ( 
.A1(n_3753),
.A2(n_288),
.B(n_289),
.Y(n_4001)
);

OAI21x1_ASAP7_75t_L g4002 ( 
.A1(n_3735),
.A2(n_288),
.B(n_290),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3663),
.B(n_290),
.Y(n_4003)
);

BUFx6f_ASAP7_75t_L g4004 ( 
.A(n_3656),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3791),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3855),
.A2(n_291),
.B(n_292),
.Y(n_4006)
);

INVx4_ASAP7_75t_L g4007 ( 
.A(n_3656),
.Y(n_4007)
);

INVx3_ASAP7_75t_SL g4008 ( 
.A(n_3680),
.Y(n_4008)
);

OAI22xp33_ASAP7_75t_L g4009 ( 
.A1(n_3784),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4009)
);

INVx1_ASAP7_75t_SL g4010 ( 
.A(n_3803),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3749),
.Y(n_4011)
);

AOI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3855),
.A2(n_295),
.B(n_296),
.Y(n_4012)
);

AO31x2_ASAP7_75t_L g4013 ( 
.A1(n_3857),
.A2(n_299),
.A3(n_297),
.B(n_298),
.Y(n_4013)
);

INVx5_ASAP7_75t_L g4014 ( 
.A(n_3784),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_L g4015 ( 
.A(n_3737),
.B(n_298),
.Y(n_4015)
);

BUFx3_ASAP7_75t_L g4016 ( 
.A(n_3802),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_L g4017 ( 
.A(n_3818),
.B(n_299),
.Y(n_4017)
);

NOR2xp33_ASAP7_75t_L g4018 ( 
.A(n_3728),
.B(n_300),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3695),
.B(n_302),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3679),
.B(n_303),
.Y(n_4020)
);

A2O1A1Ixp33_ASAP7_75t_L g4021 ( 
.A1(n_3816),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_4021)
);

OAI21xp33_ASAP7_75t_L g4022 ( 
.A1(n_3858),
.A2(n_304),
.B(n_305),
.Y(n_4022)
);

NAND2xp33_ASAP7_75t_L g4023 ( 
.A(n_3751),
.B(n_306),
.Y(n_4023)
);

AO31x2_ASAP7_75t_L g4024 ( 
.A1(n_3807),
.A2(n_308),
.A3(n_306),
.B(n_307),
.Y(n_4024)
);

AOI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3672),
.A2(n_307),
.B(n_309),
.Y(n_4025)
);

OA21x2_ASAP7_75t_L g4026 ( 
.A1(n_3820),
.A2(n_310),
.B(n_311),
.Y(n_4026)
);

AO31x2_ASAP7_75t_L g4027 ( 
.A1(n_3674),
.A2(n_3732),
.A3(n_3747),
.B(n_3700),
.Y(n_4027)
);

INVx4_ASAP7_75t_L g4028 ( 
.A(n_3656),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3830),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3695),
.B(n_310),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3700),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3732),
.Y(n_4032)
);

OR2x2_ASAP7_75t_L g4033 ( 
.A(n_3710),
.B(n_311),
.Y(n_4033)
);

HB1xp67_ASAP7_75t_L g4034 ( 
.A(n_3644),
.Y(n_4034)
);

AO31x2_ASAP7_75t_L g4035 ( 
.A1(n_3732),
.A2(n_314),
.A3(n_312),
.B(n_313),
.Y(n_4035)
);

A2O1A1Ixp33_ASAP7_75t_L g4036 ( 
.A1(n_3831),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3665),
.A2(n_315),
.B(n_316),
.Y(n_4037)
);

NOR2xp33_ASAP7_75t_L g4038 ( 
.A(n_3744),
.B(n_3797),
.Y(n_4038)
);

A2O1A1Ixp33_ASAP7_75t_L g4039 ( 
.A1(n_3789),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_4039)
);

OAI21x1_ASAP7_75t_L g4040 ( 
.A1(n_3770),
.A2(n_317),
.B(n_318),
.Y(n_4040)
);

OAI21x1_ASAP7_75t_L g4041 ( 
.A1(n_3792),
.A2(n_319),
.B(n_321),
.Y(n_4041)
);

OAI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3804),
.A2(n_321),
.B(n_322),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3748),
.B(n_322),
.Y(n_4043)
);

OAI21x1_ASAP7_75t_L g4044 ( 
.A1(n_3888),
.A2(n_3859),
.B(n_3747),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3891),
.A2(n_3859),
.B(n_3851),
.Y(n_4045)
);

OAI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_4014),
.A2(n_3750),
.B1(n_3825),
.B2(n_3842),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3917),
.A2(n_3813),
.B1(n_3774),
.B2(n_3787),
.Y(n_4047)
);

OAI21x1_ASAP7_75t_L g4048 ( 
.A1(n_3984),
.A2(n_3806),
.B(n_3774),
.Y(n_4048)
);

AOI221xp5_ASAP7_75t_SL g4049 ( 
.A1(n_3870),
.A2(n_3701),
.B1(n_3800),
.B2(n_3799),
.C(n_3736),
.Y(n_4049)
);

AO21x2_ASAP7_75t_L g4050 ( 
.A1(n_4031),
.A2(n_3729),
.B(n_3812),
.Y(n_4050)
);

BUFx2_ASAP7_75t_L g4051 ( 
.A(n_3933),
.Y(n_4051)
);

OAI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_4014),
.A2(n_3812),
.B1(n_3811),
.B2(n_3817),
.Y(n_4052)
);

OA21x2_ASAP7_75t_L g4053 ( 
.A1(n_4029),
.A2(n_3833),
.B(n_3780),
.Y(n_4053)
);

AOI221xp5_ASAP7_75t_L g4054 ( 
.A1(n_3869),
.A2(n_3750),
.B1(n_3836),
.B2(n_3727),
.C(n_3716),
.Y(n_4054)
);

INVx6_ASAP7_75t_L g4055 ( 
.A(n_3948),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3901),
.B(n_3740),
.Y(n_4056)
);

OA21x2_ASAP7_75t_L g4057 ( 
.A1(n_4032),
.A2(n_4034),
.B(n_3974),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_4011),
.B(n_3933),
.Y(n_4058)
);

NOR2xp33_ASAP7_75t_L g4059 ( 
.A(n_3969),
.B(n_3781),
.Y(n_4059)
);

AND2x4_ASAP7_75t_L g4060 ( 
.A(n_3970),
.B(n_3835),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3889),
.Y(n_4061)
);

OAI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3953),
.A2(n_3772),
.B(n_3771),
.Y(n_4062)
);

OAI221xp5_ASAP7_75t_L g4063 ( 
.A1(n_3976),
.A2(n_3766),
.B1(n_3778),
.B2(n_3763),
.C(n_3752),
.Y(n_4063)
);

OAI21x1_ASAP7_75t_L g4064 ( 
.A1(n_3932),
.A2(n_3817),
.B(n_3762),
.Y(n_4064)
);

CKINVDCx8_ASAP7_75t_R g4065 ( 
.A(n_3865),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_L g4066 ( 
.A(n_4038),
.B(n_3802),
.Y(n_4066)
);

OAI21x1_ASAP7_75t_L g4067 ( 
.A1(n_3924),
.A2(n_3814),
.B(n_3769),
.Y(n_4067)
);

BUFx2_ASAP7_75t_L g4068 ( 
.A(n_4008),
.Y(n_4068)
);

OAI21x1_ASAP7_75t_L g4069 ( 
.A1(n_3937),
.A2(n_3827),
.B(n_3682),
.Y(n_4069)
);

HB1xp67_ASAP7_75t_L g4070 ( 
.A(n_3989),
.Y(n_4070)
);

OAI21x1_ASAP7_75t_L g4071 ( 
.A1(n_3949),
.A2(n_3913),
.B(n_3920),
.Y(n_4071)
);

OAI22xp5_ASAP7_75t_SL g4072 ( 
.A1(n_4014),
.A2(n_3844),
.B1(n_3813),
.B2(n_3835),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_L g4073 ( 
.A1(n_3938),
.A2(n_3673),
.B(n_3843),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3898),
.Y(n_4074)
);

AO31x2_ASAP7_75t_L g4075 ( 
.A1(n_3875),
.A2(n_3793),
.A3(n_3849),
.B(n_3821),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3934),
.Y(n_4076)
);

OAI21x1_ASAP7_75t_L g4077 ( 
.A1(n_3862),
.A2(n_3673),
.B(n_3773),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_3902),
.B(n_3821),
.Y(n_4078)
);

OAI21xp33_ASAP7_75t_SL g4079 ( 
.A1(n_3965),
.A2(n_3692),
.B(n_3688),
.Y(n_4079)
);

AND2x4_ASAP7_75t_L g4080 ( 
.A(n_3997),
.B(n_3644),
.Y(n_4080)
);

OAI21x1_ASAP7_75t_L g4081 ( 
.A1(n_3906),
.A2(n_3644),
.B(n_3821),
.Y(n_4081)
);

OAI21x1_ASAP7_75t_L g4082 ( 
.A1(n_3927),
.A2(n_3849),
.B(n_3745),
.Y(n_4082)
);

OA21x2_ASAP7_75t_L g4083 ( 
.A1(n_3921),
.A2(n_3849),
.B(n_3745),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3900),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3909),
.Y(n_4085)
);

INVx6_ASAP7_75t_L g4086 ( 
.A(n_3948),
.Y(n_4086)
);

BUFx6f_ASAP7_75t_L g4087 ( 
.A(n_4016),
.Y(n_4087)
);

BUFx5_ASAP7_75t_L g4088 ( 
.A(n_4005),
.Y(n_4088)
);

BUFx2_ASAP7_75t_L g4089 ( 
.A(n_3960),
.Y(n_4089)
);

BUFx4f_ASAP7_75t_L g4090 ( 
.A(n_3964),
.Y(n_4090)
);

OAI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_3895),
.A2(n_323),
.B(n_324),
.Y(n_4091)
);

OAI21x1_ASAP7_75t_L g4092 ( 
.A1(n_4037),
.A2(n_3745),
.B(n_3667),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3910),
.Y(n_4093)
);

BUFx12f_ASAP7_75t_L g4094 ( 
.A(n_3879),
.Y(n_4094)
);

CKINVDCx11_ASAP7_75t_R g4095 ( 
.A(n_3886),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3926),
.Y(n_4096)
);

OR2x6_ASAP7_75t_L g4097 ( 
.A(n_3873),
.B(n_3667),
.Y(n_4097)
);

AO32x2_ASAP7_75t_L g4098 ( 
.A1(n_3892),
.A2(n_3908),
.A3(n_3887),
.B1(n_4028),
.B2(n_4007),
.Y(n_4098)
);

INVx1_ASAP7_75t_SL g4099 ( 
.A(n_3911),
.Y(n_4099)
);

AO21x2_ASAP7_75t_L g4100 ( 
.A1(n_3884),
.A2(n_3667),
.B(n_323),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3929),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3958),
.B(n_324),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3951),
.Y(n_4103)
);

OAI21x1_ASAP7_75t_L g4104 ( 
.A1(n_4040),
.A2(n_325),
.B(n_326),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_SL g4105 ( 
.A1(n_3883),
.A2(n_325),
.B(n_326),
.Y(n_4105)
);

AOI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_4023),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3956),
.Y(n_4107)
);

AO21x2_ASAP7_75t_L g4108 ( 
.A1(n_3946),
.A2(n_328),
.B(n_329),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3868),
.A2(n_3998),
.B(n_3923),
.Y(n_4109)
);

AOI22x1_ASAP7_75t_L g4110 ( 
.A1(n_3955),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_4110)
);

AO21x2_ASAP7_75t_L g4111 ( 
.A1(n_3950),
.A2(n_332),
.B(n_333),
.Y(n_4111)
);

HB1xp67_ASAP7_75t_L g4112 ( 
.A(n_3915),
.Y(n_4112)
);

AOI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_3967),
.A2(n_709),
.B(n_334),
.Y(n_4113)
);

HB1xp67_ASAP7_75t_L g4114 ( 
.A(n_3962),
.Y(n_4114)
);

AOI22xp33_ASAP7_75t_SL g4115 ( 
.A1(n_3991),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3973),
.Y(n_4116)
);

BUFx6f_ASAP7_75t_L g4117 ( 
.A(n_4004),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_4000),
.Y(n_4118)
);

OAI21xp5_ASAP7_75t_SL g4119 ( 
.A1(n_3877),
.A2(n_335),
.B(n_337),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_4010),
.B(n_338),
.Y(n_4120)
);

AO21x2_ASAP7_75t_L g4121 ( 
.A1(n_3931),
.A2(n_3954),
.B(n_3979),
.Y(n_4121)
);

OAI21x1_ASAP7_75t_L g4122 ( 
.A1(n_4002),
.A2(n_338),
.B(n_339),
.Y(n_4122)
);

OAI21x1_ASAP7_75t_L g4123 ( 
.A1(n_3986),
.A2(n_4041),
.B(n_4001),
.Y(n_4123)
);

AO31x2_ASAP7_75t_L g4124 ( 
.A1(n_3992),
.A2(n_341),
.A3(n_339),
.B(n_340),
.Y(n_4124)
);

INVxp67_ASAP7_75t_L g4125 ( 
.A(n_3880),
.Y(n_4125)
);

OR2x6_ASAP7_75t_L g4126 ( 
.A(n_3988),
.B(n_340),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3961),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3972),
.B(n_701),
.Y(n_4128)
);

AND2x2_ASAP7_75t_SL g4129 ( 
.A(n_3980),
.B(n_341),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_4027),
.Y(n_4130)
);

BUFx2_ASAP7_75t_L g4131 ( 
.A(n_3941),
.Y(n_4131)
);

OAI21x1_ASAP7_75t_L g4132 ( 
.A1(n_3968),
.A2(n_342),
.B(n_343),
.Y(n_4132)
);

INVx3_ASAP7_75t_L g4133 ( 
.A(n_3993),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4027),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_4027),
.Y(n_4135)
);

OAI21x1_ASAP7_75t_L g4136 ( 
.A1(n_4006),
.A2(n_342),
.B(n_343),
.Y(n_4136)
);

AND2x4_ASAP7_75t_L g4137 ( 
.A(n_4004),
.B(n_344),
.Y(n_4137)
);

OAI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3936),
.A2(n_344),
.B(n_346),
.Y(n_4138)
);

INVxp67_ASAP7_75t_SL g4139 ( 
.A(n_3994),
.Y(n_4139)
);

AND2x4_ASAP7_75t_L g4140 ( 
.A(n_3942),
.B(n_347),
.Y(n_4140)
);

BUFx6f_ASAP7_75t_L g4141 ( 
.A(n_3871),
.Y(n_4141)
);

OAI21x1_ASAP7_75t_SL g4142 ( 
.A1(n_3878),
.A2(n_347),
.B(n_348),
.Y(n_4142)
);

OAI21x1_ASAP7_75t_L g4143 ( 
.A1(n_4012),
.A2(n_349),
.B(n_350),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_SL g4144 ( 
.A(n_3982),
.B(n_349),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4035),
.Y(n_4145)
);

AO31x2_ASAP7_75t_L g4146 ( 
.A1(n_3904),
.A2(n_353),
.A3(n_350),
.B(n_352),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4035),
.Y(n_4147)
);

A2O1A1Ixp33_ASAP7_75t_L g4148 ( 
.A1(n_3945),
.A2(n_700),
.B(n_354),
.C(n_352),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4035),
.Y(n_4149)
);

CKINVDCx6p67_ASAP7_75t_R g4150 ( 
.A(n_3964),
.Y(n_4150)
);

OAI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_3863),
.A2(n_356),
.B1(n_353),
.B2(n_355),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3864),
.Y(n_4152)
);

OAI21x1_ASAP7_75t_L g4153 ( 
.A1(n_3903),
.A2(n_355),
.B(n_356),
.Y(n_4153)
);

OAI22xp5_ASAP7_75t_L g4154 ( 
.A1(n_3867),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.Y(n_4154)
);

OAI21x1_ASAP7_75t_SL g4155 ( 
.A1(n_3981),
.A2(n_359),
.B(n_360),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3864),
.Y(n_4156)
);

AOI22xp5_ASAP7_75t_L g4157 ( 
.A1(n_3983),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3996),
.Y(n_4158)
);

HB1xp67_ASAP7_75t_L g4159 ( 
.A(n_3996),
.Y(n_4159)
);

BUFx12f_ASAP7_75t_L g4160 ( 
.A(n_3897),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3996),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3944),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3905),
.B(n_699),
.Y(n_4163)
);

BUFx2_ASAP7_75t_L g4164 ( 
.A(n_3959),
.Y(n_4164)
);

OAI21x1_ASAP7_75t_L g4165 ( 
.A1(n_3907),
.A2(n_362),
.B(n_363),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_3985),
.Y(n_4166)
);

INVx6_ASAP7_75t_L g4167 ( 
.A(n_3978),
.Y(n_4167)
);

INVx2_ASAP7_75t_SL g4168 ( 
.A(n_3990),
.Y(n_4168)
);

AND2x4_ASAP7_75t_L g4169 ( 
.A(n_3944),
.B(n_3919),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_L g4170 ( 
.A1(n_3963),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3944),
.Y(n_4171)
);

NOR2xp67_ASAP7_75t_L g4172 ( 
.A(n_4033),
.B(n_4043),
.Y(n_4172)
);

BUFx6f_ASAP7_75t_L g4173 ( 
.A(n_3881),
.Y(n_4173)
);

NOR2xp67_ASAP7_75t_SL g4174 ( 
.A(n_4025),
.B(n_364),
.Y(n_4174)
);

AO31x2_ASAP7_75t_L g4175 ( 
.A1(n_4036),
.A2(n_368),
.A3(n_366),
.B(n_367),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3939),
.B(n_699),
.Y(n_4176)
);

BUFx3_ASAP7_75t_L g4177 ( 
.A(n_4019),
.Y(n_4177)
);

AOI22x1_ASAP7_75t_L g4178 ( 
.A1(n_3899),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_4178)
);

NOR2xp67_ASAP7_75t_L g4179 ( 
.A(n_4020),
.B(n_370),
.Y(n_4179)
);

BUFx2_ASAP7_75t_SL g4180 ( 
.A(n_3947),
.Y(n_4180)
);

OAI22x1_ASAP7_75t_L g4181 ( 
.A1(n_4017),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_4181)
);

AOI22x1_ASAP7_75t_L g4182 ( 
.A1(n_3971),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3864),
.Y(n_4183)
);

AOI21x1_ASAP7_75t_L g4184 ( 
.A1(n_4003),
.A2(n_374),
.B(n_375),
.Y(n_4184)
);

INVx4_ASAP7_75t_L g4185 ( 
.A(n_3964),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3872),
.A2(n_376),
.B(n_377),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_SL g4187 ( 
.A1(n_3966),
.A2(n_376),
.B(n_377),
.Y(n_4187)
);

BUFx2_ASAP7_75t_R g4188 ( 
.A(n_3882),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3925),
.Y(n_4189)
);

OAI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_3928),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_4190)
);

OR2x6_ASAP7_75t_L g4191 ( 
.A(n_4042),
.B(n_378),
.Y(n_4191)
);

OA21x2_ASAP7_75t_L g4192 ( 
.A1(n_4039),
.A2(n_3914),
.B(n_4021),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3922),
.Y(n_4193)
);

BUFx12f_ASAP7_75t_L g4194 ( 
.A(n_4030),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_3987),
.B(n_380),
.Y(n_4195)
);

OA21x2_ASAP7_75t_L g4196 ( 
.A1(n_3874),
.A2(n_3957),
.B(n_3918),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4013),
.Y(n_4197)
);

AND2x4_ASAP7_75t_L g4198 ( 
.A(n_4048),
.B(n_3919),
.Y(n_4198)
);

A2O1A1Ixp33_ASAP7_75t_L g4199 ( 
.A1(n_4109),
.A2(n_3930),
.B(n_4022),
.C(n_3975),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4159),
.B(n_3922),
.Y(n_4200)
);

OR2x2_ASAP7_75t_L g4201 ( 
.A(n_4078),
.B(n_4058),
.Y(n_4201)
);

HB1xp67_ASAP7_75t_L g4202 ( 
.A(n_4070),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_4045),
.A2(n_3952),
.B(n_3890),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4101),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4101),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_4158),
.B(n_4161),
.Y(n_4206)
);

OAI21x1_ASAP7_75t_L g4207 ( 
.A1(n_4081),
.A2(n_3935),
.B(n_4026),
.Y(n_4207)
);

OR2x6_ASAP7_75t_L g4208 ( 
.A(n_4097),
.B(n_4185),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4088),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4103),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_4196),
.A2(n_3896),
.B(n_3995),
.Y(n_4211)
);

AO21x2_ASAP7_75t_L g4212 ( 
.A1(n_4130),
.A2(n_4009),
.B(n_3876),
.Y(n_4212)
);

AOI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_4196),
.A2(n_3971),
.B(n_3893),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4088),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4139),
.B(n_3922),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4103),
.Y(n_4216)
);

INVxp33_ASAP7_75t_L g4217 ( 
.A(n_4095),
.Y(n_4217)
);

OA21x2_ASAP7_75t_L g4218 ( 
.A1(n_4134),
.A2(n_3999),
.B(n_4015),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4107),
.Y(n_4219)
);

INVx2_ASAP7_75t_SL g4220 ( 
.A(n_4087),
.Y(n_4220)
);

OAI21x1_ASAP7_75t_L g4221 ( 
.A1(n_4044),
.A2(n_3935),
.B(n_4026),
.Y(n_4221)
);

INVx3_ASAP7_75t_L g4222 ( 
.A(n_4080),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4116),
.B(n_3893),
.Y(n_4223)
);

AOI21x1_ASAP7_75t_L g4224 ( 
.A1(n_4135),
.A2(n_3940),
.B(n_3925),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4107),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4068),
.B(n_3919),
.Y(n_4226)
);

AOI21xp5_ASAP7_75t_L g4227 ( 
.A1(n_4187),
.A2(n_4018),
.B(n_3977),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_4088),
.Y(n_4228)
);

AOI21xp5_ASAP7_75t_L g4229 ( 
.A1(n_4148),
.A2(n_3977),
.B(n_3916),
.Y(n_4229)
);

BUFx6f_ASAP7_75t_L g4230 ( 
.A(n_4087),
.Y(n_4230)
);

NOR2x1_ASAP7_75t_SL g4231 ( 
.A(n_4050),
.B(n_3943),
.Y(n_4231)
);

OAI21x1_ASAP7_75t_L g4232 ( 
.A1(n_4197),
.A2(n_4082),
.B(n_4147),
.Y(n_4232)
);

BUFx6f_ASAP7_75t_L g4233 ( 
.A(n_4087),
.Y(n_4233)
);

NOR2xp33_ASAP7_75t_L g4234 ( 
.A(n_4188),
.B(n_381),
.Y(n_4234)
);

OAI21x1_ASAP7_75t_SL g4235 ( 
.A1(n_4185),
.A2(n_3894),
.B(n_3912),
.Y(n_4235)
);

AO31x2_ASAP7_75t_L g4236 ( 
.A1(n_4147),
.A2(n_3912),
.A3(n_3925),
.B(n_3866),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4051),
.B(n_4013),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4060),
.B(n_4013),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4116),
.Y(n_4239)
);

OAI21x1_ASAP7_75t_L g4240 ( 
.A1(n_4149),
.A2(n_4145),
.B(n_4064),
.Y(n_4240)
);

OA21x2_ASAP7_75t_L g4241 ( 
.A1(n_4149),
.A2(n_3912),
.B(n_3977),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_4088),
.Y(n_4242)
);

AOI21x1_ASAP7_75t_L g4243 ( 
.A1(n_4172),
.A2(n_4128),
.B(n_4102),
.Y(n_4243)
);

AOI21xp5_ASAP7_75t_L g4244 ( 
.A1(n_4186),
.A2(n_3916),
.B(n_3885),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_SL g4245 ( 
.A(n_4090),
.B(n_4097),
.Y(n_4245)
);

OAI21x1_ASAP7_75t_L g4246 ( 
.A1(n_4162),
.A2(n_4024),
.B(n_3916),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4061),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4088),
.Y(n_4248)
);

AOI21xp33_ASAP7_75t_SL g4249 ( 
.A1(n_4144),
.A2(n_382),
.B(n_383),
.Y(n_4249)
);

OAI21x1_ASAP7_75t_L g4250 ( 
.A1(n_4171),
.A2(n_4024),
.B(n_382),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4114),
.B(n_4024),
.Y(n_4251)
);

AOI21xp5_ASAP7_75t_L g4252 ( 
.A1(n_4138),
.A2(n_383),
.B(n_384),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4074),
.Y(n_4253)
);

OA21x2_ASAP7_75t_L g4254 ( 
.A1(n_4189),
.A2(n_384),
.B(n_385),
.Y(n_4254)
);

AOI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_4119),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_4118),
.B(n_386),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4084),
.Y(n_4257)
);

OAI21x1_ASAP7_75t_L g4258 ( 
.A1(n_4193),
.A2(n_387),
.B(n_389),
.Y(n_4258)
);

AOI21x1_ASAP7_75t_L g4259 ( 
.A1(n_4163),
.A2(n_390),
.B(n_391),
.Y(n_4259)
);

CKINVDCx20_ASAP7_75t_R g4260 ( 
.A(n_4160),
.Y(n_4260)
);

AO31x2_ASAP7_75t_L g4261 ( 
.A1(n_4193),
.A2(n_394),
.A3(n_392),
.B(n_393),
.Y(n_4261)
);

NOR2xp33_ASAP7_75t_L g4262 ( 
.A(n_4125),
.B(n_392),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4085),
.B(n_395),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4093),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4096),
.Y(n_4265)
);

BUFx6f_ASAP7_75t_L g4266 ( 
.A(n_4094),
.Y(n_4266)
);

BUFx2_ASAP7_75t_L g4267 ( 
.A(n_4060),
.Y(n_4267)
);

OAI21x1_ASAP7_75t_L g4268 ( 
.A1(n_4057),
.A2(n_395),
.B(n_397),
.Y(n_4268)
);

AOI22xp33_ASAP7_75t_L g4269 ( 
.A1(n_4192),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_4269)
);

OAI21x1_ASAP7_75t_SL g4270 ( 
.A1(n_4182),
.A2(n_398),
.B(n_399),
.Y(n_4270)
);

NAND3xp33_ASAP7_75t_L g4271 ( 
.A(n_4157),
.B(n_400),
.C(n_401),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4127),
.Y(n_4272)
);

CKINVDCx5p33_ASAP7_75t_R g4273 ( 
.A(n_4180),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4152),
.B(n_400),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4112),
.Y(n_4275)
);

OAI21x1_ASAP7_75t_L g4276 ( 
.A1(n_4057),
.A2(n_401),
.B(n_402),
.Y(n_4276)
);

INVx4_ASAP7_75t_L g4277 ( 
.A(n_4126),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4152),
.B(n_402),
.Y(n_4278)
);

A2O1A1Ixp33_ASAP7_75t_L g4279 ( 
.A1(n_4090),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_4279)
);

OA21x2_ASAP7_75t_L g4280 ( 
.A1(n_4080),
.A2(n_403),
.B(n_404),
.Y(n_4280)
);

BUFx3_ASAP7_75t_L g4281 ( 
.A(n_4133),
.Y(n_4281)
);

AOI22x1_ASAP7_75t_L g4282 ( 
.A1(n_4181),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_4282)
);

AOI21xp33_ASAP7_75t_L g4283 ( 
.A1(n_4191),
.A2(n_406),
.B(n_408),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4076),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4131),
.Y(n_4285)
);

AO21x2_ASAP7_75t_L g4286 ( 
.A1(n_4156),
.A2(n_409),
.B(n_410),
.Y(n_4286)
);

INVx3_ASAP7_75t_L g4287 ( 
.A(n_4141),
.Y(n_4287)
);

OAI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_4113),
.A2(n_409),
.B(n_410),
.Y(n_4288)
);

OA21x2_ASAP7_75t_L g4289 ( 
.A1(n_4156),
.A2(n_413),
.B(n_414),
.Y(n_4289)
);

BUFx4f_ASAP7_75t_SL g4290 ( 
.A(n_4099),
.Y(n_4290)
);

BUFx2_ASAP7_75t_L g4291 ( 
.A(n_4089),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4164),
.Y(n_4292)
);

BUFx2_ASAP7_75t_L g4293 ( 
.A(n_4133),
.Y(n_4293)
);

BUFx3_ASAP7_75t_L g4294 ( 
.A(n_4194),
.Y(n_4294)
);

OAI21x1_ASAP7_75t_L g4295 ( 
.A1(n_4073),
.A2(n_413),
.B(n_414),
.Y(n_4295)
);

OA21x2_ASAP7_75t_L g4296 ( 
.A1(n_4183),
.A2(n_415),
.B(n_416),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4083),
.Y(n_4297)
);

BUFx3_ASAP7_75t_L g4298 ( 
.A(n_4173),
.Y(n_4298)
);

OA21x2_ASAP7_75t_L g4299 ( 
.A1(n_4169),
.A2(n_415),
.B(n_417),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4083),
.Y(n_4300)
);

INVxp67_ASAP7_75t_L g4301 ( 
.A(n_4108),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4169),
.Y(n_4302)
);

HB1xp67_ASAP7_75t_L g4303 ( 
.A(n_4053),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4053),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_4150),
.Y(n_4305)
);

AOI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_4195),
.A2(n_417),
.B(n_418),
.Y(n_4306)
);

BUFx12f_ASAP7_75t_L g4307 ( 
.A(n_4126),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4166),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4177),
.B(n_419),
.Y(n_4309)
);

AND2x4_ASAP7_75t_L g4310 ( 
.A(n_4092),
.B(n_420),
.Y(n_4310)
);

INVx3_ASAP7_75t_L g4311 ( 
.A(n_4141),
.Y(n_4311)
);

OAI21x1_ASAP7_75t_L g4312 ( 
.A1(n_4123),
.A2(n_421),
.B(n_422),
.Y(n_4312)
);

OAI21x1_ASAP7_75t_L g4313 ( 
.A1(n_4071),
.A2(n_4077),
.B(n_4062),
.Y(n_4313)
);

CKINVDCx11_ASAP7_75t_R g4314 ( 
.A(n_4065),
.Y(n_4314)
);

AOI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_4191),
.A2(n_421),
.B(n_422),
.Y(n_4315)
);

AO31x2_ASAP7_75t_L g4316 ( 
.A1(n_4046),
.A2(n_425),
.A3(n_423),
.B(n_424),
.Y(n_4316)
);

OAI21x1_ASAP7_75t_L g4317 ( 
.A1(n_4067),
.A2(n_423),
.B(n_424),
.Y(n_4317)
);

OR2x6_ASAP7_75t_L g4318 ( 
.A(n_4141),
.B(n_426),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4117),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_4192),
.A2(n_4182),
.B1(n_4121),
.B2(n_4110),
.Y(n_4320)
);

BUFx3_ASAP7_75t_L g4321 ( 
.A(n_4173),
.Y(n_4321)
);

NAND2x1p5_ASAP7_75t_L g4322 ( 
.A(n_4117),
.B(n_427),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4117),
.Y(n_4323)
);

OAI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4091),
.A2(n_428),
.B(n_429),
.Y(n_4324)
);

CKINVDCx11_ASAP7_75t_R g4325 ( 
.A(n_4140),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4055),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4049),
.B(n_428),
.Y(n_4327)
);

OAI21x1_ASAP7_75t_SL g4328 ( 
.A1(n_4105),
.A2(n_430),
.B(n_431),
.Y(n_4328)
);

AOI21xp33_ASAP7_75t_SL g4329 ( 
.A1(n_4129),
.A2(n_430),
.B(n_431),
.Y(n_4329)
);

OA21x2_ASAP7_75t_L g4330 ( 
.A1(n_4069),
.A2(n_432),
.B(n_433),
.Y(n_4330)
);

AND2x4_ASAP7_75t_L g4331 ( 
.A(n_4168),
.B(n_432),
.Y(n_4331)
);

OAI21x1_ASAP7_75t_L g4332 ( 
.A1(n_4104),
.A2(n_433),
.B(n_434),
.Y(n_4332)
);

AOI21xp5_ASAP7_75t_L g4333 ( 
.A1(n_4190),
.A2(n_435),
.B(n_436),
.Y(n_4333)
);

OA21x2_ASAP7_75t_L g4334 ( 
.A1(n_4054),
.A2(n_436),
.B(n_438),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4055),
.Y(n_4335)
);

OAI21xp33_ASAP7_75t_L g4336 ( 
.A1(n_4106),
.A2(n_438),
.B(n_439),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_4086),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4111),
.Y(n_4338)
);

OA21x2_ASAP7_75t_L g4339 ( 
.A1(n_4122),
.A2(n_439),
.B(n_440),
.Y(n_4339)
);

BUFx6f_ASAP7_75t_L g4340 ( 
.A(n_4137),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4059),
.B(n_440),
.Y(n_4341)
);

OAI21x1_ASAP7_75t_L g4342 ( 
.A1(n_4136),
.A2(n_442),
.B(n_443),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4100),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4086),
.Y(n_4344)
);

HB1xp67_ASAP7_75t_L g4345 ( 
.A(n_4075),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_4173),
.Y(n_4346)
);

A2O1A1Ixp33_ASAP7_75t_L g4347 ( 
.A1(n_4179),
.A2(n_4079),
.B(n_4174),
.C(n_4153),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4098),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4075),
.B(n_442),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4110),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4056),
.B(n_445),
.Y(n_4351)
);

AO21x2_ASAP7_75t_L g4352 ( 
.A1(n_4052),
.A2(n_4142),
.B(n_4155),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_4143),
.A2(n_446),
.B(n_447),
.Y(n_4353)
);

CKINVDCx16_ASAP7_75t_R g4354 ( 
.A(n_4072),
.Y(n_4354)
);

OA21x2_ASAP7_75t_L g4355 ( 
.A1(n_4176),
.A2(n_449),
.B(n_450),
.Y(n_4355)
);

NAND2x1p5_ASAP7_75t_L g4356 ( 
.A(n_4137),
.B(n_449),
.Y(n_4356)
);

AOI21xp5_ASAP7_75t_L g4357 ( 
.A1(n_4151),
.A2(n_450),
.B(n_451),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_4167),
.Y(n_4358)
);

OR2x2_ASAP7_75t_L g4359 ( 
.A(n_4120),
.B(n_451),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_4066),
.B(n_452),
.Y(n_4360)
);

OAI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_4047),
.A2(n_4132),
.B(n_4165),
.Y(n_4361)
);

OAI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_4178),
.A2(n_4115),
.B1(n_4170),
.B2(n_4154),
.Y(n_4362)
);

AOI22xp33_ASAP7_75t_L g4363 ( 
.A1(n_4229),
.A2(n_4178),
.B1(n_4063),
.B2(n_4167),
.Y(n_4363)
);

AOI222xp33_ASAP7_75t_L g4364 ( 
.A1(n_4324),
.A2(n_4140),
.B1(n_4098),
.B2(n_4146),
.C1(n_4124),
.C2(n_4075),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4293),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4267),
.B(n_4098),
.Y(n_4366)
);

AOI22xp33_ASAP7_75t_L g4367 ( 
.A1(n_4229),
.A2(n_4124),
.B1(n_4146),
.B2(n_4175),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4204),
.Y(n_4368)
);

AOI22xp33_ASAP7_75t_L g4369 ( 
.A1(n_4227),
.A2(n_4124),
.B1(n_4146),
.B2(n_4175),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4205),
.Y(n_4370)
);

INVx3_ASAP7_75t_L g4371 ( 
.A(n_4230),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4210),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4216),
.Y(n_4373)
);

OAI22xp33_ASAP7_75t_L g4374 ( 
.A1(n_4354),
.A2(n_4184),
.B1(n_4175),
.B2(n_454),
.Y(n_4374)
);

OAI22xp5_ASAP7_75t_L g4375 ( 
.A1(n_4227),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_4375)
);

BUFx4f_ASAP7_75t_SL g4376 ( 
.A(n_4260),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4219),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4343),
.B(n_455),
.Y(n_4378)
);

OAI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_4320),
.A2(n_4255),
.B1(n_4199),
.B2(n_4271),
.Y(n_4379)
);

AOI22xp33_ASAP7_75t_L g4380 ( 
.A1(n_4211),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_4380)
);

INVx3_ASAP7_75t_L g4381 ( 
.A(n_4230),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_4211),
.A2(n_460),
.B1(n_457),
.B2(n_458),
.Y(n_4382)
);

AOI22xp33_ASAP7_75t_SL g4383 ( 
.A1(n_4231),
.A2(n_463),
.B1(n_460),
.B2(n_462),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4291),
.Y(n_4384)
);

AOI222xp33_ASAP7_75t_L g4385 ( 
.A1(n_4324),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.C1(n_466),
.C2(n_467),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4225),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_L g4387 ( 
.A(n_4266),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4222),
.Y(n_4388)
);

NOR2xp33_ASAP7_75t_L g4389 ( 
.A(n_4217),
.B(n_465),
.Y(n_4389)
);

INVx5_ASAP7_75t_SL g4390 ( 
.A(n_4318),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4222),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4239),
.Y(n_4392)
);

INVx4_ASAP7_75t_L g4393 ( 
.A(n_4318),
.Y(n_4393)
);

OAI22xp33_ASAP7_75t_L g4394 ( 
.A1(n_4245),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_4394)
);

OAI21xp33_ASAP7_75t_L g4395 ( 
.A1(n_4203),
.A2(n_469),
.B(n_470),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_4310),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_L g4397 ( 
.A1(n_4271),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_4397)
);

AOI22xp33_ASAP7_75t_L g4398 ( 
.A1(n_4218),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_4398)
);

BUFx2_ASAP7_75t_L g4399 ( 
.A(n_4208),
.Y(n_4399)
);

AOI22xp33_ASAP7_75t_L g4400 ( 
.A1(n_4218),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4272),
.Y(n_4401)
);

BUFx12f_ASAP7_75t_L g4402 ( 
.A(n_4314),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_4362),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4247),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4253),
.Y(n_4405)
);

INVx3_ASAP7_75t_L g4406 ( 
.A(n_4230),
.Y(n_4406)
);

OAI22xp33_ASAP7_75t_L g4407 ( 
.A1(n_4245),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4257),
.Y(n_4408)
);

OAI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_4255),
.A2(n_482),
.B1(n_479),
.B2(n_480),
.Y(n_4409)
);

INVx2_ASAP7_75t_SL g4410 ( 
.A(n_4233),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4362),
.A2(n_483),
.B1(n_479),
.B2(n_480),
.Y(n_4411)
);

AOI22xp33_ASAP7_75t_L g4412 ( 
.A1(n_4203),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_4412)
);

OAI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_4315),
.A2(n_4252),
.B1(n_4244),
.B2(n_4269),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4264),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4252),
.A2(n_487),
.B1(n_484),
.B2(n_486),
.Y(n_4415)
);

OAI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4315),
.A2(n_486),
.B1(n_488),
.B2(n_489),
.Y(n_4416)
);

BUFx2_ASAP7_75t_L g4417 ( 
.A(n_4208),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4265),
.Y(n_4418)
);

HB1xp67_ASAP7_75t_L g4419 ( 
.A(n_4280),
.Y(n_4419)
);

BUFx3_ASAP7_75t_L g4420 ( 
.A(n_4266),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4310),
.Y(n_4421)
);

AOI22xp33_ASAP7_75t_SL g4422 ( 
.A1(n_4235),
.A2(n_697),
.B1(n_490),
.B2(n_491),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4206),
.Y(n_4423)
);

OAI21xp5_ASAP7_75t_SL g4424 ( 
.A1(n_4283),
.A2(n_489),
.B(n_490),
.Y(n_4424)
);

AOI22xp5_ASAP7_75t_L g4425 ( 
.A1(n_4336),
.A2(n_491),
.B1(n_492),
.B2(n_493),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4206),
.Y(n_4426)
);

OAI21xp5_ASAP7_75t_SL g4427 ( 
.A1(n_4283),
.A2(n_493),
.B(n_494),
.Y(n_4427)
);

AOI22xp33_ASAP7_75t_SL g4428 ( 
.A1(n_4348),
.A2(n_696),
.B1(n_495),
.B2(n_496),
.Y(n_4428)
);

INVxp67_ASAP7_75t_L g4429 ( 
.A(n_4355),
.Y(n_4429)
);

BUFx2_ASAP7_75t_L g4430 ( 
.A(n_4208),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_4212),
.A2(n_494),
.B1(n_497),
.B2(n_498),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4338),
.B(n_499),
.Y(n_4432)
);

AOI22xp33_ASAP7_75t_L g4433 ( 
.A1(n_4212),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_4433)
);

AOI22xp33_ASAP7_75t_L g4434 ( 
.A1(n_4336),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4292),
.B(n_502),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4299),
.Y(n_4436)
);

OAI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4349),
.A2(n_505),
.B1(n_507),
.B2(n_508),
.Y(n_4437)
);

INVx3_ASAP7_75t_L g4438 ( 
.A(n_4233),
.Y(n_4438)
);

AND2x2_ASAP7_75t_L g4439 ( 
.A(n_4285),
.B(n_505),
.Y(n_4439)
);

BUFx6f_ASAP7_75t_L g4440 ( 
.A(n_4266),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4238),
.B(n_507),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4299),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_L g4443 ( 
.A1(n_4352),
.A2(n_510),
.B1(n_511),
.B2(n_513),
.Y(n_4443)
);

OAI22xp5_ASAP7_75t_L g4444 ( 
.A1(n_4244),
.A2(n_4347),
.B1(n_4349),
.B2(n_4279),
.Y(n_4444)
);

AOI22xp33_ASAP7_75t_L g4445 ( 
.A1(n_4352),
.A2(n_511),
.B1(n_513),
.B2(n_514),
.Y(n_4445)
);

OAI22xp5_ASAP7_75t_L g4446 ( 
.A1(n_4282),
.A2(n_4301),
.B1(n_4318),
.B2(n_4350),
.Y(n_4446)
);

AND2x2_ASAP7_75t_L g4447 ( 
.A(n_4358),
.B(n_514),
.Y(n_4447)
);

AOI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_4213),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4301),
.B(n_515),
.Y(n_4449)
);

AOI22xp33_ASAP7_75t_L g4450 ( 
.A1(n_4213),
.A2(n_516),
.B1(n_517),
.B2(n_519),
.Y(n_4450)
);

OR2x2_ASAP7_75t_L g4451 ( 
.A(n_4201),
.B(n_519),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_L g4452 ( 
.A1(n_4361),
.A2(n_4334),
.B1(n_4288),
.B2(n_4357),
.Y(n_4452)
);

AOI22xp33_ASAP7_75t_SL g4453 ( 
.A1(n_4361),
.A2(n_696),
.B1(n_521),
.B2(n_522),
.Y(n_4453)
);

AOI22xp33_ASAP7_75t_L g4454 ( 
.A1(n_4334),
.A2(n_520),
.B1(n_521),
.B2(n_524),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_4243),
.B(n_525),
.Y(n_4455)
);

BUFx3_ASAP7_75t_L g4456 ( 
.A(n_4290),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4223),
.Y(n_4457)
);

AOI22xp33_ASAP7_75t_L g4458 ( 
.A1(n_4288),
.A2(n_4357),
.B1(n_4333),
.B2(n_4277),
.Y(n_4458)
);

CKINVDCx5p33_ASAP7_75t_R g4459 ( 
.A(n_4273),
.Y(n_4459)
);

OAI21xp5_ASAP7_75t_SL g4460 ( 
.A1(n_4249),
.A2(n_525),
.B(n_526),
.Y(n_4460)
);

AOI22xp33_ASAP7_75t_L g4461 ( 
.A1(n_4333),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.Y(n_4461)
);

AND2x4_ASAP7_75t_SL g4462 ( 
.A(n_4233),
.B(n_527),
.Y(n_4462)
);

OAI21xp5_ASAP7_75t_L g4463 ( 
.A1(n_4306),
.A2(n_528),
.B(n_529),
.Y(n_4463)
);

BUFx6f_ASAP7_75t_L g4464 ( 
.A(n_4322),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4223),
.Y(n_4465)
);

AOI22xp33_ASAP7_75t_L g4466 ( 
.A1(n_4277),
.A2(n_530),
.B1(n_531),
.B2(n_532),
.Y(n_4466)
);

AOI22xp33_ASAP7_75t_L g4467 ( 
.A1(n_4241),
.A2(n_530),
.B1(n_531),
.B2(n_532),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4241),
.A2(n_533),
.B1(n_535),
.B2(n_536),
.Y(n_4468)
);

AOI22xp33_ASAP7_75t_SL g4469 ( 
.A1(n_4307),
.A2(n_693),
.B1(n_535),
.B2(n_537),
.Y(n_4469)
);

INVx2_ASAP7_75t_SL g4470 ( 
.A(n_4340),
.Y(n_4470)
);

OAI222xp33_ASAP7_75t_L g4471 ( 
.A1(n_4345),
.A2(n_533),
.B1(n_537),
.B2(n_538),
.C1(n_539),
.C2(n_540),
.Y(n_4471)
);

OAI21xp5_ASAP7_75t_SL g4472 ( 
.A1(n_4329),
.A2(n_538),
.B(n_541),
.Y(n_4472)
);

OAI21xp33_ASAP7_75t_L g4473 ( 
.A1(n_4327),
.A2(n_541),
.B(n_542),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4251),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4254),
.Y(n_4475)
);

OAI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_4306),
.A2(n_542),
.B(n_544),
.Y(n_4476)
);

CKINVDCx11_ASAP7_75t_R g4477 ( 
.A(n_4305),
.Y(n_4477)
);

CKINVDCx20_ASAP7_75t_R g4478 ( 
.A(n_4325),
.Y(n_4478)
);

AOI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4226),
.A2(n_544),
.B1(n_545),
.B2(n_546),
.Y(n_4479)
);

BUFx6f_ASAP7_75t_L g4480 ( 
.A(n_4322),
.Y(n_4480)
);

AOI22xp33_ASAP7_75t_L g4481 ( 
.A1(n_4270),
.A2(n_4298),
.B1(n_4321),
.B2(n_4328),
.Y(n_4481)
);

INVx3_ASAP7_75t_L g4482 ( 
.A(n_4287),
.Y(n_4482)
);

AOI22xp33_ASAP7_75t_L g4483 ( 
.A1(n_4330),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4254),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4289),
.Y(n_4485)
);

AOI22xp33_ASAP7_75t_L g4486 ( 
.A1(n_4330),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.Y(n_4486)
);

OAI22xp5_ASAP7_75t_L g4487 ( 
.A1(n_4220),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.Y(n_4487)
);

BUFx6f_ASAP7_75t_L g4488 ( 
.A(n_4312),
.Y(n_4488)
);

INVx3_ASAP7_75t_L g4489 ( 
.A(n_4287),
.Y(n_4489)
);

HB1xp67_ASAP7_75t_L g4490 ( 
.A(n_4280),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4289),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4296),
.Y(n_4492)
);

CKINVDCx5p33_ASAP7_75t_R g4493 ( 
.A(n_4294),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4346),
.B(n_551),
.Y(n_4494)
);

OR2x2_ASAP7_75t_L g4495 ( 
.A(n_4215),
.B(n_552),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4326),
.B(n_4335),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4296),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4284),
.Y(n_4498)
);

OAI22xp5_ASAP7_75t_SL g4499 ( 
.A1(n_4234),
.A2(n_553),
.B1(n_554),
.B2(n_555),
.Y(n_4499)
);

AOI22xp33_ASAP7_75t_SL g4500 ( 
.A1(n_4355),
.A2(n_553),
.B1(n_554),
.B2(n_556),
.Y(n_4500)
);

AOI22xp33_ASAP7_75t_L g4501 ( 
.A1(n_4339),
.A2(n_556),
.B1(n_557),
.B2(n_558),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4337),
.B(n_558),
.Y(n_4502)
);

BUFx6f_ASAP7_75t_L g4503 ( 
.A(n_4340),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4311),
.Y(n_4504)
);

NOR2x1_ASAP7_75t_SL g4505 ( 
.A(n_4237),
.B(n_559),
.Y(n_4505)
);

OAI22xp5_ASAP7_75t_L g4506 ( 
.A1(n_4327),
.A2(n_559),
.B1(n_560),
.B2(n_561),
.Y(n_4506)
);

HB1xp67_ASAP7_75t_L g4507 ( 
.A(n_4202),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4311),
.B(n_560),
.Y(n_4508)
);

OAI22xp5_ASAP7_75t_L g4509 ( 
.A1(n_4344),
.A2(n_561),
.B1(n_562),
.B2(n_563),
.Y(n_4509)
);

CKINVDCx5p33_ASAP7_75t_R g4510 ( 
.A(n_4340),
.Y(n_4510)
);

AOI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_4339),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4511)
);

BUFx2_ASAP7_75t_L g4512 ( 
.A(n_4281),
.Y(n_4512)
);

INVx1_ASAP7_75t_SL g4513 ( 
.A(n_4215),
.Y(n_4513)
);

AOI22xp33_ASAP7_75t_L g4514 ( 
.A1(n_4262),
.A2(n_565),
.B1(n_567),
.B2(n_568),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4232),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4275),
.Y(n_4516)
);

OAI21xp5_ASAP7_75t_L g4517 ( 
.A1(n_4268),
.A2(n_567),
.B(n_568),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4276),
.Y(n_4518)
);

BUFx3_ASAP7_75t_L g4519 ( 
.A(n_4331),
.Y(n_4519)
);

OAI21xp5_ASAP7_75t_SL g4520 ( 
.A1(n_4356),
.A2(n_569),
.B(n_570),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4507),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4503),
.Y(n_4522)
);

OA21x2_ASAP7_75t_L g4523 ( 
.A1(n_4485),
.A2(n_4240),
.B(n_4297),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4366),
.B(n_4302),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4368),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4370),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4503),
.Y(n_4527)
);

INVx2_ASAP7_75t_SL g4528 ( 
.A(n_4503),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4399),
.B(n_4313),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_4393),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4372),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4417),
.B(n_4319),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4393),
.Y(n_4533)
);

BUFx2_ASAP7_75t_L g4534 ( 
.A(n_4402),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_4488),
.Y(n_4535)
);

OA21x2_ASAP7_75t_L g4536 ( 
.A1(n_4491),
.A2(n_4300),
.B(n_4304),
.Y(n_4536)
);

INVx2_ASAP7_75t_SL g4537 ( 
.A(n_4420),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4373),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4377),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4363),
.B(n_4274),
.Y(n_4540)
);

BUFx5_ASAP7_75t_L g4541 ( 
.A(n_4475),
.Y(n_4541)
);

INVx2_ASAP7_75t_L g4542 ( 
.A(n_4488),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4452),
.B(n_4274),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4386),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4379),
.A2(n_4200),
.B(n_4278),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4430),
.B(n_4323),
.Y(n_4546)
);

AO21x2_ASAP7_75t_L g4547 ( 
.A1(n_4449),
.A2(n_4303),
.B(n_4200),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_4488),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_4396),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4421),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4482),
.B(n_4198),
.Y(n_4551)
);

NAND2x1p5_ASAP7_75t_L g4552 ( 
.A(n_4464),
.B(n_4250),
.Y(n_4552)
);

AOI22xp33_ASAP7_75t_SL g4553 ( 
.A1(n_4379),
.A2(n_4286),
.B1(n_4198),
.B2(n_4356),
.Y(n_4553)
);

OR2x6_ASAP7_75t_L g4554 ( 
.A(n_4520),
.B(n_4317),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4482),
.B(n_4308),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4489),
.B(n_4316),
.Y(n_4556)
);

AO21x2_ASAP7_75t_L g4557 ( 
.A1(n_4455),
.A2(n_4286),
.B(n_4278),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4392),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4401),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4453),
.B(n_4256),
.Y(n_4560)
);

INVx2_ASAP7_75t_L g4561 ( 
.A(n_4384),
.Y(n_4561)
);

BUFx4f_ASAP7_75t_L g4562 ( 
.A(n_4387),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4404),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4405),
.Y(n_4564)
);

BUFx3_ASAP7_75t_L g4565 ( 
.A(n_4478),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4489),
.B(n_4316),
.Y(n_4566)
);

INVx2_ASAP7_75t_SL g4567 ( 
.A(n_4387),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4408),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4504),
.B(n_4316),
.Y(n_4569)
);

INVx2_ASAP7_75t_SL g4570 ( 
.A(n_4387),
.Y(n_4570)
);

INVx3_ASAP7_75t_L g4571 ( 
.A(n_4390),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4419),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4365),
.Y(n_4573)
);

INVxp67_ASAP7_75t_L g4574 ( 
.A(n_4505),
.Y(n_4574)
);

BUFx2_ASAP7_75t_L g4575 ( 
.A(n_4512),
.Y(n_4575)
);

OR2x2_ASAP7_75t_L g4576 ( 
.A(n_4429),
.B(n_4246),
.Y(n_4576)
);

HB1xp67_ASAP7_75t_L g4577 ( 
.A(n_4490),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4414),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4496),
.Y(n_4579)
);

AND2x2_ASAP7_75t_L g4580 ( 
.A(n_4388),
.B(n_4209),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4391),
.B(n_4214),
.Y(n_4581)
);

AOI21x1_ASAP7_75t_L g4582 ( 
.A1(n_4375),
.A2(n_4259),
.B(n_4256),
.Y(n_4582)
);

NAND2x1_ASAP7_75t_L g4583 ( 
.A(n_4436),
.B(n_4228),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4371),
.B(n_4242),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4418),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4464),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4498),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4516),
.Y(n_4588)
);

HB1xp67_ASAP7_75t_L g4589 ( 
.A(n_4518),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4442),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4458),
.B(n_4263),
.Y(n_4591)
);

AO21x2_ASAP7_75t_L g4592 ( 
.A1(n_4484),
.A2(n_4263),
.B(n_4207),
.Y(n_4592)
);

INVx3_ASAP7_75t_L g4593 ( 
.A(n_4390),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4371),
.B(n_4248),
.Y(n_4594)
);

INVx6_ASAP7_75t_L g4595 ( 
.A(n_4440),
.Y(n_4595)
);

OR2x6_ASAP7_75t_L g4596 ( 
.A(n_4520),
.B(n_4444),
.Y(n_4596)
);

OA21x2_ASAP7_75t_L g4597 ( 
.A1(n_4492),
.A2(n_4221),
.B(n_4295),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4381),
.B(n_4406),
.Y(n_4598)
);

AND2x4_ASAP7_75t_L g4599 ( 
.A(n_4470),
.B(n_4381),
.Y(n_4599)
);

BUFx3_ASAP7_75t_L g4600 ( 
.A(n_4477),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4464),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4480),
.Y(n_4602)
);

INVx2_ASAP7_75t_SL g4603 ( 
.A(n_4440),
.Y(n_4603)
);

BUFx3_ASAP7_75t_L g4604 ( 
.A(n_4456),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4480),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4480),
.Y(n_4606)
);

OA21x2_ASAP7_75t_L g4607 ( 
.A1(n_4497),
.A2(n_4258),
.B(n_4224),
.Y(n_4607)
);

AND2x2_ASAP7_75t_L g4608 ( 
.A(n_4406),
.B(n_4309),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4423),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4441),
.B(n_4444),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4438),
.B(n_4341),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4426),
.Y(n_4612)
);

NOR2xp33_ASAP7_75t_L g4613 ( 
.A(n_4440),
.B(n_4359),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4438),
.Y(n_4614)
);

OR2x2_ASAP7_75t_L g4615 ( 
.A(n_4474),
.B(n_4236),
.Y(n_4615)
);

OR2x6_ASAP7_75t_L g4616 ( 
.A(n_4463),
.B(n_4342),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4378),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4495),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4515),
.Y(n_4619)
);

AO21x2_ASAP7_75t_L g4620 ( 
.A1(n_4375),
.A2(n_4332),
.B(n_4353),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4410),
.B(n_4351),
.Y(n_4621)
);

HB1xp67_ASAP7_75t_L g4622 ( 
.A(n_4457),
.Y(n_4622)
);

HB1xp67_ASAP7_75t_L g4623 ( 
.A(n_4465),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4432),
.Y(n_4624)
);

OA21x2_ASAP7_75t_L g4625 ( 
.A1(n_4431),
.A2(n_4360),
.B(n_4331),
.Y(n_4625)
);

AO21x2_ASAP7_75t_L g4626 ( 
.A1(n_4468),
.A2(n_4261),
.B(n_4236),
.Y(n_4626)
);

INVx3_ASAP7_75t_L g4627 ( 
.A(n_4390),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4513),
.B(n_4261),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4519),
.Y(n_4629)
);

HB1xp67_ASAP7_75t_L g4630 ( 
.A(n_4451),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4508),
.Y(n_4631)
);

AOI22xp33_ASAP7_75t_L g4632 ( 
.A1(n_4413),
.A2(n_4395),
.B1(n_4364),
.B2(n_4446),
.Y(n_4632)
);

INVx3_ASAP7_75t_L g4633 ( 
.A(n_4510),
.Y(n_4633)
);

INVx3_ASAP7_75t_L g4634 ( 
.A(n_4493),
.Y(n_4634)
);

OAI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4433),
.A2(n_4261),
.B1(n_4236),
.B2(n_572),
.Y(n_4635)
);

AOI22xp33_ASAP7_75t_L g4636 ( 
.A1(n_4413),
.A2(n_569),
.B1(n_571),
.B2(n_573),
.Y(n_4636)
);

BUFx3_ASAP7_75t_L g4637 ( 
.A(n_4376),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4435),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4374),
.B(n_571),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4439),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4494),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4513),
.B(n_575),
.Y(n_4642)
);

HB1xp67_ASAP7_75t_L g4643 ( 
.A(n_4446),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4447),
.Y(n_4644)
);

HB1xp67_ASAP7_75t_L g4645 ( 
.A(n_4517),
.Y(n_4645)
);

CKINVDCx11_ASAP7_75t_R g4646 ( 
.A(n_4409),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4481),
.B(n_575),
.Y(n_4647)
);

AND2x4_ASAP7_75t_L g4648 ( 
.A(n_4517),
.B(n_576),
.Y(n_4648)
);

AO21x2_ASAP7_75t_L g4649 ( 
.A1(n_4471),
.A2(n_576),
.B(n_577),
.Y(n_4649)
);

INVx5_ASAP7_75t_L g4650 ( 
.A(n_4502),
.Y(n_4650)
);

BUFx3_ASAP7_75t_L g4651 ( 
.A(n_4459),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4437),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4506),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4364),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4462),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_4389),
.Y(n_4656)
);

HB1xp67_ASAP7_75t_L g4657 ( 
.A(n_4463),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4473),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4398),
.B(n_578),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_SL g4660 ( 
.A(n_4383),
.B(n_578),
.Y(n_4660)
);

INVx3_ASAP7_75t_L g4661 ( 
.A(n_4422),
.Y(n_4661)
);

AND2x4_ASAP7_75t_L g4662 ( 
.A(n_4367),
.B(n_579),
.Y(n_4662)
);

INVx4_ASAP7_75t_L g4663 ( 
.A(n_4385),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4369),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4416),
.Y(n_4665)
);

BUFx3_ASAP7_75t_L g4666 ( 
.A(n_4499),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4416),
.Y(n_4667)
);

NOR2x1_ASAP7_75t_SL g4668 ( 
.A(n_4554),
.B(n_4460),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4575),
.B(n_4400),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4575),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4633),
.B(n_4443),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4572),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4633),
.B(n_4445),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4633),
.B(n_4479),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4577),
.Y(n_4675)
);

OR2x2_ASAP7_75t_L g4676 ( 
.A(n_4667),
.B(n_4467),
.Y(n_4676)
);

NOR2x1_ASAP7_75t_L g4677 ( 
.A(n_4600),
.B(n_4424),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4537),
.B(n_4476),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4521),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4541),
.Y(n_4680)
);

OR2x2_ASAP7_75t_L g4681 ( 
.A(n_4667),
.B(n_4454),
.Y(n_4681)
);

AND2x4_ASAP7_75t_L g4682 ( 
.A(n_4571),
.B(n_4476),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4662),
.B(n_4500),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4590),
.Y(n_4684)
);

INVx2_ASAP7_75t_SL g4685 ( 
.A(n_4600),
.Y(n_4685)
);

AND2x2_ASAP7_75t_L g4686 ( 
.A(n_4537),
.B(n_4403),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4571),
.B(n_4411),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4525),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4541),
.Y(n_4689)
);

CKINVDCx20_ASAP7_75t_R g4690 ( 
.A(n_4534),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4541),
.Y(n_4691)
);

OR2x2_ASAP7_75t_L g4692 ( 
.A(n_4645),
.B(n_4424),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4526),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4531),
.Y(n_4694)
);

INVx2_ASAP7_75t_L g4695 ( 
.A(n_4541),
.Y(n_4695)
);

BUFx2_ASAP7_75t_L g4696 ( 
.A(n_4534),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4541),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4571),
.B(n_4483),
.Y(n_4698)
);

OA21x2_ASAP7_75t_L g4699 ( 
.A1(n_4632),
.A2(n_4427),
.B(n_4472),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4538),
.Y(n_4700)
);

INVx5_ASAP7_75t_L g4701 ( 
.A(n_4595),
.Y(n_4701)
);

AND2x4_ASAP7_75t_L g4702 ( 
.A(n_4593),
.B(n_4425),
.Y(n_4702)
);

BUFx3_ASAP7_75t_L g4703 ( 
.A(n_4565),
.Y(n_4703)
);

AO21x2_ASAP7_75t_L g4704 ( 
.A1(n_4654),
.A2(n_4427),
.B(n_4409),
.Y(n_4704)
);

OA21x2_ASAP7_75t_L g4705 ( 
.A1(n_4545),
.A2(n_4472),
.B(n_4382),
.Y(n_4705)
);

OR2x2_ASAP7_75t_L g4706 ( 
.A(n_4643),
.B(n_4486),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4539),
.Y(n_4707)
);

INVx2_ASAP7_75t_SL g4708 ( 
.A(n_4595),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4544),
.Y(n_4709)
);

BUFx8_ASAP7_75t_SL g4710 ( 
.A(n_4565),
.Y(n_4710)
);

OR2x2_ASAP7_75t_L g4711 ( 
.A(n_4549),
.B(n_4501),
.Y(n_4711)
);

NOR2x1_ASAP7_75t_SL g4712 ( 
.A(n_4554),
.B(n_4460),
.Y(n_4712)
);

AND2x2_ASAP7_75t_SL g4713 ( 
.A(n_4663),
.B(n_4397),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4598),
.B(n_4511),
.Y(n_4714)
);

BUFx2_ASAP7_75t_L g4715 ( 
.A(n_4604),
.Y(n_4715)
);

AOI211xp5_ASAP7_75t_L g4716 ( 
.A1(n_4635),
.A2(n_4394),
.B(n_4407),
.C(n_4509),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4558),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4559),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4662),
.B(n_4380),
.Y(n_4719)
);

INVx2_ASAP7_75t_SL g4720 ( 
.A(n_4595),
.Y(n_4720)
);

AOI221xp5_ASAP7_75t_L g4721 ( 
.A1(n_4663),
.A2(n_4412),
.B1(n_4448),
.B2(n_4450),
.C(n_4415),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_4541),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4563),
.Y(n_4723)
);

HB1xp67_ASAP7_75t_L g4724 ( 
.A(n_4657),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4598),
.B(n_4428),
.Y(n_4725)
);

AOI221xp5_ASAP7_75t_L g4726 ( 
.A1(n_4663),
.A2(n_4469),
.B1(n_4434),
.B2(n_4487),
.C(n_4461),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4541),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4593),
.B(n_4466),
.Y(n_4728)
);

BUFx2_ASAP7_75t_L g4729 ( 
.A(n_4604),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4564),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4662),
.B(n_4385),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4650),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4593),
.B(n_4514),
.Y(n_4733)
);

INVx2_ASAP7_75t_L g4734 ( 
.A(n_4650),
.Y(n_4734)
);

INVxp67_ASAP7_75t_SL g4735 ( 
.A(n_4661),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4661),
.B(n_579),
.Y(n_4736)
);

AND2x4_ASAP7_75t_L g4737 ( 
.A(n_4627),
.B(n_580),
.Y(n_4737)
);

NOR2xp33_ASAP7_75t_L g4738 ( 
.A(n_4661),
.B(n_581),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4627),
.B(n_581),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4650),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4627),
.B(n_582),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4568),
.Y(n_4742)
);

BUFx3_ASAP7_75t_L g4743 ( 
.A(n_4637),
.Y(n_4743)
);

HB1xp67_ASAP7_75t_L g4744 ( 
.A(n_4596),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4578),
.Y(n_4745)
);

OR2x2_ASAP7_75t_L g4746 ( 
.A(n_4549),
.B(n_582),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4644),
.B(n_583),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4611),
.B(n_584),
.Y(n_4748)
);

OR2x2_ASAP7_75t_L g4749 ( 
.A(n_4550),
.B(n_4561),
.Y(n_4749)
);

HB1xp67_ASAP7_75t_L g4750 ( 
.A(n_4596),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4611),
.B(n_4532),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4532),
.B(n_584),
.Y(n_4752)
);

HB1xp67_ASAP7_75t_L g4753 ( 
.A(n_4596),
.Y(n_4753)
);

AND2x4_ASAP7_75t_L g4754 ( 
.A(n_4599),
.B(n_585),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4585),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4644),
.B(n_586),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4650),
.Y(n_4757)
);

HB1xp67_ASAP7_75t_L g4758 ( 
.A(n_4596),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4650),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4587),
.Y(n_4760)
);

INVxp67_ASAP7_75t_SL g4761 ( 
.A(n_4666),
.Y(n_4761)
);

INVx4_ASAP7_75t_L g4762 ( 
.A(n_4595),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4546),
.B(n_586),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4588),
.Y(n_4764)
);

AO21x2_ASAP7_75t_L g4765 ( 
.A1(n_4642),
.A2(n_587),
.B(n_588),
.Y(n_4765)
);

AOI33xp33_ASAP7_75t_L g4766 ( 
.A1(n_4553),
.A2(n_587),
.A3(n_589),
.B1(n_590),
.B2(n_591),
.B3(n_592),
.Y(n_4766)
);

INVx1_ASAP7_75t_SL g4767 ( 
.A(n_4637),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4630),
.Y(n_4768)
);

AO31x2_ASAP7_75t_L g4769 ( 
.A1(n_4664),
.A2(n_589),
.A3(n_590),
.B(n_591),
.Y(n_4769)
);

OAI21xp5_ASAP7_75t_SL g4770 ( 
.A1(n_4543),
.A2(n_592),
.B(n_593),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4550),
.Y(n_4771)
);

AOI22xp33_ASAP7_75t_SL g4772 ( 
.A1(n_4666),
.A2(n_691),
.B1(n_594),
.B2(n_595),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4642),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4583),
.Y(n_4774)
);

AND2x2_ASAP7_75t_L g4775 ( 
.A(n_4546),
.B(n_593),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4583),
.Y(n_4776)
);

INVx3_ASAP7_75t_L g4777 ( 
.A(n_4634),
.Y(n_4777)
);

OR2x2_ASAP7_75t_L g4778 ( 
.A(n_4561),
.B(n_594),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4567),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4567),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4641),
.B(n_595),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4641),
.B(n_596),
.Y(n_4782)
);

HB1xp67_ASAP7_75t_L g4783 ( 
.A(n_4696),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4690),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4670),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4715),
.B(n_4599),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4729),
.B(n_4599),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4670),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4690),
.Y(n_4789)
);

HB1xp67_ASAP7_75t_L g4790 ( 
.A(n_4732),
.Y(n_4790)
);

HB1xp67_ASAP7_75t_L g4791 ( 
.A(n_4732),
.Y(n_4791)
);

OR2x2_ASAP7_75t_L g4792 ( 
.A(n_4724),
.B(n_4704),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_4751),
.B(n_4530),
.Y(n_4793)
);

BUFx3_ASAP7_75t_L g4794 ( 
.A(n_4710),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4771),
.Y(n_4795)
);

OR2x2_ASAP7_75t_L g4796 ( 
.A(n_4724),
.B(n_4704),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4679),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4749),
.Y(n_4798)
);

HB1xp67_ASAP7_75t_L g4799 ( 
.A(n_4734),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4703),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4768),
.Y(n_4801)
);

OR2x2_ASAP7_75t_L g4802 ( 
.A(n_4692),
.B(n_4610),
.Y(n_4802)
);

INVx4_ASAP7_75t_L g4803 ( 
.A(n_4710),
.Y(n_4803)
);

OR2x2_ASAP7_75t_L g4804 ( 
.A(n_4735),
.B(n_4579),
.Y(n_4804)
);

AND2x2_ASAP7_75t_L g4805 ( 
.A(n_4777),
.B(n_4725),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4672),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4675),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4773),
.Y(n_4808)
);

INVx2_ASAP7_75t_L g4809 ( 
.A(n_4703),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4777),
.B(n_4530),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4746),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4743),
.Y(n_4812)
);

OR2x2_ASAP7_75t_L g4813 ( 
.A(n_4735),
.B(n_4626),
.Y(n_4813)
);

INVx1_ASAP7_75t_SL g4814 ( 
.A(n_4767),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4684),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4775),
.Y(n_4816)
);

OR2x2_ASAP7_75t_L g4817 ( 
.A(n_4676),
.B(n_4626),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4775),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4743),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_4761),
.B(n_4574),
.Y(n_4820)
);

INVxp67_ASAP7_75t_SL g4821 ( 
.A(n_4761),
.Y(n_4821)
);

OR2x2_ASAP7_75t_L g4822 ( 
.A(n_4744),
.B(n_4579),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4777),
.Y(n_4823)
);

INVx2_ASAP7_75t_SL g4824 ( 
.A(n_4701),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4774),
.Y(n_4825)
);

AND2x4_ASAP7_75t_L g4826 ( 
.A(n_4701),
.B(n_4528),
.Y(n_4826)
);

NAND2x1_ASAP7_75t_L g4827 ( 
.A(n_4762),
.B(n_4556),
.Y(n_4827)
);

INVx2_ASAP7_75t_L g4828 ( 
.A(n_4774),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4778),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_L g4830 ( 
.A(n_4725),
.B(n_4640),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4738),
.B(n_4640),
.Y(n_4831)
);

AND2x2_ASAP7_75t_L g4832 ( 
.A(n_4685),
.B(n_4533),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4734),
.Y(n_4833)
);

OR2x2_ASAP7_75t_L g4834 ( 
.A(n_4681),
.B(n_4626),
.Y(n_4834)
);

INVx3_ASAP7_75t_L g4835 ( 
.A(n_4762),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4685),
.B(n_4533),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4738),
.B(n_4631),
.Y(n_4837)
);

INVx2_ASAP7_75t_L g4838 ( 
.A(n_4776),
.Y(n_4838)
);

OR2x2_ASAP7_75t_L g4839 ( 
.A(n_4711),
.B(n_4573),
.Y(n_4839)
);

OR2x6_ASAP7_75t_L g4840 ( 
.A(n_4677),
.B(n_4744),
.Y(n_4840)
);

INVx2_ASAP7_75t_SL g4841 ( 
.A(n_4701),
.Y(n_4841)
);

HB1xp67_ASAP7_75t_L g4842 ( 
.A(n_4740),
.Y(n_4842)
);

OR2x2_ASAP7_75t_L g4843 ( 
.A(n_4706),
.B(n_4573),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_L g4844 ( 
.A(n_4713),
.B(n_4646),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4776),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4740),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4757),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4701),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4757),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4762),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4668),
.B(n_4570),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4766),
.B(n_4631),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4766),
.B(n_4665),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4712),
.B(n_4570),
.Y(n_4854)
);

INVxp67_ASAP7_75t_L g4855 ( 
.A(n_4750),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4674),
.B(n_4603),
.Y(n_4856)
);

HB1xp67_ASAP7_75t_L g4857 ( 
.A(n_4792),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4792),
.Y(n_4858)
);

OR2x2_ASAP7_75t_L g4859 ( 
.A(n_4796),
.B(n_4699),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4796),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4784),
.B(n_4678),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4821),
.B(n_4713),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4783),
.B(n_4699),
.Y(n_4863)
);

AND2x2_ASAP7_75t_L g4864 ( 
.A(n_4784),
.B(n_4714),
.Y(n_4864)
);

BUFx2_ASAP7_75t_L g4865 ( 
.A(n_4840),
.Y(n_4865)
);

HB1xp67_ASAP7_75t_L g4866 ( 
.A(n_4786),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4813),
.Y(n_4867)
);

AND2x2_ASAP7_75t_L g4868 ( 
.A(n_4789),
.B(n_4714),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4813),
.Y(n_4869)
);

INVx3_ASAP7_75t_L g4870 ( 
.A(n_4803),
.Y(n_4870)
);

NAND3xp33_ASAP7_75t_L g4871 ( 
.A(n_4844),
.B(n_4840),
.C(n_4753),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_4840),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4855),
.B(n_4699),
.Y(n_4873)
);

AND2x4_ASAP7_75t_L g4874 ( 
.A(n_4826),
.B(n_4786),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4789),
.B(n_4708),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4816),
.B(n_4731),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_SL g4877 ( 
.A(n_4814),
.B(n_4562),
.Y(n_4877)
);

HB1xp67_ASAP7_75t_L g4878 ( 
.A(n_4787),
.Y(n_4878)
);

AND2x2_ASAP7_75t_L g4879 ( 
.A(n_4787),
.B(n_4805),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4840),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4805),
.B(n_4708),
.Y(n_4881)
);

AND2x4_ASAP7_75t_L g4882 ( 
.A(n_4826),
.B(n_4794),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4817),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4804),
.Y(n_4884)
);

AND2x2_ASAP7_75t_L g4885 ( 
.A(n_4856),
.B(n_4720),
.Y(n_4885)
);

AND2x2_ASAP7_75t_L g4886 ( 
.A(n_4856),
.B(n_4720),
.Y(n_4886)
);

OR2x2_ASAP7_75t_L g4887 ( 
.A(n_4817),
.B(n_4750),
.Y(n_4887)
);

AND2x2_ASAP7_75t_L g4888 ( 
.A(n_4832),
.B(n_4753),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4790),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4791),
.Y(n_4890)
);

HB1xp67_ASAP7_75t_L g4891 ( 
.A(n_4823),
.Y(n_4891)
);

AND2x4_ASAP7_75t_L g4892 ( 
.A(n_4826),
.B(n_4759),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4799),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4842),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4834),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4785),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4788),
.Y(n_4897)
);

AND2x2_ASAP7_75t_L g4898 ( 
.A(n_4832),
.B(n_4758),
.Y(n_4898)
);

AND2x2_ASAP7_75t_L g4899 ( 
.A(n_4836),
.B(n_4758),
.Y(n_4899)
);

INVx2_ASAP7_75t_L g4900 ( 
.A(n_4834),
.Y(n_4900)
);

OR2x2_ASAP7_75t_L g4901 ( 
.A(n_4843),
.B(n_4759),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4836),
.B(n_4702),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4812),
.B(n_4702),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4822),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4812),
.B(n_4702),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4819),
.B(n_4851),
.Y(n_4906)
);

AND2x2_ASAP7_75t_SL g4907 ( 
.A(n_4844),
.B(n_4705),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4835),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4819),
.B(n_4698),
.Y(n_4909)
);

NOR2xp33_ASAP7_75t_L g4910 ( 
.A(n_4803),
.B(n_4634),
.Y(n_4910)
);

INVx2_ASAP7_75t_L g4911 ( 
.A(n_4835),
.Y(n_4911)
);

OR2x2_ASAP7_75t_L g4912 ( 
.A(n_4843),
.B(n_4779),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4851),
.B(n_4682),
.Y(n_4913)
);

NAND2xp33_ASAP7_75t_R g4914 ( 
.A(n_4820),
.B(n_4705),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4835),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4854),
.B(n_4682),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4823),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4902),
.B(n_4800),
.Y(n_4918)
);

INVxp67_ASAP7_75t_L g4919 ( 
.A(n_4902),
.Y(n_4919)
);

HB1xp67_ASAP7_75t_L g4920 ( 
.A(n_4866),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4878),
.Y(n_4921)
);

BUFx2_ASAP7_75t_L g4922 ( 
.A(n_4857),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4891),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4857),
.Y(n_4924)
);

AOI22xp33_ASAP7_75t_L g4925 ( 
.A1(n_4907),
.A2(n_4646),
.B1(n_4705),
.B2(n_4794),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4912),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4879),
.B(n_4800),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4879),
.B(n_4803),
.Y(n_4928)
);

INVx4_ASAP7_75t_L g4929 ( 
.A(n_4870),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4912),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4885),
.B(n_4809),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4901),
.Y(n_4932)
);

AND2x4_ASAP7_75t_L g4933 ( 
.A(n_4874),
.B(n_4824),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4901),
.Y(n_4934)
);

INVx1_ASAP7_75t_SL g4935 ( 
.A(n_4888),
.Y(n_4935)
);

HB1xp67_ASAP7_75t_L g4936 ( 
.A(n_4874),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4888),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4898),
.Y(n_4938)
);

INVx2_ASAP7_75t_L g4939 ( 
.A(n_4860),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4885),
.B(n_4886),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4898),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4860),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4886),
.B(n_4793),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4899),
.B(n_4809),
.Y(n_4944)
);

NOR2xp33_ASAP7_75t_L g4945 ( 
.A(n_4870),
.B(n_4853),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4899),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4882),
.B(n_4793),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4860),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4881),
.B(n_4810),
.Y(n_4949)
);

AND2x4_ASAP7_75t_L g4950 ( 
.A(n_4874),
.B(n_4824),
.Y(n_4950)
);

OR2x2_ASAP7_75t_L g4951 ( 
.A(n_4859),
.B(n_4830),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4874),
.Y(n_4952)
);

AND2x2_ASAP7_75t_L g4953 ( 
.A(n_4882),
.B(n_4854),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4889),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4881),
.B(n_4810),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4889),
.Y(n_4956)
);

OR2x2_ASAP7_75t_L g4957 ( 
.A(n_4859),
.B(n_4839),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4882),
.B(n_4779),
.Y(n_4958)
);

INVx1_ASAP7_75t_SL g4959 ( 
.A(n_4913),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4882),
.B(n_4780),
.Y(n_4960)
);

HB1xp67_ASAP7_75t_L g4961 ( 
.A(n_4870),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4890),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4913),
.B(n_4780),
.Y(n_4963)
);

INVx2_ASAP7_75t_SL g4964 ( 
.A(n_4892),
.Y(n_4964)
);

NOR2xp33_ASAP7_75t_L g4965 ( 
.A(n_4870),
.B(n_4818),
.Y(n_4965)
);

AOI22xp33_ASAP7_75t_L g4966 ( 
.A1(n_4907),
.A2(n_4802),
.B1(n_4669),
.B2(n_4721),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4916),
.B(n_4903),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4903),
.B(n_4754),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4890),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4893),
.Y(n_4970)
);

HB1xp67_ASAP7_75t_L g4971 ( 
.A(n_4865),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4893),
.Y(n_4972)
);

INVx2_ASAP7_75t_L g4973 ( 
.A(n_4865),
.Y(n_4973)
);

OR2x2_ASAP7_75t_L g4974 ( 
.A(n_4863),
.B(n_4839),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_SL g4975 ( 
.A(n_4928),
.B(n_4907),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4922),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4928),
.B(n_4916),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4940),
.B(n_4905),
.Y(n_4978)
);

INVxp67_ASAP7_75t_L g4979 ( 
.A(n_4940),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4947),
.B(n_4905),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4922),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4936),
.Y(n_4982)
);

HB1xp67_ASAP7_75t_L g4983 ( 
.A(n_4964),
.Y(n_4983)
);

INVx2_ASAP7_75t_L g4984 ( 
.A(n_4964),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4947),
.B(n_4906),
.Y(n_4985)
);

AND2x2_ASAP7_75t_L g4986 ( 
.A(n_4953),
.B(n_4906),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4953),
.B(n_4864),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4957),
.B(n_4863),
.Y(n_4988)
);

OR2x2_ASAP7_75t_L g4989 ( 
.A(n_4957),
.B(n_4873),
.Y(n_4989)
);

NOR2x1_ASAP7_75t_L g4990 ( 
.A(n_4924),
.B(n_4858),
.Y(n_4990)
);

AND2x2_ASAP7_75t_L g4991 ( 
.A(n_4943),
.B(n_4864),
.Y(n_4991)
);

OR2x2_ASAP7_75t_L g4992 ( 
.A(n_4935),
.B(n_4873),
.Y(n_4992)
);

INVx2_ASAP7_75t_L g4993 ( 
.A(n_4933),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4943),
.B(n_4868),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4933),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4961),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4967),
.B(n_4868),
.Y(n_4997)
);

NOR2x1p5_ASAP7_75t_L g4998 ( 
.A(n_4944),
.B(n_4862),
.Y(n_4998)
);

INVx1_ASAP7_75t_SL g4999 ( 
.A(n_4967),
.Y(n_4999)
);

HB1xp67_ASAP7_75t_L g5000 ( 
.A(n_4933),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4958),
.B(n_4875),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_4950),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4958),
.B(n_4875),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4960),
.B(n_4909),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4924),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_4950),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4939),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4939),
.Y(n_5008)
);

HB1xp67_ASAP7_75t_L g5009 ( 
.A(n_4950),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4974),
.B(n_4862),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4942),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4942),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4948),
.Y(n_5013)
);

AND2x2_ASAP7_75t_L g5014 ( 
.A(n_4960),
.B(n_4909),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_SL g5015 ( 
.A(n_4925),
.B(n_4682),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4959),
.B(n_4861),
.Y(n_5016)
);

AND2x2_ASAP7_75t_L g5017 ( 
.A(n_4963),
.B(n_4861),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4963),
.B(n_4892),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4948),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4920),
.Y(n_5020)
);

HB1xp67_ASAP7_75t_L g5021 ( 
.A(n_4952),
.Y(n_5021)
);

HB1xp67_ASAP7_75t_L g5022 ( 
.A(n_4952),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4937),
.B(n_4910),
.Y(n_5023)
);

NOR2xp33_ASAP7_75t_SL g5024 ( 
.A(n_4919),
.B(n_4562),
.Y(n_5024)
);

BUFx3_ASAP7_75t_L g5025 ( 
.A(n_4973),
.Y(n_5025)
);

INVx1_ASAP7_75t_SL g5026 ( 
.A(n_5003),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4997),
.B(n_4938),
.Y(n_5027)
);

HB1xp67_ASAP7_75t_L g5028 ( 
.A(n_4990),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_4997),
.B(n_4941),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_5000),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_5009),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4983),
.Y(n_5032)
);

INVxp67_ASAP7_75t_SL g5033 ( 
.A(n_4990),
.Y(n_5033)
);

AND2x2_ASAP7_75t_L g5034 ( 
.A(n_5003),
.B(n_4946),
.Y(n_5034)
);

AND2x2_ASAP7_75t_L g5035 ( 
.A(n_4987),
.B(n_4904),
.Y(n_5035)
);

AND2x2_ASAP7_75t_L g5036 ( 
.A(n_4987),
.B(n_4904),
.Y(n_5036)
);

HB1xp67_ASAP7_75t_L g5037 ( 
.A(n_4993),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_5017),
.B(n_4892),
.Y(n_5038)
);

HB1xp67_ASAP7_75t_L g5039 ( 
.A(n_4993),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_5017),
.B(n_4892),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4977),
.B(n_4949),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4995),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4977),
.B(n_4955),
.Y(n_5043)
);

INVx2_ASAP7_75t_L g5044 ( 
.A(n_4995),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_4986),
.B(n_4966),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4986),
.B(n_4921),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4991),
.B(n_4931),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_5002),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_5004),
.B(n_4926),
.Y(n_5049)
);

AND2x4_ASAP7_75t_L g5050 ( 
.A(n_5002),
.B(n_4929),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_5006),
.Y(n_5051)
);

BUFx2_ASAP7_75t_L g5052 ( 
.A(n_5006),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_5025),
.Y(n_5053)
);

NOR2x1_ASAP7_75t_SL g5054 ( 
.A(n_5004),
.B(n_4765),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_5014),
.B(n_4978),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_5014),
.B(n_4884),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_5025),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_5025),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_5021),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_5022),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_4978),
.B(n_4991),
.Y(n_5061)
);

AOI22xp33_ASAP7_75t_L g5062 ( 
.A1(n_5015),
.A2(n_4871),
.B1(n_4945),
.B2(n_4998),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_SL g5063 ( 
.A(n_4989),
.B(n_4858),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4981),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4994),
.B(n_4930),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4981),
.Y(n_5066)
);

OR2x2_ASAP7_75t_L g5067 ( 
.A(n_4999),
.B(n_4927),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_SL g5068 ( 
.A(n_4989),
.B(n_4988),
.Y(n_5068)
);

AND2x2_ASAP7_75t_SL g5069 ( 
.A(n_5010),
.B(n_4945),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_4994),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_4979),
.B(n_4850),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4976),
.Y(n_5072)
);

AND2x2_ASAP7_75t_L g5073 ( 
.A(n_5023),
.B(n_4918),
.Y(n_5073)
);

INVx1_ASAP7_75t_SL g5074 ( 
.A(n_5018),
.Y(n_5074)
);

OR2x2_ASAP7_75t_L g5075 ( 
.A(n_5001),
.B(n_4951),
.Y(n_5075)
);

NAND2x1_ASAP7_75t_L g5076 ( 
.A(n_4976),
.B(n_4929),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_5020),
.B(n_4850),
.Y(n_5077)
);

NOR2x1_ASAP7_75t_L g5078 ( 
.A(n_4988),
.B(n_4929),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_5028),
.Y(n_5079)
);

OR2x2_ASAP7_75t_L g5080 ( 
.A(n_5026),
.B(n_4985),
.Y(n_5080)
);

OR2x2_ASAP7_75t_L g5081 ( 
.A(n_5061),
.B(n_5055),
.Y(n_5081)
);

INVxp67_ASAP7_75t_L g5082 ( 
.A(n_5054),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_5033),
.B(n_4971),
.Y(n_5083)
);

AND2x2_ASAP7_75t_L g5084 ( 
.A(n_5047),
.B(n_5023),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_5041),
.B(n_5043),
.Y(n_5085)
);

OR2x2_ASAP7_75t_L g5086 ( 
.A(n_5038),
.B(n_4980),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_5027),
.B(n_5016),
.Y(n_5087)
);

HB1xp67_ASAP7_75t_L g5088 ( 
.A(n_5028),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_5033),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_5037),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_5037),
.Y(n_5091)
);

OR2x2_ASAP7_75t_L g5092 ( 
.A(n_5040),
.B(n_4992),
.Y(n_5092)
);

HB1xp67_ASAP7_75t_L g5093 ( 
.A(n_5039),
.Y(n_5093)
);

OR2x2_ASAP7_75t_L g5094 ( 
.A(n_5070),
.B(n_4992),
.Y(n_5094)
);

AOI21xp33_ASAP7_75t_L g5095 ( 
.A1(n_5068),
.A2(n_4914),
.B(n_5010),
.Y(n_5095)
);

OR2x2_ASAP7_75t_L g5096 ( 
.A(n_5065),
.B(n_4951),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5039),
.Y(n_5097)
);

OR2x2_ASAP7_75t_L g5098 ( 
.A(n_5030),
.B(n_4975),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5078),
.Y(n_5099)
);

AND2x2_ASAP7_75t_L g5100 ( 
.A(n_5029),
.B(n_4968),
.Y(n_5100)
);

INVx3_ASAP7_75t_L g5101 ( 
.A(n_5050),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_5073),
.B(n_4998),
.Y(n_5102)
);

OR2x2_ASAP7_75t_L g5103 ( 
.A(n_5031),
.B(n_4974),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5050),
.Y(n_5104)
);

INVx2_ASAP7_75t_L g5105 ( 
.A(n_5050),
.Y(n_5105)
);

OR2x2_ASAP7_75t_L g5106 ( 
.A(n_5049),
.B(n_4982),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_5076),
.Y(n_5107)
);

NAND3xp33_ASAP7_75t_SL g5108 ( 
.A(n_5062),
.B(n_4871),
.C(n_5024),
.Y(n_5108)
);

INVx1_ASAP7_75t_SL g5109 ( 
.A(n_5069),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_5069),
.B(n_4982),
.Y(n_5110)
);

INVx1_ASAP7_75t_SL g5111 ( 
.A(n_5035),
.Y(n_5111)
);

NOR2xp33_ASAP7_75t_L g5112 ( 
.A(n_5074),
.B(n_4877),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_5035),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_5036),
.Y(n_5114)
);

AND2x2_ASAP7_75t_L g5115 ( 
.A(n_5046),
.B(n_4811),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5053),
.B(n_4973),
.Y(n_5116)
);

OAI322xp33_ASAP7_75t_L g5117 ( 
.A1(n_5068),
.A2(n_4880),
.A3(n_4872),
.B1(n_4894),
.B2(n_5020),
.C1(n_4887),
.C2(n_4956),
.Y(n_5117)
);

INVx2_ASAP7_75t_SL g5118 ( 
.A(n_5056),
.Y(n_5118)
);

OR2x2_ASAP7_75t_L g5119 ( 
.A(n_5067),
.B(n_4837),
.Y(n_5119)
);

AND2x2_ASAP7_75t_L g5120 ( 
.A(n_5046),
.B(n_4829),
.Y(n_5120)
);

INVx2_ASAP7_75t_SL g5121 ( 
.A(n_5056),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_5036),
.Y(n_5122)
);

NAND2xp5_ASAP7_75t_L g5123 ( 
.A(n_5034),
.B(n_4932),
.Y(n_5123)
);

OR2x2_ASAP7_75t_L g5124 ( 
.A(n_5057),
.B(n_4876),
.Y(n_5124)
);

HB1xp67_ASAP7_75t_L g5125 ( 
.A(n_5058),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_5034),
.B(n_4984),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_5032),
.B(n_4884),
.Y(n_5127)
);

AND2x2_ASAP7_75t_L g5128 ( 
.A(n_5052),
.B(n_4634),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_5101),
.Y(n_5129)
);

AND2x2_ASAP7_75t_L g5130 ( 
.A(n_5128),
.B(n_4934),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_5101),
.Y(n_5131)
);

BUFx2_ASAP7_75t_L g5132 ( 
.A(n_5118),
.Y(n_5132)
);

NOR2xp67_ASAP7_75t_L g5133 ( 
.A(n_5121),
.B(n_4872),
.Y(n_5133)
);

OR2x2_ASAP7_75t_L g5134 ( 
.A(n_5111),
.B(n_5045),
.Y(n_5134)
);

NAND2x1p5_ASAP7_75t_L g5135 ( 
.A(n_5111),
.B(n_5104),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_5093),
.B(n_4984),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_5126),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_5126),
.Y(n_5138)
);

OR2x2_ASAP7_75t_L g5139 ( 
.A(n_5113),
.B(n_4876),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_5110),
.Y(n_5140)
);

AND2x2_ASAP7_75t_L g5141 ( 
.A(n_5084),
.B(n_4894),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_5095),
.B(n_4872),
.Y(n_5142)
);

OR2x2_ASAP7_75t_L g5143 ( 
.A(n_5114),
.B(n_4831),
.Y(n_5143)
);

OR2x2_ASAP7_75t_L g5144 ( 
.A(n_5122),
.B(n_4887),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_5095),
.B(n_4880),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_5110),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_5085),
.B(n_4923),
.Y(n_5147)
);

INVx3_ASAP7_75t_L g5148 ( 
.A(n_5105),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_5115),
.Y(n_5149)
);

AND2x2_ASAP7_75t_L g5150 ( 
.A(n_5087),
.B(n_4880),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_5088),
.Y(n_5151)
);

AND2x2_ASAP7_75t_L g5152 ( 
.A(n_5100),
.B(n_5044),
.Y(n_5152)
);

AND2x4_ASAP7_75t_L g5153 ( 
.A(n_5120),
.B(n_5044),
.Y(n_5153)
);

AND2x2_ASAP7_75t_L g5154 ( 
.A(n_5102),
.B(n_5059),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_5090),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_5091),
.Y(n_5156)
);

OAI221xp5_ASAP7_75t_L g5157 ( 
.A1(n_5109),
.A2(n_5062),
.B1(n_5063),
.B2(n_4736),
.C(n_5005),
.Y(n_5157)
);

INVxp33_ASAP7_75t_L g5158 ( 
.A(n_5112),
.Y(n_5158)
);

INVxp67_ASAP7_75t_L g5159 ( 
.A(n_5094),
.Y(n_5159)
);

NOR2xp33_ASAP7_75t_SL g5160 ( 
.A(n_5117),
.B(n_5060),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_5097),
.Y(n_5161)
);

XOR2x2_ASAP7_75t_L g5162 ( 
.A(n_5108),
.B(n_5063),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_5109),
.B(n_4908),
.Y(n_5163)
);

INVxp67_ASAP7_75t_SL g5164 ( 
.A(n_5083),
.Y(n_5164)
);

INVx1_ASAP7_75t_SL g5165 ( 
.A(n_5103),
.Y(n_5165)
);

OR2x2_ASAP7_75t_L g5166 ( 
.A(n_5123),
.B(n_5075),
.Y(n_5166)
);

AND2x2_ASAP7_75t_L g5167 ( 
.A(n_5127),
.B(n_4801),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_L g5168 ( 
.A(n_5125),
.B(n_4908),
.Y(n_5168)
);

INVx2_ASAP7_75t_L g5169 ( 
.A(n_5080),
.Y(n_5169)
);

INVx1_ASAP7_75t_SL g5170 ( 
.A(n_5083),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_5116),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_5116),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_5153),
.B(n_4965),
.Y(n_5173)
);

NOR2xp33_ASAP7_75t_L g5174 ( 
.A(n_5165),
.B(n_5117),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_5135),
.Y(n_5175)
);

OAI322xp33_ASAP7_75t_L g5176 ( 
.A1(n_5160),
.A2(n_5089),
.A3(n_5079),
.B1(n_5098),
.B2(n_4969),
.C1(n_4970),
.C2(n_4962),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_5135),
.Y(n_5177)
);

OAI21xp5_ASAP7_75t_SL g5178 ( 
.A1(n_5165),
.A2(n_4965),
.B(n_5107),
.Y(n_5178)
);

OAI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_5159),
.A2(n_4852),
.B1(n_5081),
.B2(n_5092),
.Y(n_5179)
);

INVx2_ASAP7_75t_L g5180 ( 
.A(n_5153),
.Y(n_5180)
);

CKINVDCx16_ASAP7_75t_R g5181 ( 
.A(n_5160),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_5133),
.Y(n_5182)
);

OAI21xp33_ASAP7_75t_L g5183 ( 
.A1(n_5158),
.A2(n_5086),
.B(n_5071),
.Y(n_5183)
);

AOI31xp33_ASAP7_75t_L g5184 ( 
.A1(n_5134),
.A2(n_5096),
.A3(n_5106),
.B(n_5124),
.Y(n_5184)
);

AOI22xp33_ASAP7_75t_L g5185 ( 
.A1(n_5132),
.A2(n_5162),
.B1(n_5169),
.B2(n_5147),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_5148),
.B(n_5042),
.Y(n_5186)
);

INVxp67_ASAP7_75t_L g5187 ( 
.A(n_5136),
.Y(n_5187)
);

AOI22xp5_ASAP7_75t_L g5188 ( 
.A1(n_5154),
.A2(n_4841),
.B1(n_4806),
.B2(n_4807),
.Y(n_5188)
);

OAI22xp5_ASAP7_75t_L g5189 ( 
.A1(n_5149),
.A2(n_4797),
.B1(n_5119),
.B2(n_4562),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_5144),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_5136),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5168),
.Y(n_5192)
);

INVxp67_ASAP7_75t_L g5193 ( 
.A(n_5141),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_L g5194 ( 
.A(n_5148),
.B(n_5048),
.Y(n_5194)
);

OAI32xp33_ASAP7_75t_L g5195 ( 
.A1(n_5170),
.A2(n_5077),
.A3(n_4895),
.B1(n_4883),
.B2(n_4900),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_5168),
.Y(n_5196)
);

OAI21xp5_ASAP7_75t_L g5197 ( 
.A1(n_5152),
.A2(n_5066),
.B(n_5064),
.Y(n_5197)
);

AOI21xp5_ASAP7_75t_L g5198 ( 
.A1(n_5157),
.A2(n_5082),
.B(n_5099),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_5130),
.B(n_5051),
.Y(n_5199)
);

BUFx2_ASAP7_75t_SL g5200 ( 
.A(n_5129),
.Y(n_5200)
);

AOI21xp33_ASAP7_75t_L g5201 ( 
.A1(n_5170),
.A2(n_4841),
.B(n_4996),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5131),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5163),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5163),
.Y(n_5204)
);

AOI22xp5_ASAP7_75t_L g5205 ( 
.A1(n_5150),
.A2(n_4808),
.B1(n_4848),
.B2(n_4798),
.Y(n_5205)
);

AOI31xp33_ASAP7_75t_L g5206 ( 
.A1(n_5175),
.A2(n_5005),
.A3(n_4996),
.B(n_5166),
.Y(n_5206)
);

NOR2xp33_ASAP7_75t_L g5207 ( 
.A(n_5193),
.B(n_5157),
.Y(n_5207)
);

NOR2xp33_ASAP7_75t_L g5208 ( 
.A(n_5178),
.B(n_5139),
.Y(n_5208)
);

INVxp67_ASAP7_75t_SL g5209 ( 
.A(n_5173),
.Y(n_5209)
);

A2O1A1Ixp33_ASAP7_75t_L g5210 ( 
.A1(n_5174),
.A2(n_4911),
.B(n_4915),
.C(n_4908),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_5199),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5186),
.Y(n_5212)
);

AOI32xp33_ASAP7_75t_L g5213 ( 
.A1(n_5177),
.A2(n_5151),
.A3(n_5167),
.B1(n_4911),
.B2(n_4915),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_5180),
.B(n_5072),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_5194),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_5182),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_5205),
.Y(n_5217)
);

NAND2xp5_ASAP7_75t_L g5218 ( 
.A(n_5181),
.B(n_4954),
.Y(n_5218)
);

O2A1O1Ixp33_ASAP7_75t_L g5219 ( 
.A1(n_5195),
.A2(n_5145),
.B(n_5142),
.C(n_5007),
.Y(n_5219)
);

OAI211xp5_ASAP7_75t_L g5220 ( 
.A1(n_5178),
.A2(n_5142),
.B(n_5145),
.C(n_5164),
.Y(n_5220)
);

INVxp67_ASAP7_75t_SL g5221 ( 
.A(n_5203),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_5200),
.Y(n_5222)
);

OR2x2_ASAP7_75t_L g5223 ( 
.A(n_5190),
.B(n_5143),
.Y(n_5223)
);

OAI21xp33_ASAP7_75t_L g5224 ( 
.A1(n_5185),
.A2(n_4848),
.B(n_4846),
.Y(n_5224)
);

AOI22xp33_ASAP7_75t_L g5225 ( 
.A1(n_5202),
.A2(n_4847),
.B1(n_4849),
.B2(n_4833),
.Y(n_5225)
);

INVxp67_ASAP7_75t_L g5226 ( 
.A(n_5184),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_5188),
.B(n_4972),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5204),
.Y(n_5228)
);

AOI22xp33_ASAP7_75t_SL g5229 ( 
.A1(n_5179),
.A2(n_4915),
.B1(n_4911),
.B2(n_4895),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5176),
.Y(n_5230)
);

AOI33xp33_ASAP7_75t_L g5231 ( 
.A1(n_5191),
.A2(n_5146),
.A3(n_5140),
.B1(n_5161),
.B2(n_5156),
.B3(n_5155),
.Y(n_5231)
);

OAI22xp33_ASAP7_75t_L g5232 ( 
.A1(n_5187),
.A2(n_4827),
.B1(n_4895),
.B2(n_4883),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_5198),
.B(n_4896),
.Y(n_5233)
);

AOI322xp5_ASAP7_75t_L g5234 ( 
.A1(n_5183),
.A2(n_5172),
.A3(n_5171),
.B1(n_5138),
.B2(n_5137),
.C1(n_5019),
.C2(n_5013),
.Y(n_5234)
);

OAI21xp5_ASAP7_75t_L g5235 ( 
.A1(n_5197),
.A2(n_5008),
.B(n_5007),
.Y(n_5235)
);

INVx2_ASAP7_75t_SL g5236 ( 
.A(n_5192),
.Y(n_5236)
);

NAND2xp5_ASAP7_75t_L g5237 ( 
.A(n_5201),
.B(n_4896),
.Y(n_5237)
);

OAI21xp33_ASAP7_75t_L g5238 ( 
.A1(n_5189),
.A2(n_4917),
.B(n_4897),
.Y(n_5238)
);

AND2x2_ASAP7_75t_L g5239 ( 
.A(n_5196),
.B(n_5008),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_5176),
.Y(n_5240)
);

INVx2_ASAP7_75t_L g5241 ( 
.A(n_5214),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_5214),
.Y(n_5242)
);

NOR3xp33_ASAP7_75t_L g5243 ( 
.A(n_5226),
.B(n_5012),
.C(n_5011),
.Y(n_5243)
);

AOI21xp5_ASAP7_75t_L g5244 ( 
.A1(n_5208),
.A2(n_5012),
.B(n_5011),
.Y(n_5244)
);

NOR2xp33_ASAP7_75t_L g5245 ( 
.A(n_5224),
.B(n_5013),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_5233),
.Y(n_5246)
);

INVx2_ASAP7_75t_SL g5247 ( 
.A(n_5223),
.Y(n_5247)
);

OAI21xp5_ASAP7_75t_L g5248 ( 
.A1(n_5207),
.A2(n_5210),
.B(n_5206),
.Y(n_5248)
);

O2A1O1Ixp5_ASAP7_75t_L g5249 ( 
.A1(n_5232),
.A2(n_5019),
.B(n_4900),
.C(n_4883),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_SL g5250 ( 
.A(n_5213),
.B(n_4900),
.Y(n_5250)
);

OAI22xp33_ASAP7_75t_L g5251 ( 
.A1(n_5240),
.A2(n_4825),
.B1(n_4838),
.B2(n_4828),
.Y(n_5251)
);

AOI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_5219),
.A2(n_4869),
.B(n_4867),
.Y(n_5252)
);

OAI21xp5_ASAP7_75t_SL g5253 ( 
.A1(n_5220),
.A2(n_4897),
.B(n_4917),
.Y(n_5253)
);

INVx1_ASAP7_75t_SL g5254 ( 
.A(n_5218),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5239),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5225),
.B(n_4671),
.Y(n_5256)
);

OR2x2_ASAP7_75t_L g5257 ( 
.A(n_5211),
.B(n_4815),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5231),
.Y(n_5258)
);

AOI22xp5_ASAP7_75t_L g5259 ( 
.A1(n_5222),
.A2(n_4825),
.B1(n_4838),
.B2(n_4828),
.Y(n_5259)
);

AOI21xp33_ASAP7_75t_L g5260 ( 
.A1(n_5221),
.A2(n_4869),
.B(n_4867),
.Y(n_5260)
);

OR2x2_ASAP7_75t_L g5261 ( 
.A(n_5230),
.B(n_4795),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5237),
.Y(n_5262)
);

INVxp67_ASAP7_75t_L g5263 ( 
.A(n_5227),
.Y(n_5263)
);

OAI21xp5_ASAP7_75t_L g5264 ( 
.A1(n_5217),
.A2(n_4741),
.B(n_4739),
.Y(n_5264)
);

OAI21xp5_ASAP7_75t_L g5265 ( 
.A1(n_5209),
.A2(n_4741),
.B(n_4739),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_5235),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5229),
.Y(n_5267)
);

AOI22xp5_ASAP7_75t_L g5268 ( 
.A1(n_5236),
.A2(n_4845),
.B1(n_4603),
.B2(n_4754),
.Y(n_5268)
);

OAI21xp33_ASAP7_75t_L g5269 ( 
.A1(n_5238),
.A2(n_4845),
.B(n_4687),
.Y(n_5269)
);

AOI322xp5_ASAP7_75t_L g5270 ( 
.A1(n_5216),
.A2(n_4639),
.A3(n_4772),
.B1(n_4726),
.B2(n_4636),
.C1(n_4669),
.C2(n_4647),
.Y(n_5270)
);

AOI322xp5_ASAP7_75t_L g5271 ( 
.A1(n_5212),
.A2(n_4647),
.A3(n_4683),
.B1(n_4719),
.B2(n_4673),
.C1(n_4733),
.C2(n_4728),
.Y(n_5271)
);

OAI211xp5_ASAP7_75t_L g5272 ( 
.A1(n_5234),
.A2(n_4770),
.B(n_4781),
.C(n_4782),
.Y(n_5272)
);

AOI221xp5_ASAP7_75t_SL g5273 ( 
.A1(n_5228),
.A2(n_4747),
.B1(n_4756),
.B2(n_4695),
.C(n_4722),
.Y(n_5273)
);

AOI22xp33_ASAP7_75t_L g5274 ( 
.A1(n_5215),
.A2(n_4548),
.B1(n_4542),
.B2(n_4535),
.Y(n_5274)
);

AOI221xp5_ASAP7_75t_SL g5275 ( 
.A1(n_5251),
.A2(n_4680),
.B1(n_4689),
.B2(n_4691),
.C(n_4695),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5268),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_5264),
.B(n_4651),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_SL g5278 ( 
.A(n_5265),
.B(n_4737),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_L g5279 ( 
.A(n_5271),
.B(n_4656),
.Y(n_5279)
);

AOI221xp5_ASAP7_75t_L g5280 ( 
.A1(n_5260),
.A2(n_4737),
.B1(n_4754),
.B2(n_4764),
.C(n_4730),
.Y(n_5280)
);

XNOR2x1_ASAP7_75t_SL g5281 ( 
.A(n_5247),
.B(n_4528),
.Y(n_5281)
);

OAI221xp5_ASAP7_75t_L g5282 ( 
.A1(n_5269),
.A2(n_4688),
.B1(n_4709),
.B2(n_4717),
.C(n_4760),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_5259),
.Y(n_5283)
);

AOI21xp5_ASAP7_75t_L g5284 ( 
.A1(n_5244),
.A2(n_5250),
.B(n_5252),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5249),
.Y(n_5285)
);

OAI32xp33_ASAP7_75t_L g5286 ( 
.A1(n_5261),
.A2(n_4576),
.A3(n_4542),
.B1(n_4535),
.B2(n_4548),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_5270),
.B(n_4656),
.Y(n_5287)
);

AOI21xp33_ASAP7_75t_L g5288 ( 
.A1(n_5242),
.A2(n_4737),
.B(n_4694),
.Y(n_5288)
);

AOI221xp5_ASAP7_75t_L g5289 ( 
.A1(n_5243),
.A2(n_4693),
.B1(n_4723),
.B2(n_4700),
.C(n_4755),
.Y(n_5289)
);

AO21x1_ASAP7_75t_L g5290 ( 
.A1(n_5253),
.A2(n_5245),
.B(n_5267),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_5241),
.B(n_4686),
.Y(n_5291)
);

AND2x4_ASAP7_75t_L g5292 ( 
.A(n_5255),
.B(n_4651),
.Y(n_5292)
);

AND2x2_ASAP7_75t_L g5293 ( 
.A(n_5254),
.B(n_4629),
.Y(n_5293)
);

OAI21xp5_ASAP7_75t_L g5294 ( 
.A1(n_5256),
.A2(n_4748),
.B(n_4752),
.Y(n_5294)
);

NOR2xp67_ASAP7_75t_L g5295 ( 
.A(n_5253),
.B(n_4763),
.Y(n_5295)
);

AOI22xp33_ASAP7_75t_SL g5296 ( 
.A1(n_5272),
.A2(n_4765),
.B1(n_4722),
.B2(n_4697),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5257),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_5266),
.Y(n_5298)
);

AOI21xp5_ASAP7_75t_L g5299 ( 
.A1(n_5248),
.A2(n_4591),
.B(n_4707),
.Y(n_5299)
);

HB1xp67_ASAP7_75t_L g5300 ( 
.A(n_5258),
.Y(n_5300)
);

HB1xp67_ASAP7_75t_L g5301 ( 
.A(n_5246),
.Y(n_5301)
);

INVxp67_ASAP7_75t_SL g5302 ( 
.A(n_5263),
.Y(n_5302)
);

OAI21xp33_ASAP7_75t_L g5303 ( 
.A1(n_5274),
.A2(n_4742),
.B(n_4718),
.Y(n_5303)
);

INVxp67_ASAP7_75t_L g5304 ( 
.A(n_5262),
.Y(n_5304)
);

NAND4xp25_ASAP7_75t_L g5305 ( 
.A(n_5273),
.B(n_4716),
.C(n_4613),
.D(n_4745),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_SL g5306 ( 
.A1(n_5247),
.A2(n_4660),
.B(n_4648),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5268),
.Y(n_5307)
);

OAI221xp5_ASAP7_75t_L g5308 ( 
.A1(n_5296),
.A2(n_4576),
.B1(n_4727),
.B2(n_4697),
.C(n_4691),
.Y(n_5308)
);

NAND3xp33_ASAP7_75t_L g5309 ( 
.A(n_5284),
.B(n_4589),
.C(n_4586),
.Y(n_5309)
);

NOR3xp33_ASAP7_75t_L g5310 ( 
.A(n_5298),
.B(n_4660),
.C(n_4624),
.Y(n_5310)
);

AOI211xp5_ASAP7_75t_L g5311 ( 
.A1(n_5288),
.A2(n_4680),
.B(n_4727),
.C(n_4689),
.Y(n_5311)
);

AOI211xp5_ASAP7_75t_L g5312 ( 
.A1(n_5290),
.A2(n_4606),
.B(n_4605),
.C(n_4602),
.Y(n_5312)
);

INVxp67_ASAP7_75t_SL g5313 ( 
.A(n_5281),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5295),
.Y(n_5314)
);

OAI22xp5_ASAP7_75t_L g5315 ( 
.A1(n_5291),
.A2(n_4605),
.B1(n_4586),
.B2(n_4601),
.Y(n_5315)
);

AND2x2_ASAP7_75t_L g5316 ( 
.A(n_5293),
.B(n_4629),
.Y(n_5316)
);

AOI21xp5_ASAP7_75t_L g5317 ( 
.A1(n_5278),
.A2(n_4540),
.B(n_4547),
.Y(n_5317)
);

NAND4xp25_ASAP7_75t_L g5318 ( 
.A(n_5287),
.B(n_4606),
.C(n_4601),
.D(n_4602),
.Y(n_5318)
);

OAI211xp5_ASAP7_75t_L g5319 ( 
.A1(n_5300),
.A2(n_4522),
.B(n_4527),
.C(n_4622),
.Y(n_5319)
);

NOR2xp33_ASAP7_75t_L g5320 ( 
.A(n_5292),
.B(n_4618),
.Y(n_5320)
);

AOI22xp5_ASAP7_75t_L g5321 ( 
.A1(n_5292),
.A2(n_4522),
.B1(n_4527),
.B2(n_4547),
.Y(n_5321)
);

AOI221xp5_ASAP7_75t_L g5322 ( 
.A1(n_5286),
.A2(n_4547),
.B1(n_4619),
.B2(n_4653),
.C(n_4658),
.Y(n_5322)
);

NOR2x1_ASAP7_75t_L g5323 ( 
.A(n_5285),
.B(n_4655),
.Y(n_5323)
);

NOR3x1_ASAP7_75t_L g5324 ( 
.A(n_5279),
.B(n_4617),
.C(n_4560),
.Y(n_5324)
);

AOI221xp5_ASAP7_75t_L g5325 ( 
.A1(n_5303),
.A2(n_4619),
.B1(n_4652),
.B2(n_4623),
.C(n_4529),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5280),
.B(n_4655),
.Y(n_5326)
);

NOR2xp33_ASAP7_75t_L g5327 ( 
.A(n_5305),
.B(n_4638),
.Y(n_5327)
);

OA21x2_ASAP7_75t_SL g5328 ( 
.A1(n_5282),
.A2(n_4648),
.B(n_4659),
.Y(n_5328)
);

AOI221x1_ASAP7_75t_L g5329 ( 
.A1(n_5276),
.A2(n_4614),
.B1(n_4529),
.B2(n_4628),
.C(n_4612),
.Y(n_5329)
);

AOI21xp5_ASAP7_75t_L g5330 ( 
.A1(n_5299),
.A2(n_4592),
.B(n_4615),
.Y(n_5330)
);

OAI211xp5_ASAP7_75t_SL g5331 ( 
.A1(n_5307),
.A2(n_4615),
.B(n_4609),
.C(n_4614),
.Y(n_5331)
);

OAI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_5304),
.A2(n_4569),
.B(n_4628),
.Y(n_5332)
);

OAI211xp5_ASAP7_75t_SL g5333 ( 
.A1(n_5283),
.A2(n_4769),
.B(n_598),
.C(n_600),
.Y(n_5333)
);

AOI21xp5_ASAP7_75t_L g5334 ( 
.A1(n_5302),
.A2(n_4592),
.B(n_4523),
.Y(n_5334)
);

NOR3xp33_ASAP7_75t_L g5335 ( 
.A(n_5297),
.B(n_4582),
.C(n_4648),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_5277),
.Y(n_5336)
);

AOI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_5301),
.A2(n_4592),
.B(n_4523),
.Y(n_5337)
);

INVxp67_ASAP7_75t_L g5338 ( 
.A(n_5323),
.Y(n_5338)
);

OAI21xp33_ASAP7_75t_L g5339 ( 
.A1(n_5318),
.A2(n_5294),
.B(n_5289),
.Y(n_5339)
);

NOR2xp67_ASAP7_75t_L g5340 ( 
.A(n_5309),
.B(n_597),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_5310),
.B(n_5306),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5316),
.B(n_5312),
.Y(n_5342)
);

AOI21xp5_ASAP7_75t_L g5343 ( 
.A1(n_5326),
.A2(n_5275),
.B(n_4523),
.Y(n_5343)
);

AND3x1_ASAP7_75t_L g5344 ( 
.A(n_5314),
.B(n_4556),
.C(n_4566),
.Y(n_5344)
);

NAND4xp25_ASAP7_75t_L g5345 ( 
.A(n_5327),
.B(n_4569),
.C(n_4566),
.D(n_4608),
.Y(n_5345)
);

OAI211xp5_ASAP7_75t_SL g5346 ( 
.A1(n_5336),
.A2(n_4769),
.B(n_602),
.C(n_603),
.Y(n_5346)
);

AOI21xp5_ASAP7_75t_L g5347 ( 
.A1(n_5313),
.A2(n_4536),
.B(n_4597),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_SL g5348 ( 
.A(n_5315),
.B(n_4608),
.Y(n_5348)
);

AOI22xp33_ASAP7_75t_L g5349 ( 
.A1(n_5335),
.A2(n_4536),
.B1(n_4649),
.B2(n_4557),
.Y(n_5349)
);

NAND4xp25_ASAP7_75t_L g5350 ( 
.A(n_5324),
.B(n_4621),
.C(n_4524),
.D(n_4551),
.Y(n_5350)
);

AOI21xp5_ASAP7_75t_L g5351 ( 
.A1(n_5317),
.A2(n_4536),
.B(n_4597),
.Y(n_5351)
);

NAND3xp33_ASAP7_75t_SL g5352 ( 
.A(n_5322),
.B(n_5319),
.C(n_5334),
.Y(n_5352)
);

OAI211xp5_ASAP7_75t_L g5353 ( 
.A1(n_5332),
.A2(n_4582),
.B(n_4607),
.C(n_4597),
.Y(n_5353)
);

AOI221xp5_ASAP7_75t_L g5354 ( 
.A1(n_5331),
.A2(n_4557),
.B1(n_4649),
.B2(n_4551),
.C(n_4524),
.Y(n_5354)
);

AOI21xp5_ASAP7_75t_L g5355 ( 
.A1(n_5320),
.A2(n_4616),
.B(n_4607),
.Y(n_5355)
);

OAI211xp5_ASAP7_75t_SL g5356 ( 
.A1(n_5330),
.A2(n_4769),
.B(n_604),
.C(n_605),
.Y(n_5356)
);

NAND2xp5_ASAP7_75t_SL g5357 ( 
.A(n_5337),
.B(n_4621),
.Y(n_5357)
);

AOI22xp33_ASAP7_75t_L g5358 ( 
.A1(n_5325),
.A2(n_4649),
.B1(n_4557),
.B2(n_4554),
.Y(n_5358)
);

AOI211xp5_ASAP7_75t_L g5359 ( 
.A1(n_5339),
.A2(n_5333),
.B(n_5308),
.C(n_5311),
.Y(n_5359)
);

NAND4xp25_ASAP7_75t_L g5360 ( 
.A(n_5340),
.B(n_5328),
.C(n_5329),
.D(n_5321),
.Y(n_5360)
);

NAND3xp33_ASAP7_75t_SL g5361 ( 
.A(n_5338),
.B(n_4552),
.C(n_4769),
.Y(n_5361)
);

AOI21xp5_ASAP7_75t_L g5362 ( 
.A1(n_5341),
.A2(n_4616),
.B(n_4554),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5344),
.Y(n_5363)
);

NOR3xp33_ASAP7_75t_L g5364 ( 
.A(n_5342),
.B(n_601),
.C(n_605),
.Y(n_5364)
);

AND2x2_ASAP7_75t_L g5365 ( 
.A(n_5348),
.B(n_4555),
.Y(n_5365)
);

NAND4xp25_ASAP7_75t_L g5366 ( 
.A(n_5343),
.B(n_4594),
.C(n_4584),
.D(n_4555),
.Y(n_5366)
);

NAND4xp25_ASAP7_75t_SL g5367 ( 
.A(n_5347),
.B(n_4584),
.C(n_4594),
.D(n_4581),
.Y(n_5367)
);

OAI211xp5_ASAP7_75t_L g5368 ( 
.A1(n_5352),
.A2(n_4607),
.B(n_4625),
.C(n_608),
.Y(n_5368)
);

AOI221xp5_ASAP7_75t_L g5369 ( 
.A1(n_5356),
.A2(n_4552),
.B1(n_4581),
.B2(n_4580),
.C(n_4620),
.Y(n_5369)
);

NAND5xp2_ASAP7_75t_L g5370 ( 
.A(n_5351),
.B(n_4552),
.C(n_607),
.D(n_608),
.E(n_609),
.Y(n_5370)
);

AOI21xp33_ASAP7_75t_L g5371 ( 
.A1(n_5357),
.A2(n_5346),
.B(n_5353),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_5345),
.Y(n_5372)
);

NAND3xp33_ASAP7_75t_L g5373 ( 
.A(n_5354),
.B(n_4616),
.C(n_4625),
.Y(n_5373)
);

NAND4xp25_ASAP7_75t_L g5374 ( 
.A(n_5350),
.B(n_606),
.C(n_607),
.D(n_609),
.Y(n_5374)
);

NAND3xp33_ASAP7_75t_SL g5375 ( 
.A(n_5358),
.B(n_606),
.C(n_610),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_5362),
.B(n_5355),
.Y(n_5376)
);

NAND4xp25_ASAP7_75t_SL g5377 ( 
.A(n_5368),
.B(n_5349),
.C(n_4580),
.D(n_612),
.Y(n_5377)
);

AND4x1_ASAP7_75t_L g5378 ( 
.A(n_5359),
.B(n_610),
.C(n_611),
.D(n_612),
.Y(n_5378)
);

NOR3xp33_ASAP7_75t_L g5379 ( 
.A(n_5372),
.B(n_611),
.C(n_613),
.Y(n_5379)
);

NAND4xp75_ASAP7_75t_L g5380 ( 
.A(n_5363),
.B(n_4625),
.C(n_615),
.D(n_616),
.Y(n_5380)
);

NAND3xp33_ASAP7_75t_L g5381 ( 
.A(n_5364),
.B(n_4616),
.C(n_615),
.Y(n_5381)
);

NAND4xp25_ASAP7_75t_L g5382 ( 
.A(n_5374),
.B(n_614),
.C(n_616),
.D(n_617),
.Y(n_5382)
);

NAND4xp25_ASAP7_75t_SL g5383 ( 
.A(n_5373),
.B(n_614),
.C(n_618),
.D(n_619),
.Y(n_5383)
);

NAND3xp33_ASAP7_75t_L g5384 ( 
.A(n_5371),
.B(n_618),
.C(n_619),
.Y(n_5384)
);

NOR3xp33_ASAP7_75t_SL g5385 ( 
.A(n_5360),
.B(n_620),
.C(n_621),
.Y(n_5385)
);

AOI21xp33_ASAP7_75t_L g5386 ( 
.A1(n_5365),
.A2(n_620),
.B(n_621),
.Y(n_5386)
);

NOR3xp33_ASAP7_75t_SL g5387 ( 
.A(n_5375),
.B(n_622),
.C(n_623),
.Y(n_5387)
);

NOR3xp33_ASAP7_75t_SL g5388 ( 
.A(n_5370),
.B(n_622),
.C(n_623),
.Y(n_5388)
);

OAI211xp5_ASAP7_75t_SL g5389 ( 
.A1(n_5369),
.A2(n_624),
.B(n_625),
.C(n_626),
.Y(n_5389)
);

NOR2x1_ASAP7_75t_L g5390 ( 
.A(n_5366),
.B(n_5361),
.Y(n_5390)
);

HB1xp67_ASAP7_75t_L g5391 ( 
.A(n_5367),
.Y(n_5391)
);

NOR3xp33_ASAP7_75t_L g5392 ( 
.A(n_5372),
.B(n_624),
.C(n_626),
.Y(n_5392)
);

AND4x1_ASAP7_75t_L g5393 ( 
.A(n_5359),
.B(n_627),
.C(n_628),
.D(n_629),
.Y(n_5393)
);

NAND3xp33_ASAP7_75t_SL g5394 ( 
.A(n_5359),
.B(n_629),
.C(n_630),
.Y(n_5394)
);

NOR2x1_ASAP7_75t_L g5395 ( 
.A(n_5384),
.B(n_4620),
.Y(n_5395)
);

OA22x2_ASAP7_75t_L g5396 ( 
.A1(n_5391),
.A2(n_630),
.B1(n_631),
.B2(n_632),
.Y(n_5396)
);

AOI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_5380),
.A2(n_4620),
.B1(n_632),
.B2(n_634),
.Y(n_5397)
);

AND2x4_ASAP7_75t_L g5398 ( 
.A(n_5388),
.B(n_631),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5378),
.Y(n_5399)
);

AOI22xp5_ASAP7_75t_L g5400 ( 
.A1(n_5379),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5393),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5385),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_5394),
.Y(n_5403)
);

NOR2xp33_ASAP7_75t_L g5404 ( 
.A(n_5382),
.B(n_635),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5392),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_L g5406 ( 
.A(n_5386),
.B(n_636),
.Y(n_5406)
);

AOI22xp5_ASAP7_75t_L g5407 ( 
.A1(n_5381),
.A2(n_638),
.B1(n_639),
.B2(n_640),
.Y(n_5407)
);

AOI22xp5_ASAP7_75t_L g5408 ( 
.A1(n_5383),
.A2(n_638),
.B1(n_639),
.B2(n_641),
.Y(n_5408)
);

NOR2x1_ASAP7_75t_L g5409 ( 
.A(n_5390),
.B(n_641),
.Y(n_5409)
);

AOI22xp5_ASAP7_75t_L g5410 ( 
.A1(n_5377),
.A2(n_642),
.B1(n_643),
.B2(n_645),
.Y(n_5410)
);

AND3x4_ASAP7_75t_L g5411 ( 
.A(n_5387),
.B(n_642),
.C(n_645),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5389),
.Y(n_5412)
);

AO22x2_ASAP7_75t_L g5413 ( 
.A1(n_5403),
.A2(n_5376),
.B1(n_647),
.B2(n_649),
.Y(n_5413)
);

NAND4xp75_ASAP7_75t_L g5414 ( 
.A(n_5409),
.B(n_646),
.C(n_647),
.D(n_649),
.Y(n_5414)
);

NAND3xp33_ASAP7_75t_L g5415 ( 
.A(n_5410),
.B(n_646),
.C(n_650),
.Y(n_5415)
);

NOR3xp33_ASAP7_75t_L g5416 ( 
.A(n_5405),
.B(n_650),
.C(n_651),
.Y(n_5416)
);

OAI211xp5_ASAP7_75t_SL g5417 ( 
.A1(n_5402),
.A2(n_652),
.B(n_653),
.C(n_654),
.Y(n_5417)
);

NOR4xp75_ASAP7_75t_L g5418 ( 
.A(n_5406),
.B(n_5411),
.C(n_5404),
.D(n_5396),
.Y(n_5418)
);

NOR3xp33_ASAP7_75t_L g5419 ( 
.A(n_5399),
.B(n_652),
.C(n_654),
.Y(n_5419)
);

OAI211xp5_ASAP7_75t_L g5420 ( 
.A1(n_5407),
.A2(n_655),
.B(n_656),
.C(n_657),
.Y(n_5420)
);

AOI221xp5_ASAP7_75t_L g5421 ( 
.A1(n_5412),
.A2(n_5398),
.B1(n_5401),
.B2(n_5397),
.C(n_5408),
.Y(n_5421)
);

NAND3xp33_ASAP7_75t_SL g5422 ( 
.A(n_5400),
.B(n_655),
.C(n_657),
.Y(n_5422)
);

NAND3xp33_ASAP7_75t_SL g5423 ( 
.A(n_5395),
.B(n_658),
.C(n_659),
.Y(n_5423)
);

NOR3xp33_ASAP7_75t_L g5424 ( 
.A(n_5409),
.B(n_658),
.C(n_659),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5413),
.Y(n_5425)
);

NOR2xp33_ASAP7_75t_L g5426 ( 
.A(n_5415),
.B(n_660),
.Y(n_5426)
);

HB1xp67_ASAP7_75t_L g5427 ( 
.A(n_5414),
.Y(n_5427)
);

NOR2xp33_ASAP7_75t_R g5428 ( 
.A(n_5423),
.B(n_661),
.Y(n_5428)
);

NOR3xp33_ASAP7_75t_L g5429 ( 
.A(n_5421),
.B(n_661),
.C(n_662),
.Y(n_5429)
);

OAI21xp33_ASAP7_75t_L g5430 ( 
.A1(n_5420),
.A2(n_662),
.B(n_663),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5413),
.Y(n_5431)
);

NOR2xp33_ASAP7_75t_SL g5432 ( 
.A(n_5427),
.B(n_5424),
.Y(n_5432)
);

INVx3_ASAP7_75t_L g5433 ( 
.A(n_5425),
.Y(n_5433)
);

NAND4xp75_ASAP7_75t_L g5434 ( 
.A(n_5431),
.B(n_5426),
.C(n_5418),
.D(n_5428),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5433),
.Y(n_5435)
);

AOI221xp5_ASAP7_75t_SL g5436 ( 
.A1(n_5432),
.A2(n_5430),
.B1(n_5422),
.B2(n_5429),
.C(n_5417),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5435),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5437),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5438),
.Y(n_5439)
);

AOI21xp5_ASAP7_75t_L g5440 ( 
.A1(n_5439),
.A2(n_5434),
.B(n_5436),
.Y(n_5440)
);

XNOR2xp5_ASAP7_75t_L g5441 ( 
.A(n_5440),
.B(n_5416),
.Y(n_5441)
);

AOI22xp33_ASAP7_75t_L g5442 ( 
.A1(n_5441),
.A2(n_5419),
.B1(n_665),
.B2(n_666),
.Y(n_5442)
);

OR2x2_ASAP7_75t_L g5443 ( 
.A(n_5442),
.B(n_664),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5443),
.Y(n_5444)
);

AOI21xp5_ASAP7_75t_L g5445 ( 
.A1(n_5444),
.A2(n_665),
.B(n_666),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_5445),
.Y(n_5446)
);

INVxp67_ASAP7_75t_L g5447 ( 
.A(n_5445),
.Y(n_5447)
);

AND2x2_ASAP7_75t_L g5448 ( 
.A(n_5446),
.B(n_669),
.Y(n_5448)
);

OA22x2_ASAP7_75t_L g5449 ( 
.A1(n_5447),
.A2(n_670),
.B1(n_671),
.B2(n_672),
.Y(n_5449)
);

AOI32xp33_ASAP7_75t_L g5450 ( 
.A1(n_5448),
.A2(n_670),
.A3(n_671),
.B1(n_673),
.B2(n_674),
.Y(n_5450)
);

AOI221xp5_ASAP7_75t_L g5451 ( 
.A1(n_5449),
.A2(n_675),
.B1(n_676),
.B2(n_677),
.C(n_678),
.Y(n_5451)
);

AOI221xp5_ASAP7_75t_L g5452 ( 
.A1(n_5451),
.A2(n_5450),
.B1(n_677),
.B2(n_679),
.C(n_680),
.Y(n_5452)
);

AOI211xp5_ASAP7_75t_L g5453 ( 
.A1(n_5452),
.A2(n_675),
.B(n_679),
.C(n_680),
.Y(n_5453)
);


endmodule