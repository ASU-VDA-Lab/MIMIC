module real_jpeg_29489_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_11),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_17),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_3),
.B(n_13),
.CON(n_18),
.SN(n_18)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_9),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_5),
.B(n_8),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_8),
.Y(n_35)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_14),
.B(n_20),
.C(n_27),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_9),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_12),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_32),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);


endmodule