module fake_aes_5071_n_10 (n_1, n_2, n_0, n_10);
input n_1;
input n_2;
input n_0;
output n_10;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
BUFx3_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
AND2x4_ASAP7_75t_L g4 ( .A(n_1), .B(n_0), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
OAI33xp33_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .A3(n_1), .B1(n_3), .B2(n_4), .B3(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_7), .B(n_4), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
INVxp67_ASAP7_75t_SL g10 ( .A(n_9), .Y(n_10) );
endmodule