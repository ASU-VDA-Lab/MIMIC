module fake_jpeg_3705_n_591 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_591);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_591;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_10),
.B(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx8_ASAP7_75t_SL g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_57),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_64),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_83),
.Y(n_141)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_72),
.Y(n_206)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g148 ( 
.A(n_76),
.Y(n_148)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_1),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_22),
.Y(n_86)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_88),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_26),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_1),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_103),
.Y(n_211)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_29),
.Y(n_126)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_29),
.Y(n_127)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_49),
.B1(n_29),
.B2(n_50),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_132),
.A2(n_136),
.B1(n_142),
.B2(n_150),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_42),
.B1(n_52),
.B2(n_36),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_83),
.A2(n_56),
.B1(n_50),
.B2(n_52),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_143),
.B(n_145),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_90),
.B(n_56),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_65),
.B(n_26),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_149),
.B(n_170),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_77),
.A2(n_49),
.B1(n_29),
.B2(n_44),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_49),
.B1(n_46),
.B2(n_44),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_161),
.A2(n_163),
.B1(n_171),
.B2(n_199),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_86),
.A2(n_46),
.B(n_43),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_162),
.B(n_14),
.C(n_15),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_61),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_37),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_115),
.A2(n_29),
.B1(n_36),
.B2(n_20),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_67),
.B(n_20),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_176),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_2),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_174),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_3),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_87),
.B(n_3),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_193),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_70),
.B(n_4),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_72),
.B(n_5),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_213),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_114),
.A2(n_22),
.B1(n_7),
.B2(n_8),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_79),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_245)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_82),
.B(n_5),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_5),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_9),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_88),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_171),
.B1(n_150),
.B2(n_199),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_161),
.A2(n_108),
.B1(n_103),
.B2(n_101),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_221),
.A2(n_245),
.B1(n_248),
.B2(n_284),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_222),
.B(n_241),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_100),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_223),
.B(n_270),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_146),
.A2(n_141),
.B(n_145),
.C(n_149),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_224),
.B(n_269),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_226),
.Y(n_327)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_229),
.Y(n_310)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

INVx11_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_231),
.Y(n_334)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_146),
.A2(n_98),
.B1(n_92),
.B2(n_89),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_240),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_176),
.A2(n_84),
.B1(n_12),
.B2(n_13),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_132),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_244),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_131),
.B(n_13),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_247),
.B(n_250),
.Y(n_332)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_249),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_159),
.B(n_14),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_253),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_157),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_133),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_260),
.Y(n_344)
);

NAND2x1_ASAP7_75t_L g346 ( 
.A(n_261),
.B(n_231),
.Y(n_346)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_262),
.Y(n_331)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_153),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_187),
.B(n_15),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_265),
.B(n_288),
.Y(n_355)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_181),
.Y(n_266)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_129),
.B(n_17),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_135),
.B(n_17),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_138),
.B(n_15),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_139),
.A2(n_15),
.B1(n_16),
.B2(n_166),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_274),
.A2(n_285),
.B1(n_291),
.B2(n_294),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_154),
.A2(n_16),
.B1(n_167),
.B2(n_202),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_275),
.A2(n_279),
.B1(n_292),
.B2(n_293),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_218),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_140),
.B(n_156),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_174),
.A2(n_169),
.B1(n_160),
.B2(n_164),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_173),
.B(n_130),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_283),
.Y(n_319)
);

BUFx6f_ASAP7_75t_SL g281 ( 
.A(n_137),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_281),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_155),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_205),
.A2(n_194),
.B1(n_217),
.B2(n_189),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_165),
.A2(n_200),
.B1(n_210),
.B2(n_158),
.Y(n_285)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_190),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_287),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_203),
.B(n_207),
.Y(n_287)
);

AO22x1_ASAP7_75t_SL g288 ( 
.A1(n_179),
.A2(n_206),
.B1(n_191),
.B2(n_220),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_178),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_184),
.B(n_208),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_209),
.A2(n_191),
.B1(n_179),
.B2(n_206),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_190),
.A2(n_205),
.B1(n_151),
.B2(n_134),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_189),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_194),
.A2(n_163),
.B1(n_136),
.B2(n_172),
.Y(n_294)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_217),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_295),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_134),
.B(n_146),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_272),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_134),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_128),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_148),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_243),
.A2(n_239),
.B1(n_268),
.B2(n_242),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_312),
.A2(n_323),
.B1(n_225),
.B2(n_276),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_237),
.A2(n_221),
.B1(n_234),
.B2(n_224),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_313),
.A2(n_316),
.B1(n_320),
.B2(n_342),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_245),
.A2(n_250),
.B1(n_247),
.B2(n_235),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_238),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_261),
.B1(n_296),
.B2(n_227),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_259),
.A2(n_241),
.B1(n_265),
.B2(n_285),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_288),
.A2(n_230),
.B(n_236),
.C(n_257),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_337),
.A2(n_344),
.B(n_327),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_284),
.A2(n_262),
.B1(n_263),
.B2(n_228),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_347),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_260),
.A2(n_289),
.B1(n_244),
.B2(n_286),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_229),
.A2(n_240),
.B1(n_253),
.B2(n_232),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_350),
.A2(n_256),
.B1(n_293),
.B2(n_295),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_249),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_368),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_358),
.B(n_364),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_255),
.B(n_267),
.C(n_226),
.Y(n_359)
);

OAI21xp33_ASAP7_75t_L g404 ( 
.A1(n_359),
.A2(n_389),
.B(n_329),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_264),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_360),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_340),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_365),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_318),
.B(n_258),
.C(n_246),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_366),
.C(n_372),
.Y(n_402)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_340),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_266),
.C(n_282),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_313),
.A2(n_281),
.B1(n_298),
.B2(n_307),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_367),
.A2(n_369),
.B1(n_373),
.B2(n_374),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_316),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_307),
.A2(n_325),
.B1(n_355),
.B2(n_312),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_306),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_304),
.C(n_309),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_325),
.A2(n_355),
.B1(n_323),
.B2(n_349),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_339),
.A2(n_315),
.B1(n_342),
.B2(n_303),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_319),
.B(n_309),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_306),
.Y(n_377)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_339),
.A2(n_315),
.B1(n_326),
.B2(n_337),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_383),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_314),
.B(n_324),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_379),
.B(n_382),
.Y(n_428)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_380),
.Y(n_426)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_338),
.B(n_314),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_339),
.A2(n_328),
.B1(n_305),
.B2(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_302),
.B(n_330),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_386),
.B(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_388),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_300),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_334),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_394),
.Y(n_432)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_392),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_302),
.B(n_330),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_393),
.B(n_395),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVxp67_ASAP7_75t_R g396 ( 
.A(n_327),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_396),
.A2(n_311),
.B(n_341),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_397),
.A2(n_317),
.B1(n_345),
.B2(n_341),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_305),
.A2(n_343),
.B1(n_336),
.B2(n_335),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_398),
.A2(n_311),
.B1(n_351),
.B2(n_352),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_329),
.C(n_308),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_413),
.C(n_414),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_L g438 ( 
.A1(n_404),
.A2(n_420),
.B(n_359),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_397),
.A2(n_353),
.B(n_321),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_358),
.B(n_308),
.C(n_310),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_362),
.B(n_368),
.C(n_366),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_375),
.A2(n_353),
.B(n_321),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_415),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_369),
.A2(n_335),
.B1(n_322),
.B2(n_310),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_418),
.A2(n_433),
.B1(n_363),
.B2(n_389),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_389),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_390),
.B1(n_394),
.B2(n_396),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_352),
.C(n_351),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_431),
.C(n_420),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_322),
.C(n_357),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_367),
.A2(n_373),
.B1(n_364),
.B2(n_356),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_356),
.B(n_384),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_434),
.B(n_425),
.Y(n_460)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_438),
.A2(n_430),
.B(n_423),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_439),
.A2(n_442),
.B1(n_446),
.B2(n_452),
.Y(n_490)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_440),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_408),
.A2(n_383),
.B1(n_378),
.B2(n_374),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_402),
.B(n_377),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_444),
.B(n_451),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_409),
.A2(n_361),
.B1(n_365),
.B2(n_386),
.Y(n_445)
);

AO21x1_ASAP7_75t_L g478 ( 
.A1(n_445),
.A2(n_417),
.B(n_424),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_393),
.B1(n_398),
.B2(n_370),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_381),
.Y(n_447)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_391),
.Y(n_449)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_434),
.A2(n_396),
.B1(n_387),
.B2(n_395),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_450),
.A2(n_461),
.B1(n_424),
.B2(n_425),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_402),
.B(n_371),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_400),
.A2(n_392),
.B1(n_385),
.B2(n_380),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_421),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_455),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_429),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_454),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_421),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_414),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_464),
.C(n_467),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_413),
.C(n_410),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_457),
.B(n_407),
.Y(n_486)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_433),
.A2(n_409),
.B1(n_400),
.B2(n_418),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_459),
.A2(n_422),
.B1(n_407),
.B2(n_426),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_430),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_410),
.A2(n_419),
.B1(n_411),
.B2(n_415),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_412),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_463),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_416),
.B(n_427),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_413),
.B(n_431),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_441),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_416),
.B(n_432),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_453),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_432),
.C(n_406),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_467),
.Y(n_468)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_447),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_480),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_488),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_475),
.A2(n_479),
.B1(n_485),
.B2(n_492),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_478),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_406),
.B1(n_427),
.B2(n_426),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_449),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_439),
.B1(n_437),
.B2(n_450),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_494),
.C(n_464),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_460),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_458),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_442),
.A2(n_459),
.B1(n_446),
.B2(n_443),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_456),
.B(n_451),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_496),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_441),
.B(n_444),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_498),
.A2(n_499),
.B1(n_504),
.B2(n_509),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_492),
.A2(n_445),
.B1(n_443),
.B2(n_455),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_501),
.B(n_508),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_493),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_502),
.B(n_505),
.Y(n_528)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_503),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_448),
.B1(n_465),
.B2(n_436),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_457),
.C(n_448),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_494),
.C(n_496),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_508),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_482),
.A2(n_469),
.B1(n_475),
.B2(n_491),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_486),
.C(n_476),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_515),
.Y(n_521)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_477),
.Y(n_513)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_513),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_471),
.C(n_481),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_473),
.Y(n_516)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_516),
.Y(n_535)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_474),
.Y(n_519)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_519),
.Y(n_525)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_491),
.Y(n_520)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_520),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_511),
.B(n_472),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_529),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_500),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_472),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_478),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_531),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_482),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_507),
.Y(n_532)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_532),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_514),
.A2(n_469),
.B(n_479),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_534),
.A2(n_510),
.B(n_520),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_523),
.A2(n_509),
.B1(n_514),
.B2(n_498),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_539),
.A2(n_550),
.B1(n_537),
.B2(n_536),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_506),
.Y(n_540)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_540),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_522),
.B(n_484),
.Y(n_542)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_506),
.C(n_501),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_543),
.Y(n_554)
);

INVx11_ASAP7_75t_L g544 ( 
.A(n_525),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_547),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_505),
.C(n_504),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_524),
.C(n_497),
.Y(n_555)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_532),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_535),
.Y(n_563)
);

XNOR2x1_ASAP7_75t_SL g549 ( 
.A(n_530),
.B(n_515),
.Y(n_549)
);

FAx1_ASAP7_75t_SL g558 ( 
.A(n_549),
.B(n_497),
.CI(n_521),
.CON(n_558),
.SN(n_558)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_523),
.A2(n_512),
.B1(n_499),
.B2(n_518),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_551),
.A2(n_553),
.B1(n_537),
.B2(n_536),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_555),
.B(n_561),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_560),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_534),
.C(n_510),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_488),
.C(n_513),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_561),
.B(n_563),
.Y(n_568)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_562),
.Y(n_571)
);

BUFx24_ASAP7_75t_SL g564 ( 
.A(n_542),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_546),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_565),
.B(n_547),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_554),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_570),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g569 ( 
.A1(n_557),
.A2(n_553),
.B(n_550),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_569),
.B(n_572),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_573),
.B(n_574),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_556),
.A2(n_541),
.B(n_546),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_571),
.B(n_560),
.C(n_555),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_576),
.B(n_577),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_571),
.A2(n_565),
.B1(n_551),
.B2(n_559),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_568),
.B(n_539),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_580),
.B(n_552),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_575),
.B(n_566),
.C(n_541),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_583),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g584 ( 
.A1(n_578),
.A2(n_558),
.B(n_549),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_584),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_586),
.A2(n_582),
.B(n_579),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_587),
.A2(n_585),
.B1(n_577),
.B2(n_579),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_588),
.A2(n_576),
.B(n_558),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_552),
.C(n_533),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_527),
.Y(n_591)
);


endmodule