module fake_jpeg_14021_n_426 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx12_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_65),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_66),
.Y(n_160)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_83),
.Y(n_128)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_29),
.A2(n_15),
.B(n_13),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_29),
.B(n_13),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_24),
.B(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_89),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_16),
.B(n_0),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_44),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_92),
.Y(n_145)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_97),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_100),
.Y(n_163)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_34),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_42),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_48),
.B1(n_44),
.B2(n_35),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_115),
.A2(n_119),
.B1(n_135),
.B2(n_150),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_118),
.B(n_130),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_60),
.A2(n_35),
.B1(n_23),
.B2(n_40),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_123),
.B(n_2),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_66),
.A2(n_27),
.B1(n_47),
.B2(n_34),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_144),
.B(n_26),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_81),
.A2(n_23),
.B1(n_40),
.B2(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_51),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_136),
.B(n_155),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_68),
.B(n_51),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_165),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_47),
.B(n_45),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_45),
.B1(n_18),
.B2(n_17),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_46),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_94),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_56),
.A2(n_62),
.B1(n_61),
.B2(n_73),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_85),
.A2(n_18),
.B1(n_17),
.B2(n_46),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_106),
.B1(n_104),
.B2(n_103),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_26),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_192),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_70),
.B1(n_64),
.B2(n_57),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_179),
.A2(n_195),
.B1(n_218),
.B2(n_171),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_113),
.A2(n_134),
.B1(n_162),
.B2(n_88),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_180),
.A2(n_221),
.B(n_184),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_181),
.B(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_156),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_188),
.Y(n_232)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_97),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_97),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_189),
.B(n_198),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_16),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_87),
.B1(n_79),
.B2(n_68),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_193),
.A2(n_216),
.B1(n_220),
.B2(n_230),
.Y(n_270)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_84),
.B1(n_111),
.B2(n_110),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_196),
.A2(n_197),
.B1(n_213),
.B2(n_145),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_135),
.A2(n_102),
.B1(n_96),
.B2(n_87),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_116),
.B(n_79),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_1),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_208),
.Y(n_246)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_117),
.B(n_151),
.C(n_138),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_205),
.C(n_215),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_112),
.B(n_154),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_3),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_149),
.B(n_5),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_150),
.A2(n_119),
.B1(n_115),
.B2(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_214),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_5),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_157),
.A2(n_164),
.B1(n_160),
.B2(n_131),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_6),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_223),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_164),
.A2(n_6),
.B1(n_8),
.B2(n_160),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_171),
.A2(n_6),
.B1(n_175),
.B2(n_176),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_161),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_224),
.Y(n_236)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_131),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_229),
.Y(n_256)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_129),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_228),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_234),
.B(n_244),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_185),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_186),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_180),
.A2(n_137),
.B1(n_142),
.B2(n_143),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_241),
.A2(n_254),
.B1(n_229),
.B2(n_222),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_181),
.B(n_131),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_145),
.B(n_172),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_248),
.A2(n_232),
.B(n_242),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_250),
.B(n_188),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_137),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_218),
.A2(n_142),
.B1(n_143),
.B2(n_169),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_190),
.A2(n_169),
.B1(n_197),
.B2(n_202),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_205),
.B1(n_182),
.B2(n_226),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_188),
.A2(n_217),
.B1(n_209),
.B2(n_215),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_265),
.B(n_243),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g265 ( 
.A1(n_177),
.A2(n_192),
.B(n_183),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_205),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_270),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_221),
.B1(n_206),
.B2(n_201),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_274),
.A2(n_294),
.B1(n_296),
.B2(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_206),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_277),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_219),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_214),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_280),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_271),
.C(n_245),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_297),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_266),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_287),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_188),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_283),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_237),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_178),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_223),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_187),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_289),
.B(n_305),
.Y(n_309)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_231),
.B1(n_258),
.B2(n_235),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_241),
.A2(n_194),
.B1(n_200),
.B2(n_210),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_291),
.A2(n_293),
.B1(n_302),
.B2(n_237),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_224),
.B(n_225),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_299),
.B(n_266),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_234),
.A2(n_211),
.B1(n_224),
.B2(n_244),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_260),
.A2(n_271),
.B1(n_263),
.B2(n_248),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_295),
.A2(n_301),
.B(n_269),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_243),
.A2(n_259),
.B1(n_253),
.B2(n_267),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_244),
.C(n_232),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_232),
.A2(n_245),
.B(n_264),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_239),
.B1(n_272),
.B2(n_238),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_272),
.B1(n_242),
.B2(n_231),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_240),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_329),
.B(n_331),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_311),
.A2(n_326),
.B(n_304),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_249),
.B1(n_266),
.B2(n_247),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_314),
.A2(n_323),
.B1(n_288),
.B2(n_303),
.Y(n_353)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_330),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_258),
.B1(n_240),
.B2(n_257),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_235),
.A3(n_257),
.B1(n_258),
.B2(n_269),
.C1(n_294),
.C2(n_274),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_273),
.A2(n_304),
.B1(n_281),
.B2(n_282),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_328),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_302),
.B1(n_290),
.B2(n_279),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_276),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_273),
.A2(n_284),
.B1(n_292),
.B2(n_275),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_309),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_335),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_299),
.B(n_283),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_344),
.B(n_283),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_289),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_288),
.Y(n_336)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_336),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_337),
.A2(n_339),
.B(n_340),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_304),
.B(n_280),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_319),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_353),
.B1(n_329),
.B2(n_320),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_327),
.A2(n_324),
.B(n_316),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_306),
.C(n_327),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_297),
.C(n_316),
.Y(n_363)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_364),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_312),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_363),
.C(n_365),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_275),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_319),
.B1(n_306),
.B2(n_322),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_360),
.A2(n_362),
.B1(n_338),
.B2(n_343),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_341),
.A2(n_330),
.B1(n_315),
.B2(n_308),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_315),
.B(n_283),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_337),
.C(n_297),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_344),
.C(n_351),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_346),
.C(n_335),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_338),
.A2(n_323),
.B1(n_314),
.B2(n_308),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_369),
.A2(n_370),
.B1(n_341),
.B2(n_346),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_338),
.A2(n_308),
.B1(n_321),
.B2(n_310),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_356),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_372),
.B(n_376),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_336),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_377),
.C(n_378),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_355),
.B(n_307),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_334),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_334),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_383),
.C(n_366),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_380),
.A2(n_382),
.B1(n_385),
.B2(n_338),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_360),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_355),
.A2(n_332),
.B1(n_340),
.B2(n_350),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_343),
.C(n_342),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_356),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_384),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_394),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_370),
.B1(n_369),
.B2(n_371),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_338),
.B1(n_354),
.B2(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_392),
.A2(n_338),
.B1(n_358),
.B2(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_393),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_381),
.A2(n_366),
.B(n_364),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_395),
.B(n_378),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_396),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_397),
.A2(n_386),
.B1(n_389),
.B2(n_394),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_399),
.A2(n_390),
.B1(n_359),
.B2(n_361),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_401),
.B(n_404),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_374),
.C(n_377),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_398),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_396),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_407),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_400),
.A2(n_388),
.B(n_395),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_409),
.A2(n_410),
.B1(n_411),
.B2(n_397),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_398),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_399),
.A2(n_367),
.B1(n_374),
.B2(n_361),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_412),
.B(n_413),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_408),
.A2(n_400),
.B(n_404),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_415),
.B(n_416),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_387),
.C(n_402),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_410),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_419),
.A2(n_359),
.B(n_368),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_373),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_420),
.A2(n_421),
.B(n_417),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_L g423 ( 
.A1(n_422),
.A2(n_409),
.B1(n_347),
.B2(n_368),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_342),
.B(n_313),
.Y(n_424)
);

AOI32xp33_ASAP7_75t_L g425 ( 
.A1(n_424),
.A2(n_313),
.A3(n_318),
.B1(n_308),
.B2(n_345),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_345),
.B(n_283),
.Y(n_426)
);


endmodule