module real_jpeg_7123_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_1),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_1),
.A2(n_124),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_1),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_1),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_25),
.B1(n_43),
.B2(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_2),
.A2(n_46),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_46),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_2),
.A2(n_46),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_2),
.A2(n_266),
.B(n_269),
.C(n_272),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_2),
.B(n_51),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_2),
.B(n_308),
.C(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_2),
.B(n_109),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_2),
.B(n_74),
.C(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_2),
.B(n_27),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_3),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_3),
.A2(n_76),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_3),
.A2(n_76),
.B1(n_179),
.B2(n_183),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_4),
.A2(n_24),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_4),
.A2(n_24),
.B1(n_71),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_4),
.A2(n_24),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_8),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_11),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_13),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_407),
.B(n_409),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_146),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_18),
.B(n_125),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_115),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_48),
.C(n_78),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_20),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_20),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_20),
.A2(n_127),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_20),
.B(n_155),
.C(n_162),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_20),
.B(n_247),
.C(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_20),
.A2(n_127),
.B1(n_247),
.B2(n_346),
.Y(n_369)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_42),
.B2(n_47),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_21),
.A2(n_26),
.B1(n_42),
.B2(n_47),
.Y(n_132)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_25),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_26),
.A2(n_42),
.B1(n_47),
.B2(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_26),
.A2(n_42),
.B(n_47),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_27)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_28),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_29),
.Y(n_143)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_30),
.Y(n_161)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_46),
.A2(n_139),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_48),
.A2(n_78),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_48),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_48),
.B(n_132),
.C(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_48),
.A2(n_131),
.B1(n_134),
.B2(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_73),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_49),
.B(n_197),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_50),
.A2(n_61),
.B1(n_191),
.B2(n_196),
.Y(n_190)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_51),
.A2(n_205),
.B(n_212),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_51),
.B(n_192),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_51),
.A2(n_62),
.B1(n_73),
.B2(n_205),
.Y(n_246)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_64),
.B1(n_67),
.B2(n_70),
.Y(n_63)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_55),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_55),
.Y(n_234)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_55),
.Y(n_279)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_57),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_58),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_58),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_62),
.B(n_197),
.Y(n_213)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_66),
.Y(n_211)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_72),
.Y(n_201)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_86),
.B1(n_109),
.B2(n_110),
.Y(n_78)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_86),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_101),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_87),
.A2(n_101),
.B1(n_138),
.B2(n_156),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_87),
.A2(n_101),
.B1(n_138),
.B2(n_156),
.Y(n_247)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_98),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_117),
.B(n_137),
.Y(n_235)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.C(n_133),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_126),
.A2(n_132),
.B1(n_259),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_126),
.Y(n_391)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_132),
.B(n_221),
.C(n_235),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_132),
.A2(n_235),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_132),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_132),
.A2(n_259),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_132),
.B(n_155),
.C(n_356),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_132),
.A2(n_259),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_133),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_134),
.Y(n_396)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_387),
.B(n_404),
.Y(n_147)
);

OAI211xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_283),
.B(n_381),
.C(n_386),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_252),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_150),
.A2(n_252),
.B(n_382),
.C(n_385),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_236),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_151),
.B(n_236),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_202),
.C(n_220),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_152),
.B(n_202),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_154),
.A2(n_155),
.B1(n_223),
.B2(n_302),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_154),
.B(n_302),
.C(n_323),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_154),
.A2(n_155),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_161),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_189),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_163),
.A2(n_189),
.B1(n_190),
.B2(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_169),
.B1(n_177),
.B2(n_186),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_165),
.A2(n_226),
.B(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_168),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_169),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_169),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_170),
.A2(n_231),
.B1(n_275),
.B2(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_170),
.A2(n_227),
.B1(n_231),
.B2(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_176),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_183),
.Y(n_309)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_189),
.A2(n_190),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_189),
.A2(n_190),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_190),
.B(n_274),
.C(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_190),
.B(n_338),
.C(n_340),
.Y(n_351)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_214),
.B2(n_219),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_214),
.Y(n_243)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_211),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_219),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_214),
.A2(n_242),
.B(n_243),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_215),
.B(n_231),
.Y(n_331)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_258),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_223),
.A2(n_302),
.B1(n_303),
.B2(n_310),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_223),
.A2(n_225),
.B1(n_302),
.B2(n_372),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_225),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_250),
.B2(n_251),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_244),
.B1(n_245),
.B2(n_249),
.Y(n_238)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_244),
.B(n_249),
.C(n_251),
.Y(n_403)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_247),
.A2(n_342),
.B1(n_343),
.B2(n_346),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_247),
.Y(n_346)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_248),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_248),
.A2(n_393),
.B1(n_397),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_253),
.B(n_255),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.C(n_263),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_263),
.B(n_379),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_264),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_265),
.A2(n_273),
.B1(n_274),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_273),
.A2(n_274),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_365),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_350),
.B(n_364),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_335),
.B(n_349),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_320),
.B(n_334),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_312),
.B(n_319),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_299),
.B(n_311),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_296),
.B(n_298),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_300),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_344),
.C(n_346),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_310),
.Y(n_318)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_322),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_333),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_332),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_332),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_348),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_348),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_340),
.B1(n_341),
.B2(n_347),
.Y(n_336)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_352),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_358),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_360),
.C(n_361),
.Y(n_374)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_375),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_374),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_374),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_373),
.C(n_377),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_383),
.B(n_384),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_378),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_399),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_405),
.B(n_406),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_392),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.C(n_398),
.Y(n_392)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_403),
.Y(n_405)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx13_ASAP7_75t_L g411 ( 
.A(n_408),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);


endmodule