module real_aes_9337_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_0), .A2(n_333), .B(n_521), .Y(n_663) );
INVx1_ASAP7_75t_L g700 ( .A(n_0), .Y(n_700) );
INVx1_ASAP7_75t_L g350 ( .A(n_1), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_1), .A2(n_77), .B1(n_434), .B2(n_440), .C(n_444), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_2), .A2(n_276), .B1(n_333), .B2(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g464 ( .A(n_2), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g1346 ( .A1(n_3), .A2(n_4), .B1(n_1322), .B2(n_1335), .Y(n_1346) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_5), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_5), .B(n_210), .Y(n_396) );
AND2x2_ASAP7_75t_L g413 ( .A(n_5), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g477 ( .A(n_5), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_6), .A2(n_18), .B1(n_742), .B2(n_1186), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_6), .A2(n_211), .B1(n_755), .B2(n_1212), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_7), .A2(n_169), .B1(n_364), .B2(n_498), .C(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g542 ( .A(n_7), .Y(n_542) );
INVxp67_ASAP7_75t_L g1010 ( .A(n_8), .Y(n_1010) );
OAI222xp33_ASAP7_75t_L g1025 ( .A1(n_8), .A2(n_42), .B1(n_267), .B2(n_754), .C1(n_1026), .C2(n_1028), .Y(n_1025) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_9), .A2(n_862), .B1(n_864), .B2(n_870), .C(n_877), .Y(n_861) );
INVx1_ASAP7_75t_L g904 ( .A(n_9), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g1328 ( .A1(n_10), .A2(n_56), .B1(n_1329), .B2(n_1332), .Y(n_1328) );
XNOR2xp5_ASAP7_75t_L g1525 ( .A(n_11), .B(n_1526), .Y(n_1525) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_12), .A2(n_55), .B1(n_417), .B2(n_853), .C(n_854), .Y(n_852) );
INVx1_ASAP7_75t_L g919 ( .A(n_12), .Y(n_919) );
INVx1_ASAP7_75t_L g843 ( .A(n_13), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_13), .A2(n_58), .B1(n_386), .B2(n_644), .Y(n_906) );
AO22x2_ASAP7_75t_L g926 ( .A1(n_14), .A2(n_927), .B1(n_984), .B2(n_985), .Y(n_926) );
CKINVDCx14_ASAP7_75t_R g984 ( .A(n_14), .Y(n_984) );
INVx1_ASAP7_75t_L g1552 ( .A(n_15), .Y(n_1552) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_16), .A2(n_36), .B1(n_362), .B2(n_363), .C(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g470 ( .A(n_16), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_17), .A2(n_265), .B1(n_577), .B2(n_787), .C(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g812 ( .A(n_17), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g1208 ( .A1(n_18), .A2(n_93), .B1(n_974), .B2(n_1209), .C(n_1210), .Y(n_1208) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_19), .A2(n_574), .B1(n_639), .B2(n_646), .C(n_653), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_19), .A2(n_190), .B1(n_674), .B2(n_686), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_20), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g1641 ( .A1(n_21), .A2(n_79), .B1(n_1642), .B2(n_1643), .Y(n_1641) );
AOI22xp33_ASAP7_75t_L g1656 ( .A1(n_21), .A2(n_79), .B1(n_515), .B2(n_1657), .Y(n_1656) );
INVx2_ASAP7_75t_L g341 ( .A(n_22), .Y(n_341) );
OR2x2_ASAP7_75t_L g359 ( .A(n_22), .B(n_346), .Y(n_359) );
AO22x1_ASAP7_75t_L g834 ( .A1(n_23), .A2(n_835), .B1(n_924), .B2(n_925), .Y(n_834) );
INVx1_ASAP7_75t_L g925 ( .A(n_23), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_24), .A2(n_246), .B1(n_592), .B2(n_594), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_24), .A2(n_246), .B1(n_440), .B2(n_444), .C(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g1013 ( .A(n_25), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_26), .A2(n_108), .B1(n_338), .B2(n_1054), .C(n_1055), .Y(n_1053) );
INVx1_ASAP7_75t_L g1081 ( .A(n_26), .Y(n_1081) );
BUFx2_ASAP7_75t_L g390 ( .A(n_27), .Y(n_390) );
OR2x2_ASAP7_75t_L g395 ( .A(n_27), .B(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g399 ( .A(n_27), .Y(n_399) );
INVx1_ASAP7_75t_L g412 ( .A(n_27), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g1189 ( .A1(n_28), .A2(n_166), .B1(n_1188), .B2(n_1190), .Y(n_1189) );
INVxp33_ASAP7_75t_SL g1216 ( .A(n_28), .Y(n_1216) );
INVx1_ASAP7_75t_L g562 ( .A(n_29), .Y(n_562) );
OAI22xp33_ASAP7_75t_L g1252 ( .A1(n_30), .A2(n_185), .B1(n_1253), .B2(n_1255), .Y(n_1252) );
INVx1_ASAP7_75t_L g1284 ( .A(n_30), .Y(n_1284) );
CKINVDCx16_ASAP7_75t_R g1323 ( .A(n_31), .Y(n_1323) );
INVx1_ASAP7_75t_L g930 ( .A(n_32), .Y(n_930) );
AOI21xp33_ASAP7_75t_L g973 ( .A1(n_32), .A2(n_386), .B(n_974), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_33), .A2(n_171), .B1(n_578), .B2(n_1064), .C(n_1066), .Y(n_1063) );
INVx1_ASAP7_75t_L g1092 ( .A(n_33), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_34), .Y(n_941) );
INVxp33_ASAP7_75t_SL g1181 ( .A(n_35), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_35), .A2(n_220), .B1(n_1057), .B2(n_1157), .C(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g455 ( .A(n_36), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_37), .Y(n_374) );
INVx1_ASAP7_75t_L g1307 ( .A(n_38), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_38), .B(n_1305), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_39), .A2(n_151), .B1(n_386), .B2(n_644), .Y(n_662) );
INVx1_ASAP7_75t_L g701 ( .A(n_39), .Y(n_701) );
INVx1_ASAP7_75t_L g999 ( .A(n_40), .Y(n_999) );
INVx1_ASAP7_75t_L g1553 ( .A(n_41), .Y(n_1553) );
INVxp67_ASAP7_75t_L g1008 ( .A(n_42), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_43), .A2(n_216), .B1(n_501), .B2(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g613 ( .A(n_43), .Y(n_613) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_44), .A2(n_111), .B1(n_736), .B2(n_737), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_44), .A2(n_70), .B1(n_652), .B2(n_765), .C(n_767), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_45), .A2(n_229), .B1(n_976), .B2(n_977), .C(n_979), .Y(n_975) );
INVx1_ASAP7_75t_L g982 ( .A(n_45), .Y(n_982) );
INVxp33_ASAP7_75t_SL g1584 ( .A(n_46), .Y(n_1584) );
AOI22xp33_ASAP7_75t_SL g1663 ( .A1(n_46), .A2(n_51), .B1(n_755), .B2(n_1034), .Y(n_1663) );
INVx1_ASAP7_75t_L g1629 ( .A(n_47), .Y(n_1629) );
AOI22xp33_ASAP7_75t_L g1649 ( .A1(n_47), .A2(n_195), .B1(n_1193), .B2(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g869 ( .A(n_48), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_48), .A2(n_159), .B1(n_499), .B2(n_644), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_49), .A2(n_172), .B1(n_856), .B2(n_860), .Y(n_855) );
OAI22xp5_ASAP7_75t_SL g888 ( .A1(n_49), .A2(n_172), .B1(n_889), .B2(n_893), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_50), .Y(n_1059) );
INVxp33_ASAP7_75t_SL g1587 ( .A(n_51), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_52), .A2(n_78), .B1(n_322), .B2(n_1250), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_52), .A2(n_78), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
INVxp33_ASAP7_75t_SL g1601 ( .A(n_53), .Y(n_1601) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_53), .A2(n_57), .B1(n_1054), .B2(n_1662), .Y(n_1661) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_54), .A2(n_190), .B1(n_376), .B2(n_382), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_54), .A2(n_273), .B1(n_677), .B2(n_682), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_55), .A2(n_117), .B1(n_921), .B2(n_922), .Y(n_920) );
INVx1_ASAP7_75t_L g1592 ( .A(n_57), .Y(n_1592) );
INVx1_ASAP7_75t_L g845 ( .A(n_58), .Y(n_845) );
AOI22xp33_ASAP7_75t_SL g1126 ( .A1(n_59), .A2(n_118), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_59), .A2(n_143), .B1(n_652), .B2(n_1153), .C(n_1155), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_60), .A2(n_71), .B1(n_362), .B2(n_577), .C(n_578), .Y(n_576) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_60), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_61), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1334 ( .A1(n_62), .A2(n_90), .B1(n_1322), .B2(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1533 ( .A(n_63), .Y(n_1533) );
INVxp33_ASAP7_75t_SL g1618 ( .A(n_64), .Y(n_1618) );
AOI22xp33_ASAP7_75t_L g1647 ( .A1(n_64), .A2(n_164), .B1(n_1642), .B2(n_1648), .Y(n_1647) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_65), .A2(n_156), .B1(n_1239), .B2(n_1241), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_65), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1535 ( .A1(n_66), .A2(n_223), .B1(n_535), .B2(n_994), .C(n_1087), .Y(n_1535) );
OAI22xp5_ASAP7_75t_L g1558 ( .A1(n_66), .A2(n_223), .B1(n_977), .B2(n_1559), .Y(n_1558) );
INVxp67_ASAP7_75t_L g1546 ( .A(n_67), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_67), .A2(n_132), .B1(n_1069), .B2(n_1568), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_68), .A2(n_198), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
INVx1_ASAP7_75t_L g1079 ( .A(n_68), .Y(n_1079) );
AOI22xp5_ASAP7_75t_SL g1342 ( .A1(n_69), .A2(n_81), .B1(n_1316), .B2(n_1322), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_70), .A2(n_136), .B1(n_730), .B2(n_733), .Y(n_729) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_71), .Y(n_621) );
INVxp33_ASAP7_75t_SL g1119 ( .A(n_72), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_72), .A2(n_212), .B1(n_499), .B2(n_644), .Y(n_1146) );
CKINVDCx16_ASAP7_75t_R g1320 ( .A(n_73), .Y(n_1320) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_74), .A2(n_88), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g763 ( .A(n_74), .Y(n_763) );
INVxp67_ASAP7_75t_SL g1117 ( .A(n_75), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_75), .A2(n_219), .B1(n_793), .B2(n_977), .C(n_1144), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_76), .A2(n_243), .B1(n_584), .B2(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g813 ( .A(n_76), .Y(n_813) );
INVx1_ASAP7_75t_L g354 ( .A(n_77), .Y(n_354) );
INVx1_ASAP7_75t_L g724 ( .A(n_80), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_80), .A2(n_105), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_82), .A2(n_162), .B1(n_787), .B2(n_788), .C(n_1040), .Y(n_1039) );
OAI221xp5_ASAP7_75t_L g1042 ( .A1(n_82), .A2(n_180), .B1(n_1043), .B2(n_1044), .C(n_1046), .Y(n_1042) );
CKINVDCx5p33_ASAP7_75t_R g1070 ( .A(n_83), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_84), .A2(n_221), .B1(n_737), .B2(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g780 ( .A(n_84), .Y(n_780) );
INVx1_ASAP7_75t_L g342 ( .A(n_85), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_85), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_86), .A2(n_259), .B1(n_501), .B2(n_504), .Y(n_500) );
INVx1_ASAP7_75t_L g553 ( .A(n_86), .Y(n_553) );
INVx1_ASAP7_75t_L g571 ( .A(n_87), .Y(n_571) );
INVx1_ASAP7_75t_L g779 ( .A(n_88), .Y(n_779) );
INVx1_ASAP7_75t_L g1245 ( .A(n_89), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_89), .A2(n_862), .B1(n_1261), .B2(n_1265), .C(n_1272), .Y(n_1260) );
INVx1_ASAP7_75t_L g647 ( .A(n_91), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_91), .A2(n_170), .B1(n_673), .B2(n_674), .Y(n_672) );
NAND2xp33_ASAP7_75t_SL g327 ( .A(n_92), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g415 ( .A(n_92), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g1187 ( .A1(n_93), .A2(n_211), .B1(n_730), .B2(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1276 ( .A(n_94), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_94), .A2(n_123), .B1(n_921), .B2(n_922), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_95), .A2(n_102), .B1(n_1193), .B2(n_1645), .Y(n_1644) );
AOI22xp33_ASAP7_75t_L g1652 ( .A1(n_95), .A2(n_102), .B1(n_1653), .B2(n_1655), .Y(n_1652) );
INVx1_ASAP7_75t_L g710 ( .A(n_96), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g989 ( .A(n_97), .B(n_990), .Y(n_989) );
INVxp67_ASAP7_75t_L g1541 ( .A(n_98), .Y(n_1541) );
AOI221xp5_ASAP7_75t_L g1564 ( .A1(n_98), .A2(n_126), .B1(n_652), .B2(n_1565), .C(n_1566), .Y(n_1564) );
INVxp33_ASAP7_75t_SL g1123 ( .A(n_99), .Y(n_1123) );
AOI21xp33_ASAP7_75t_L g1147 ( .A1(n_99), .A2(n_1148), .B(n_1149), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_100), .A2(n_635), .B1(n_705), .B2(n_706), .Y(n_634) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_100), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_101), .Y(n_803) );
INVxp67_ASAP7_75t_L g997 ( .A(n_103), .Y(n_997) );
AOI221xp5_ASAP7_75t_L g1031 ( .A1(n_103), .A2(n_178), .B1(n_362), .B2(n_363), .C(n_578), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_104), .Y(n_312) );
INVx1_ASAP7_75t_L g720 ( .A(n_105), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_106), .A2(n_1166), .B1(n_1167), .B2(n_1217), .Y(n_1165) );
INVx1_ASAP7_75t_L g1217 ( .A(n_106), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_106), .A2(n_249), .B1(n_1329), .B2(n_1386), .Y(n_1385) );
CKINVDCx5p33_ASAP7_75t_R g1196 ( .A(n_107), .Y(n_1196) );
INVx1_ASAP7_75t_L g1083 ( .A(n_108), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_109), .A2(n_231), .B1(n_577), .B2(n_652), .C(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g821 ( .A(n_109), .Y(n_821) );
INVx1_ASAP7_75t_L g1594 ( .A(n_110), .Y(n_1594) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_111), .A2(n_136), .B1(n_770), .B2(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g1180 ( .A(n_112), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_113), .A2(n_123), .B1(n_743), .B2(n_1136), .C(n_1278), .Y(n_1277) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_113), .A2(n_207), .B1(n_1288), .B2(n_1290), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_114), .A2(n_238), .B1(n_588), .B2(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g606 ( .A(n_114), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_115), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_116), .A2(n_173), .B1(n_743), .B2(n_1136), .Y(n_1135) );
INVxp33_ASAP7_75t_SL g1159 ( .A(n_116), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_117), .A2(n_134), .B1(n_849), .B2(n_850), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_118), .A2(n_122), .B1(n_1069), .B2(n_1157), .Y(n_1156) );
AOI22xp33_ASAP7_75t_SL g1192 ( .A1(n_119), .A2(n_139), .B1(n_742), .B2(n_1193), .Y(n_1192) );
INVxp33_ASAP7_75t_L g1215 ( .A(n_119), .Y(n_1215) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_120), .A2(n_222), .B1(n_333), .B2(n_521), .C(n_577), .Y(n_586) );
INVx1_ASAP7_75t_L g605 ( .A(n_120), .Y(n_605) );
INVxp33_ASAP7_75t_L g1530 ( .A(n_121), .Y(n_1530) );
AOI221xp5_ASAP7_75t_L g1560 ( .A1(n_121), .A2(n_158), .B1(n_790), .B2(n_1561), .C(n_1562), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_122), .A2(n_143), .B1(n_1131), .B2(n_1132), .Y(n_1130) );
INVx1_ASAP7_75t_L g287 ( .A(n_124), .Y(n_287) );
INVx1_ASAP7_75t_L g1162 ( .A(n_125), .Y(n_1162) );
INVxp67_ASAP7_75t_L g1543 ( .A(n_126), .Y(n_1543) );
INVx1_ASAP7_75t_L g391 ( .A(n_127), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_128), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_129), .Y(n_938) );
OA22x2_ASAP7_75t_L g781 ( .A1(n_130), .A2(n_782), .B1(n_827), .B2(n_828), .Y(n_781) );
INVx1_ASAP7_75t_L g828 ( .A(n_130), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_131), .A2(n_192), .B1(n_1131), .B2(n_1132), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_131), .Y(n_1142) );
INVx1_ASAP7_75t_L g1538 ( .A(n_132), .Y(n_1538) );
INVxp67_ASAP7_75t_SL g1172 ( .A(n_133), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_133), .A2(n_280), .B1(n_750), .B2(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g917 ( .A(n_134), .Y(n_917) );
INVx1_ASAP7_75t_L g1531 ( .A(n_135), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1341 ( .A1(n_137), .A2(n_235), .B1(n_1329), .B2(n_1332), .Y(n_1341) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_138), .A2(n_227), .B1(n_318), .B2(n_322), .Y(n_317) );
INVx1_ASAP7_75t_L g426 ( .A(n_138), .Y(n_426) );
INVxp67_ASAP7_75t_SL g1213 ( .A(n_139), .Y(n_1213) );
INVx1_ASAP7_75t_L g1121 ( .A(n_140), .Y(n_1121) );
OAI222xp33_ASAP7_75t_L g992 ( .A1(n_141), .A2(n_179), .B1(n_270), .B2(n_394), .C1(n_993), .C2(n_994), .Y(n_992) );
INVx1_ASAP7_75t_L g1019 ( .A(n_141), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_142), .A2(n_146), .B1(n_1316), .B2(n_1388), .Y(n_1387) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_144), .Y(n_523) );
INVx1_ASAP7_75t_L g1178 ( .A(n_145), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_147), .Y(n_943) );
CKINVDCx14_ASAP7_75t_R g1338 ( .A(n_148), .Y(n_1338) );
AOI22xp5_ASAP7_75t_L g1345 ( .A1(n_149), .A2(n_237), .B1(n_1329), .B2(n_1332), .Y(n_1345) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_150), .A2(n_277), .B1(n_498), .B2(n_520), .C(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g530 ( .A(n_150), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_151), .A2(n_261), .B1(n_703), .B2(n_704), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_152), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_153), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_154), .Y(n_804) );
INVx1_ASAP7_75t_L g745 ( .A(n_155), .Y(n_745) );
INVxp67_ASAP7_75t_SL g1271 ( .A(n_156), .Y(n_1271) );
INVx1_ASAP7_75t_L g510 ( .A(n_157), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_157), .A2(n_239), .B1(n_441), .B2(n_535), .C(n_537), .Y(n_534) );
INVxp33_ASAP7_75t_L g1534 ( .A(n_158), .Y(n_1534) );
INVx1_ASAP7_75t_L g867 ( .A(n_159), .Y(n_867) );
INVx1_ASAP7_75t_L g1596 ( .A(n_160), .Y(n_1596) );
INVx1_ASAP7_75t_L g1248 ( .A(n_161), .Y(n_1248) );
OAI211xp5_ASAP7_75t_SL g1273 ( .A1(n_161), .A2(n_838), .B(n_1274), .C(n_1279), .Y(n_1273) );
OAI332xp33_ASAP7_75t_L g995 ( .A1(n_162), .A2(n_447), .A3(n_630), .B1(n_951), .B2(n_996), .B3(n_1000), .C1(n_1003), .C2(n_1009), .Y(n_995) );
INVx1_ASAP7_75t_L g931 ( .A(n_163), .Y(n_931) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_163), .A2(n_205), .B1(n_644), .B2(n_972), .Y(n_971) );
INVxp67_ASAP7_75t_SL g1626 ( .A(n_164), .Y(n_1626) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_165), .Y(n_723) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_166), .Y(n_1199) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_167), .Y(n_496) );
INVx1_ASAP7_75t_L g575 ( .A(n_168), .Y(n_575) );
INVx1_ASAP7_75t_L g548 ( .A(n_169), .Y(n_548) );
INVx1_ASAP7_75t_L g642 ( .A(n_170), .Y(n_642) );
INVx1_ASAP7_75t_L g1094 ( .A(n_171), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g1151 ( .A(n_173), .Y(n_1151) );
AO221x2_ASAP7_75t_L g1336 ( .A1(n_174), .A2(n_264), .B1(n_1322), .B2(n_1335), .C(n_1337), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_175), .A2(n_224), .B1(n_394), .B2(n_703), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g966 ( .A1(n_175), .A2(n_202), .B1(n_386), .B2(n_644), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_176), .A2(n_202), .B1(n_950), .B2(n_951), .Y(n_949) );
INVx1_ASAP7_75t_L g962 ( .A(n_176), .Y(n_962) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_177), .A2(n_499), .B(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_177), .A2(n_260), .B1(n_677), .B2(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g1001 ( .A(n_178), .Y(n_1001) );
INVx1_ASAP7_75t_L g1035 ( .A(n_179), .Y(n_1035) );
INVx1_ASAP7_75t_L g1038 ( .A(n_180), .Y(n_1038) );
CKINVDCx5p33_ASAP7_75t_R g939 ( .A(n_181), .Y(n_939) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_182), .B(n_287), .Y(n_1303) );
AND3x2_ASAP7_75t_L g1319 ( .A(n_182), .B(n_287), .C(n_1306), .Y(n_1319) );
OA332x1_ASAP7_75t_L g928 ( .A1(n_183), .A2(n_447), .A3(n_929), .B1(n_934), .B2(n_937), .B3(n_940), .C1(n_945), .C2(n_946), .Y(n_928) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_183), .A2(n_521), .B(n_968), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_184), .Y(n_1225) );
INVx1_ASAP7_75t_L g1282 ( .A(n_185), .Y(n_1282) );
AOI22xp5_ASAP7_75t_SL g1354 ( .A1(n_186), .A2(n_201), .B1(n_1316), .B2(n_1322), .Y(n_1354) );
INVx2_ASAP7_75t_L g300 ( .A(n_187), .Y(n_300) );
INVx1_ASAP7_75t_L g595 ( .A(n_188), .Y(n_595) );
AOI22xp5_ASAP7_75t_SL g1353 ( .A1(n_189), .A2(n_251), .B1(n_1329), .B2(n_1332), .Y(n_1353) );
AOI22xp5_ASAP7_75t_L g1574 ( .A1(n_189), .A2(n_1575), .B1(n_1578), .B2(n_1667), .Y(n_1574) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_189), .A2(n_1581), .B1(n_1665), .B2(n_1666), .Y(n_1580) );
INVxp67_ASAP7_75t_L g1665 ( .A(n_189), .Y(n_1665) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_191), .A2(n_252), .B1(n_787), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g818 ( .A(n_191), .Y(n_818) );
INVxp33_ASAP7_75t_SL g1160 ( .A(n_192), .Y(n_1160) );
INVx1_ASAP7_75t_L g1550 ( .A(n_193), .Y(n_1550) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_194), .Y(n_801) );
INVxp33_ASAP7_75t_SL g1613 ( .A(n_195), .Y(n_1613) );
OAI211xp5_ASAP7_75t_L g837 ( .A1(n_196), .A2(n_838), .B(n_842), .C(n_847), .Y(n_837) );
INVx1_ASAP7_75t_L g905 ( .A(n_196), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_197), .A2(n_233), .B1(n_957), .B2(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1090 ( .A(n_197), .Y(n_1090) );
INVx1_ASAP7_75t_L g1084 ( .A(n_198), .Y(n_1084) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_199), .Y(n_657) );
INVx1_ASAP7_75t_L g1306 ( .A(n_200), .Y(n_1306) );
INVx1_ASAP7_75t_L g1603 ( .A(n_203), .Y(n_1603) );
AO221x2_ASAP7_75t_L g1423 ( .A1(n_204), .A2(n_206), .B1(n_1388), .B2(n_1424), .C(n_1425), .Y(n_1423) );
INVx1_ASAP7_75t_L g935 ( .A(n_205), .Y(n_935) );
INVx1_ASAP7_75t_L g1275 ( .A(n_207), .Y(n_1275) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_208), .A2(n_209), .B1(n_977), .B2(n_1061), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1086 ( .A1(n_208), .A2(n_209), .B1(n_535), .B2(n_994), .C(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g302 ( .A(n_210), .Y(n_302) );
INVx2_ASAP7_75t_L g414 ( .A(n_210), .Y(n_414) );
INVxp33_ASAP7_75t_SL g1124 ( .A(n_212), .Y(n_1124) );
OR2x2_ASAP7_75t_L g636 ( .A(n_213), .B(n_393), .Y(n_636) );
CKINVDCx14_ASAP7_75t_R g1427 ( .A(n_214), .Y(n_1427) );
INVx1_ASAP7_75t_L g1549 ( .A(n_215), .Y(n_1549) );
INVx1_ASAP7_75t_L g623 ( .A(n_216), .Y(n_623) );
INVx1_ASAP7_75t_L g881 ( .A(n_217), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_218), .A2(n_566), .B1(n_632), .B2(n_633), .Y(n_565) );
INVx1_ASAP7_75t_L g633 ( .A(n_218), .Y(n_633) );
INVxp67_ASAP7_75t_SL g1116 ( .A(n_219), .Y(n_1116) );
INVxp33_ASAP7_75t_SL g1176 ( .A(n_220), .Y(n_1176) );
INVx1_ASAP7_75t_L g748 ( .A(n_221), .Y(n_748) );
INVx1_ASAP7_75t_L g601 ( .A(n_222), .Y(n_601) );
INVx1_ASAP7_75t_L g980 ( .A(n_224), .Y(n_980) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_225), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g1313 ( .A(n_226), .Y(n_1313) );
INVx1_ASAP7_75t_L g404 ( .A(n_227), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_228), .Y(n_508) );
INVx1_ASAP7_75t_L g983 ( .A(n_229), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_230), .Y(n_380) );
INVx1_ASAP7_75t_L g819 ( .A(n_231), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_232), .Y(n_791) );
INVx1_ASAP7_75t_L g1096 ( .A(n_233), .Y(n_1096) );
INVx1_ASAP7_75t_L g1074 ( .A(n_234), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_236), .A2(n_241), .B1(n_594), .B2(n_793), .Y(n_792) );
OAI221xp5_ASAP7_75t_L g815 ( .A1(n_236), .A2(n_241), .B1(n_434), .B2(n_440), .C(n_444), .Y(n_815) );
INVx1_ASAP7_75t_L g599 ( .A(n_238), .Y(n_599) );
INVx1_ASAP7_75t_L g511 ( .A(n_239), .Y(n_511) );
INVx1_ASAP7_75t_L g524 ( .A(n_240), .Y(n_524) );
INVx1_ASAP7_75t_L g585 ( .A(n_242), .Y(n_585) );
INVx1_ASAP7_75t_L g809 ( .A(n_243), .Y(n_809) );
INVx1_ASAP7_75t_L g718 ( .A(n_244), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_244), .A2(n_262), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g1002 ( .A(n_245), .Y(n_1002) );
INVx1_ASAP7_75t_L g1022 ( .A(n_247), .Y(n_1022) );
INVx1_ASAP7_75t_L g1222 ( .A(n_248), .Y(n_1222) );
CKINVDCx5p33_ASAP7_75t_R g1555 ( .A(n_250), .Y(n_1555) );
INVx1_ASAP7_75t_L g822 ( .A(n_252), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_253), .Y(n_1073) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_254), .Y(n_875) );
INVx2_ASAP7_75t_L g299 ( .A(n_255), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_256), .Y(n_518) );
INVx1_ASAP7_75t_L g1106 ( .A(n_257), .Y(n_1106) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_258), .A2(n_333), .B(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g421 ( .A(n_258), .Y(n_421) );
INVx1_ASAP7_75t_L g540 ( .A(n_259), .Y(n_540) );
INVx1_ASAP7_75t_L g645 ( .A(n_260), .Y(n_645) );
INVx1_ASAP7_75t_L g660 ( .A(n_261), .Y(n_660) );
INVx1_ASAP7_75t_L g715 ( .A(n_262), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_263), .Y(n_936) );
INVx1_ASAP7_75t_L g810 ( .A(n_265), .Y(n_810) );
INVx1_ASAP7_75t_L g1233 ( .A(n_266), .Y(n_1233) );
INVxp67_ASAP7_75t_L g1004 ( .A(n_267), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_268), .Y(n_1072) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_269), .Y(n_721) );
INVx1_ASAP7_75t_L g1023 ( .A(n_270), .Y(n_1023) );
INVx1_ASAP7_75t_L g1237 ( .A(n_271), .Y(n_1237) );
CKINVDCx20_ASAP7_75t_R g1308 ( .A(n_272), .Y(n_1308) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_273), .A2(n_655), .B(n_656), .C(n_659), .Y(n_654) );
BUFx3_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
INVx1_ASAP7_75t_L g326 ( .A(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g320 ( .A(n_275), .Y(n_320) );
BUFx3_ASAP7_75t_L g325 ( .A(n_275), .Y(n_325) );
INVx1_ASAP7_75t_L g459 ( .A(n_276), .Y(n_459) );
INVx1_ASAP7_75t_L g532 ( .A(n_277), .Y(n_532) );
INVx1_ASAP7_75t_L g570 ( .A(n_278), .Y(n_570) );
INVx1_ASAP7_75t_L g1139 ( .A(n_279), .Y(n_1139) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_280), .Y(n_1173) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_303), .B(n_1291), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x4_ASAP7_75t_L g1577 ( .A(n_285), .B(n_291), .Y(n_1577) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g1573 ( .A(n_286), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_286), .B(n_288), .Y(n_1670) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_288), .B(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x6_ASAP7_75t_L g1610 ( .A(n_293), .B(n_399), .Y(n_1610) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g671 ( .A(n_294), .B(n_302), .Y(n_671) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g448 ( .A(n_295), .B(n_449), .Y(n_448) );
INVx8_ASAP7_75t_L g1602 ( .A(n_296), .Y(n_1602) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x2_ASAP7_75t_L g394 ( .A(n_297), .B(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g463 ( .A(n_297), .Y(n_463) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_297), .Y(n_559) );
INVx2_ASAP7_75t_SL g612 ( .A(n_297), .Y(n_612) );
INVx2_ASAP7_75t_SL g874 ( .A(n_297), .Y(n_874) );
INVx1_ASAP7_75t_L g1012 ( .A(n_297), .Y(n_1012) );
OR2x6_ASAP7_75t_L g1605 ( .A(n_297), .B(n_1586), .Y(n_1605) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_L g409 ( .A(n_299), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g419 ( .A(n_299), .Y(n_419) );
AND2x2_ASAP7_75t_L g425 ( .A(n_299), .B(n_300), .Y(n_425) );
INVx2_ASAP7_75t_L g430 ( .A(n_299), .Y(n_430) );
INVx1_ASAP7_75t_L g469 ( .A(n_299), .Y(n_469) );
INVx2_ASAP7_75t_L g410 ( .A(n_300), .Y(n_410) );
INVx1_ASAP7_75t_L g432 ( .A(n_300), .Y(n_432) );
INVx1_ASAP7_75t_L g438 ( .A(n_300), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_300), .B(n_430), .Y(n_454) );
INVx1_ASAP7_75t_L g468 ( .A(n_300), .Y(n_468) );
AND2x4_ASAP7_75t_L g1595 ( .A(n_301), .B(n_438), .Y(n_1595) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_1109), .B2(n_1110), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
XNOR2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_707), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_563), .B2(n_564), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_486), .B2(n_487), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
XNOR2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g1425 ( .A1(n_312), .A2(n_1426), .B1(n_1427), .B2(n_1428), .Y(n_1425) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_401), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_387), .B1(n_391), .B2(n_392), .Y(n_314) );
NAND4xp25_ASAP7_75t_L g315 ( .A(n_316), .B(n_355), .C(n_373), .D(n_383), .Y(n_315) );
AOI322xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_327), .A3(n_332), .B1(n_343), .B2(n_350), .C1(n_351), .C2(n_354), .Y(n_316) );
BUFx3_ASAP7_75t_L g1250 ( .A(n_318), .Y(n_1250) );
BUFx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_319), .Y(n_386) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_319), .Y(n_499) );
BUFx2_ASAP7_75t_L g515 ( .A(n_319), .Y(n_515) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_319), .Y(n_584) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_319), .Y(n_588) );
BUFx2_ASAP7_75t_L g796 ( .A(n_319), .Y(n_796) );
INVx2_ASAP7_75t_SL g914 ( .A(n_319), .Y(n_914) );
AND2x6_ASAP7_75t_L g1619 ( .A(n_319), .B(n_1620), .Y(n_1619) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g379 ( .A(n_320), .Y(n_379) );
AND2x2_ASAP7_75t_L g331 ( .A(n_321), .B(n_325), .Y(n_331) );
INVx2_ASAP7_75t_L g336 ( .A(n_321), .Y(n_336) );
BUFx2_ASAP7_75t_L g1157 ( .A(n_322), .Y(n_1157) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x6_ASAP7_75t_L g921 ( .A(n_323), .B(n_916), .Y(n_921) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_324), .Y(n_505) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_324), .Y(n_644) );
INVx1_ASAP7_75t_L g1658 ( .A(n_324), .Y(n_1658) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx2_ASAP7_75t_L g337 ( .A(n_325), .Y(n_337) );
INVx1_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g1628 ( .A1(n_328), .A2(n_1594), .B1(n_1596), .B2(n_1629), .C1(n_1630), .C2(n_1633), .Y(n_1628) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g577 ( .A(n_329), .Y(n_577) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_330), .Y(n_498) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_330), .Y(n_777) );
INVx1_ASAP7_75t_L g909 ( .A(n_330), .Y(n_909) );
AND2x4_ASAP7_75t_L g1635 ( .A(n_330), .B(n_1636), .Y(n_1635) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
AND2x2_ASAP7_75t_L g918 ( .A(n_333), .B(n_915), .Y(n_918) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g968 ( .A(n_334), .Y(n_968) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g400 ( .A(n_335), .B(n_344), .Y(n_400) );
INVx6_ASAP7_75t_L g503 ( .A(n_335), .Y(n_503) );
AND2x4_ASAP7_75t_L g1623 ( .A(n_335), .B(n_1624), .Y(n_1623) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g353 ( .A(n_336), .Y(n_353) );
INVx1_ASAP7_75t_L g349 ( .A(n_337), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_SL g521 ( .A(n_339), .Y(n_521) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_339), .Y(n_760) );
INVx1_ASAP7_75t_L g788 ( .A(n_339), .Y(n_788) );
AND2x4_ASAP7_75t_L g902 ( .A(n_339), .B(n_399), .Y(n_902) );
INVx2_ASAP7_75t_L g1149 ( .A(n_339), .Y(n_1149) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AND2x4_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g367 ( .A(n_341), .B(n_342), .Y(n_367) );
INVx1_ASAP7_75t_L g1616 ( .A(n_341), .Y(n_1616) );
INVx1_ASAP7_75t_L g1621 ( .A(n_341), .Y(n_1621) );
HB1xp67_ASAP7_75t_L g1625 ( .A(n_341), .Y(n_1625) );
INVx1_ASAP7_75t_L g1638 ( .A(n_342), .Y(n_1638) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_343), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVx2_ASAP7_75t_L g750 ( .A(n_343), .Y(n_750) );
INVx2_ASAP7_75t_SL g976 ( .A(n_343), .Y(n_976) );
INVx1_ASAP7_75t_L g1061 ( .A(n_343), .Y(n_1061) );
INVx1_ASAP7_75t_L g1559 ( .A(n_343), .Y(n_1559) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
AND2x4_ASAP7_75t_L g351 ( .A(n_344), .B(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
AND2x2_ASAP7_75t_L g512 ( .A(n_344), .B(n_352), .Y(n_512) );
AND2x4_ASAP7_75t_L g593 ( .A(n_344), .B(n_347), .Y(n_593) );
INVx1_ASAP7_75t_L g776 ( .A(n_344), .Y(n_776) );
NAND2x1p5_ASAP7_75t_L g892 ( .A(n_344), .B(n_474), .Y(n_892) );
AND2x2_ASAP7_75t_L g978 ( .A(n_344), .B(n_352), .Y(n_978) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g890 ( .A(n_348), .Y(n_890) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g1632 ( .A(n_349), .Y(n_1632) );
INVx2_ASAP7_75t_SL g594 ( .A(n_351), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_351), .A2(n_593), .B1(n_657), .B2(n_658), .Y(n_656) );
AOI222xp33_ASAP7_75t_SL g1016 ( .A1(n_351), .A2(n_1017), .B1(n_1019), .B2(n_1020), .C1(n_1022), .C2(n_1023), .Y(n_1016) );
INVx2_ASAP7_75t_L g894 ( .A(n_352), .Y(n_894) );
BUFx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x6_ASAP7_75t_L g1633 ( .A(n_353), .B(n_1621), .Y(n_1633) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B1(n_361), .B2(n_368), .C(n_371), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_356), .A2(n_371), .B1(n_496), .B2(n_497), .C(n_500), .Y(n_495) );
INVx2_ASAP7_75t_SL g574 ( .A(n_356), .Y(n_574) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_356), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g794 ( .A1(n_356), .A2(n_371), .B1(n_795), .B2(n_797), .C(n_801), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_356), .A2(n_358), .B1(n_371), .B2(n_1013), .C(n_1025), .Y(n_1024) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
BUFx4f_ASAP7_75t_L g363 ( .A(n_357), .Y(n_363) );
AND2x4_ASAP7_75t_L g371 ( .A(n_357), .B(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g768 ( .A(n_357), .Y(n_768) );
INVx1_ASAP7_75t_L g1041 ( .A(n_357), .Y(n_1041) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_357), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1067 ( .A(n_357), .Y(n_1067) );
AND2x4_ASAP7_75t_L g385 ( .A(n_358), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g583 ( .A(n_358), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g376 ( .A(n_359), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g382 ( .A(n_359), .B(n_370), .Y(n_382) );
OR2x2_ASAP7_75t_L g916 ( .A(n_359), .B(n_412), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g954 ( .A1(n_359), .A2(n_955), .B(n_958), .C(n_959), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_360), .A2(n_374), .B1(n_479), .B2(n_480), .Y(n_478) );
BUFx3_ASAP7_75t_L g1034 ( .A(n_362), .Y(n_1034) );
INVx2_ASAP7_75t_L g1154 ( .A(n_362), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_363), .A2(n_913), .B1(n_939), .B2(n_941), .Y(n_958) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x6_ASAP7_75t_L g1230 ( .A(n_366), .B(n_389), .Y(n_1230) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g579 ( .A(n_367), .Y(n_579) );
INVx2_ASAP7_75t_SL g652 ( .A(n_367), .Y(n_652) );
INVx1_ASAP7_75t_L g897 ( .A(n_367), .Y(n_897) );
INVx1_ASAP7_75t_L g974 ( .A(n_367), .Y(n_974) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g800 ( .A(n_370), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_371), .A2(n_573), .B1(n_575), .B2(n_576), .C(n_580), .Y(n_572) );
INVx1_ASAP7_75t_L g653 ( .A(n_371), .Y(n_653) );
INVx1_ASAP7_75t_L g959 ( .A(n_371), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_371), .A2(n_762), .B1(n_1063), .B2(n_1068), .C(n_1070), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_380), .B2(n_381), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_375), .A2(n_381), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_375), .A2(n_381), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_375), .A2(n_381), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_375), .A2(n_381), .B1(n_803), .B2(n_804), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_375), .A2(n_381), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_375), .A2(n_381), .B1(n_1159), .B2(n_1160), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_375), .A2(n_381), .B1(n_1215), .B2(n_1216), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1569 ( .A1(n_375), .A2(n_381), .B1(n_1552), .B2(n_1553), .Y(n_1569) );
INVx6_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g641 ( .A(n_377), .Y(n_641) );
INVx1_ASAP7_75t_L g759 ( .A(n_377), .Y(n_759) );
INVx1_ASAP7_75t_L g1027 ( .A(n_377), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1232 ( .A(n_377), .Y(n_1232) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g650 ( .A(n_378), .B(n_379), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_380), .A2(n_384), .B1(n_451), .B2(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_385), .B(n_523), .Y(n_522) );
AOI211xp5_ASAP7_75t_SL g747 ( .A1(n_385), .A2(n_748), .B(n_749), .C(n_752), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_385), .A2(n_1053), .B1(n_1056), .B2(n_1059), .C(n_1060), .Y(n_1052) );
AOI21xp33_ASAP7_75t_SL g1141 ( .A1(n_385), .A2(n_1142), .B(n_1143), .Y(n_1141) );
AOI211xp5_ASAP7_75t_L g1198 ( .A1(n_385), .A2(n_1199), .B(n_1200), .C(n_1202), .Y(n_1198) );
AOI211xp5_ASAP7_75t_L g1557 ( .A1(n_385), .A2(n_1549), .B(n_1558), .C(n_1560), .Y(n_1557) );
INVx2_ASAP7_75t_SL g1240 ( .A(n_386), .Y(n_1240) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_387), .A2(n_392), .B1(n_568), .B2(n_595), .Y(n_567) );
INVx2_ASAP7_75t_L g1161 ( .A(n_387), .Y(n_1161) );
CKINVDCx8_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g667 ( .A(n_389), .Y(n_667) );
AND2x4_ASAP7_75t_L g670 ( .A(n_389), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g689 ( .A(n_389), .B(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g728 ( .A(n_389), .B(n_671), .Y(n_728) );
OR2x2_ASAP7_75t_L g896 ( .A(n_389), .B(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x6_ASAP7_75t_L g447 ( .A(n_390), .B(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g493 ( .A(n_390), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_392), .A2(n_667), .B1(n_784), .B2(n_805), .Y(n_783) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx5_ASAP7_75t_L g525 ( .A(n_393), .Y(n_525) );
INVx1_ASAP7_75t_L g1075 ( .A(n_393), .Y(n_1075) );
INVx1_ASAP7_75t_L g1195 ( .A(n_393), .Y(n_1195) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_397), .Y(n_393) );
INVx3_ASAP7_75t_L g439 ( .A(n_395), .Y(n_439) );
INVx1_ASAP7_75t_L g859 ( .A(n_396), .Y(n_859) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x6_ASAP7_75t_L g882 ( .A(n_398), .B(n_883), .Y(n_882) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_400), .B(n_980), .Y(n_979) );
INVx2_ASAP7_75t_L g1018 ( .A(n_400), .Y(n_1018) );
NOR3xp33_ASAP7_75t_SL g401 ( .A(n_402), .B(n_433), .C(n_446), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_420), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_415), .B2(n_416), .Y(n_403) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g529 ( .A(n_406), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_406), .A2(n_416), .B1(n_809), .B2(n_810), .Y(n_808) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_406), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1080 ( .A(n_406), .Y(n_1080) );
BUFx2_ASAP7_75t_L g1120 ( .A(n_406), .Y(n_1120) );
BUFx2_ASAP7_75t_L g1177 ( .A(n_406), .Y(n_1177) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .Y(n_406) );
BUFx3_ASAP7_75t_L g485 ( .A(n_407), .Y(n_485) );
INVx2_ASAP7_75t_L g622 ( .A(n_407), .Y(n_622) );
INVx1_ASAP7_75t_L g868 ( .A(n_407), .Y(n_868) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g552 ( .A(n_408), .Y(n_552) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_408), .Y(n_851) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g458 ( .A(n_409), .Y(n_458) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_409), .Y(n_732) );
INVx1_ASAP7_75t_L g1590 ( .A(n_409), .Y(n_1590) );
AND2x4_ASAP7_75t_L g418 ( .A(n_410), .B(n_419), .Y(n_418) );
AND2x6_ASAP7_75t_L g416 ( .A(n_411), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g422 ( .A(n_411), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g427 ( .A(n_411), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g533 ( .A(n_411), .B(n_428), .Y(n_533) );
AND2x2_ASAP7_75t_L g600 ( .A(n_411), .B(n_552), .Y(n_600) );
AND2x2_ASAP7_75t_L g602 ( .A(n_411), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g725 ( .A(n_411), .B(n_428), .Y(n_725) );
AND2x2_ASAP7_75t_L g814 ( .A(n_411), .B(n_428), .Y(n_814) );
AND2x2_ASAP7_75t_L g947 ( .A(n_411), .B(n_886), .Y(n_947) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_411), .B(n_428), .Y(n_1085) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
INVx2_ASAP7_75t_L g841 ( .A(n_413), .Y(n_841) );
AND2x2_ASAP7_75t_L g844 ( .A(n_413), .B(n_429), .Y(n_844) );
AND2x4_ASAP7_75t_L g863 ( .A(n_413), .B(n_688), .Y(n_863) );
INVx1_ASAP7_75t_L g449 ( .A(n_414), .Y(n_449) );
INVx1_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_416), .A2(n_518), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_416), .A2(n_529), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_416), .A2(n_1079), .B1(n_1080), .B2(n_1081), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_416), .A2(n_1119), .B1(n_1120), .B2(n_1121), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_416), .A2(n_1176), .B1(n_1177), .B2(n_1178), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_416), .A2(n_1177), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_417), .B(n_439), .Y(n_445) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_418), .Y(n_603) );
BUFx3_ASAP7_75t_L g675 ( .A(n_418), .Y(n_675) );
BUFx2_ASAP7_75t_L g698 ( .A(n_418), .Y(n_698) );
BUFx6f_ASAP7_75t_L g1593 ( .A(n_418), .Y(n_1593) );
AND2x4_ASAP7_75t_L g1607 ( .A(n_418), .B(n_1608), .Y(n_1607) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_426), .B2(n_427), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_422), .A2(n_516), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_422), .A2(n_427), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_422), .A2(n_533), .B1(n_700), .B2(n_701), .C(n_702), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_422), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_422), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g1043 ( .A(n_422), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_422), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_422), .A2(n_814), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_422), .A2(n_533), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_422), .A2(n_533), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
BUFx2_ASAP7_75t_L g673 ( .A(n_423), .Y(n_673) );
BUFx3_ASAP7_75t_L g742 ( .A(n_423), .Y(n_742) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g886 ( .A(n_424), .Y(n_886) );
INVx2_ASAP7_75t_L g1645 ( .A(n_424), .Y(n_1645) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_425), .Y(n_688) );
INVx1_ASAP7_75t_L g950 ( .A(n_427), .Y(n_950) );
INVx1_ASAP7_75t_L g993 ( .A(n_427), .Y(n_993) );
INVx2_ASAP7_75t_SL g738 ( .A(n_428), .Y(n_738) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g678 ( .A(n_429), .Y(n_678) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_429), .Y(n_849) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_429), .Y(n_1131) );
AND2x4_ASAP7_75t_L g1585 ( .A(n_429), .B(n_1586), .Y(n_1585) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g443 ( .A(n_430), .Y(n_443) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g536 ( .A(n_435), .Y(n_536) );
NAND2x1_ASAP7_75t_SL g435 ( .A(n_436), .B(n_439), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g856 ( .A(n_436), .B(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_438), .Y(n_693) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_439), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g692 ( .A(n_439), .B(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g694 ( .A(n_439), .B(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g697 ( .A(n_439), .B(n_698), .Y(n_697) );
BUFx4f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx4f_ASAP7_75t_L g994 ( .A(n_441), .Y(n_994) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x6_ASAP7_75t_L g860 ( .A(n_443), .B(n_858), .Y(n_860) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g537 ( .A(n_445), .Y(n_537) );
BUFx2_ASAP7_75t_L g1087 ( .A(n_445), .Y(n_1087) );
OAI33xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_450), .A3(n_460), .B1(n_471), .B2(n_478), .B3(n_483), .Y(n_446) );
OAI33xp33_ASAP7_75t_L g538 ( .A1(n_447), .A2(n_471), .A3(n_539), .B1(n_543), .B2(n_554), .B3(n_556), .Y(n_538) );
OAI33xp33_ASAP7_75t_L g609 ( .A1(n_447), .A2(n_610), .A3(n_618), .B1(n_624), .B2(n_628), .B3(n_630), .Y(n_609) );
OAI33xp33_ASAP7_75t_L g816 ( .A1(n_447), .A2(n_471), .A3(n_817), .B1(n_820), .B2(n_823), .B3(n_826), .Y(n_816) );
OAI33xp33_ASAP7_75t_L g1088 ( .A1(n_447), .A2(n_630), .A3(n_1089), .B1(n_1093), .B2(n_1098), .B3(n_1104), .Y(n_1088) );
OAI33xp33_ASAP7_75t_L g1536 ( .A1(n_447), .A2(n_471), .A3(n_1537), .B1(n_1542), .B2(n_1547), .B3(n_1551), .Y(n_1536) );
INVx1_ASAP7_75t_L g1586 ( .A(n_449), .Y(n_1586) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_455), .B1(n_456), .B2(n_459), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_451), .A2(n_551), .B1(n_821), .B2(n_822), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_451), .A2(n_791), .B1(n_804), .B2(n_824), .Y(n_823) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g942 ( .A(n_452), .Y(n_942) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_453), .Y(n_626) );
INVx1_ASAP7_75t_L g1101 ( .A(n_453), .Y(n_1101) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g547 ( .A(n_454), .Y(n_547) );
BUFx2_ASAP7_75t_L g866 ( .A(n_454), .Y(n_866) );
INVx1_ASAP7_75t_L g1648 ( .A(n_456), .Y(n_1648) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g627 ( .A(n_457), .Y(n_627) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g684 ( .A(n_458), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B1(n_465), .B2(n_470), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g479 ( .A(n_462), .Y(n_479) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g817 ( .A1(n_465), .A2(n_479), .B1(n_818), .B2(n_819), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_465), .A2(n_873), .B1(n_935), .B2(n_936), .Y(n_934) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g561 ( .A(n_466), .Y(n_561) );
BUFx3_ASAP7_75t_L g629 ( .A(n_466), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g937 ( .A1(n_466), .A2(n_559), .B1(n_938), .B2(n_939), .Y(n_937) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
AND2x2_ASAP7_75t_L g482 ( .A(n_468), .B(n_469), .Y(n_482) );
INVx1_ASAP7_75t_L g696 ( .A(n_469), .Y(n_696) );
CKINVDCx8_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g1646 ( .A(n_472), .B(n_1647), .C(n_1649), .Y(n_1646) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx6_ASAP7_75t_L g631 ( .A(n_473), .Y(n_631) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g690 ( .A(n_475), .Y(n_690) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g1599 ( .A(n_476), .Y(n_1599) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_479), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_539) );
OAI22xp33_ASAP7_75t_L g826 ( .A1(n_479), .A2(n_614), .B1(n_801), .B2(n_803), .Y(n_826) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g616 ( .A(n_482), .Y(n_616) );
INVx3_ASAP7_75t_L g871 ( .A(n_482), .Y(n_871) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
XNOR2x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_562), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_526), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_494), .B1(n_524), .B2(n_525), .Y(n_489) );
AOI21xp5_ASAP7_75t_SL g1014 ( .A1(n_490), .A2(n_1015), .B(n_1042), .Y(n_1014) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI31xp33_ASAP7_75t_L g746 ( .A1(n_491), .A2(n_747), .A3(n_761), .B(n_778), .Y(n_746) );
AOI31xp33_ASAP7_75t_L g1556 ( .A1(n_491), .A2(n_1557), .A3(n_1563), .B(n_1569), .Y(n_1556) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI31xp33_ASAP7_75t_L g953 ( .A1(n_492), .A2(n_954), .A3(n_960), .B(n_975), .Y(n_953) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g879 ( .A(n_493), .Y(n_879) );
AND2x4_ASAP7_75t_L g1637 ( .A(n_493), .B(n_1638), .Y(n_1637) );
NAND5xp2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .C(n_509), .D(n_513), .E(n_522), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_496), .A2(n_507), .B1(n_557), .B2(n_560), .Y(n_556) );
HB1xp67_ASAP7_75t_L g1566 ( .A(n_498), .Y(n_1566) );
BUFx3_ASAP7_75t_L g1057 ( .A(n_499), .Y(n_1057) );
INVx2_ASAP7_75t_L g1065 ( .A(n_499), .Y(n_1065) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g520 ( .A(n_502), .Y(n_520) );
INVx4_ASAP7_75t_L g1055 ( .A(n_502), .Y(n_1055) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g772 ( .A(n_503), .Y(n_772) );
INVx1_ASAP7_75t_L g787 ( .A(n_503), .Y(n_787) );
INVx2_ASAP7_75t_L g956 ( .A(n_503), .Y(n_956) );
INVx1_ASAP7_75t_L g972 ( .A(n_503), .Y(n_972) );
INVx2_ASAP7_75t_SL g1148 ( .A(n_503), .Y(n_1148) );
INVx2_ASAP7_75t_L g1617 ( .A(n_503), .Y(n_1617) );
INVx1_ASAP7_75t_L g517 ( .A(n_504), .Y(n_517) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_504), .Y(n_773) );
INVx1_ASAP7_75t_L g1242 ( .A(n_504), .Y(n_1242) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_505), .Y(n_581) );
INVx1_ASAP7_75t_L g590 ( .A(n_505), .Y(n_590) );
BUFx6f_ASAP7_75t_L g957 ( .A(n_505), .Y(n_957) );
INVx2_ASAP7_75t_L g1028 ( .A(n_505), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_505), .Y(n_1030) );
AND2x6_ASAP7_75t_L g1627 ( .A(n_505), .B(n_1615), .Y(n_1627) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_508), .A2(n_523), .B1(n_551), .B2(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g751 ( .A(n_512), .Y(n_751) );
OAI221xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_516), .B1(n_517), .B2(n_518), .C(n_519), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_525), .A2(n_745), .B(n_746), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_525), .A2(n_1139), .B(n_1140), .Y(n_1138) );
AOI21xp33_ASAP7_75t_SL g1554 ( .A1(n_525), .A2(n_1555), .B(n_1556), .Y(n_1554) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_534), .C(n_538), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g608 ( .A(n_536), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_548), .B1(n_549), .B2(n_553), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g555 ( .A(n_545), .Y(n_555) );
INVx2_ASAP7_75t_L g1095 ( .A(n_545), .Y(n_1095) );
INVx2_ASAP7_75t_L g1548 ( .A(n_545), .Y(n_1548) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g620 ( .A(n_547), .Y(n_620) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g1643 ( .A(n_551), .Y(n_1643) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g680 ( .A(n_552), .Y(n_680) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_552), .Y(n_933) );
INVx1_ASAP7_75t_L g1007 ( .A(n_552), .Y(n_1007) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_559), .A2(n_570), .B1(n_575), .B2(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_559), .Y(n_1105) );
OAI22xp5_ASAP7_75t_SL g1009 ( .A1(n_560), .A2(n_1010), .B1(n_1011), .B2(n_1013), .Y(n_1009) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
XOR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_634), .Y(n_564) );
INVx1_ASAP7_75t_L g632 ( .A(n_566), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_596), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .C(n_582), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_571), .A2(n_585), .B1(n_625), .B2(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B1(n_586), .B2(n_587), .C(n_591), .Y(n_582) );
INVx1_ASAP7_75t_L g655 ( .A(n_583), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_583), .A2(n_786), .B1(n_789), .B2(n_791), .C(n_792), .Y(n_785) );
INVx1_ASAP7_75t_L g754 ( .A(n_584), .Y(n_754) );
INVx1_ASAP7_75t_L g766 ( .A(n_584), .Y(n_766) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g793 ( .A(n_593), .Y(n_793) );
INVx4_ASAP7_75t_L g1021 ( .A(n_593), .Y(n_1021) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_607), .C(n_609), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_604), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_598) );
INVx2_ASAP7_75t_L g703 ( .A(n_600), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_602), .Y(n_704) );
INVxp67_ASAP7_75t_L g951 ( .A(n_602), .Y(n_951) );
INVx2_ASAP7_75t_SL g734 ( .A(n_603), .Y(n_734) );
BUFx6f_ASAP7_75t_L g1193 ( .A(n_603), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B1(n_614), .B2(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x6_ASAP7_75t_L g877 ( .A(n_616), .B(n_858), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_616), .A2(n_873), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_616), .B(n_858), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g998 ( .A(n_620), .Y(n_998) );
INVx2_ASAP7_75t_SL g1267 ( .A(n_620), .Y(n_1267) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_629), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1089) );
OAI22xp33_ASAP7_75t_L g1104 ( .A1(n_629), .A2(n_1070), .B1(n_1072), .B2(n_1105), .Y(n_1104) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI33xp33_ASAP7_75t_L g726 ( .A1(n_631), .A2(n_727), .A3(n_729), .B1(n_735), .B2(n_739), .B3(n_741), .Y(n_726) );
INVx1_ASAP7_75t_L g945 ( .A(n_631), .Y(n_945) );
AOI33xp33_ASAP7_75t_L g1125 ( .A1(n_631), .A2(n_670), .A3(n_1126), .B1(n_1130), .B2(n_1134), .B3(n_1135), .Y(n_1125) );
AOI33xp33_ASAP7_75t_L g1182 ( .A1(n_631), .A2(n_1183), .A3(n_1185), .B1(n_1187), .B2(n_1189), .B3(n_1192), .Y(n_1182) );
INVx1_ASAP7_75t_L g706 ( .A(n_635), .Y(n_706) );
NAND4xp75_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .C(n_668), .D(n_699), .Y(n_635) );
OAI31xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_654), .A3(n_664), .B(n_665), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_643), .B2(n_645), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g899 ( .A(n_641), .Y(n_899) );
INVx2_ASAP7_75t_L g1244 ( .A(n_641), .Y(n_1244) );
INVx1_ASAP7_75t_L g1289 ( .A(n_641), .Y(n_1289) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx3_ASAP7_75t_L g755 ( .A(n_644), .Y(n_755) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_644), .Y(n_790) );
OAI21xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_651), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_648), .A2(n_872), .B1(n_875), .B2(n_899), .C(n_900), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_648), .A2(n_758), .B1(n_904), .B2(n_905), .C(n_906), .Y(n_903) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g661 ( .A(n_649), .Y(n_661) );
INVx1_ASAP7_75t_L g970 ( .A(n_649), .Y(n_970) );
INVx2_ASAP7_75t_L g1145 ( .A(n_649), .Y(n_1145) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g757 ( .A(n_650), .Y(n_757) );
INVx2_ASAP7_75t_L g923 ( .A(n_650), .Y(n_923) );
INVx1_ASAP7_75t_L g965 ( .A(n_650), .Y(n_965) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_650), .Y(n_1205) );
INVx1_ASAP7_75t_L g1236 ( .A(n_650), .Y(n_1236) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_657), .A2(n_658), .B1(n_692), .B2(n_694), .C(n_697), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B(n_662), .C(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI31xp33_ASAP7_75t_SL g1256 ( .A1(n_666), .A2(n_1257), .A3(n_1260), .B(n_1273), .Y(n_1256) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp67_ASAP7_75t_L g883 ( .A(n_667), .B(n_884), .Y(n_883) );
AND2x2_ASAP7_75t_SL g668 ( .A(n_669), .B(n_691), .Y(n_668) );
AOI33xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .A3(n_676), .B1(n_681), .B2(n_685), .B3(n_689), .Y(n_669) );
BUFx2_ASAP7_75t_SL g876 ( .A(n_671), .Y(n_876) );
INVx1_ASAP7_75t_L g1264 ( .A(n_671), .Y(n_1264) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_674), .Y(n_1186) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x4_ASAP7_75t_L g839 ( .A(n_675), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g1642 ( .A(n_678), .Y(n_1642) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g825 ( .A(n_680), .Y(n_825) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g846 ( .A(n_684), .B(n_840), .Y(n_846) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_SL g736 ( .A(n_687), .Y(n_736) );
INVx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
BUFx6f_ASAP7_75t_L g853 ( .A(n_688), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_690), .Y(n_854) );
INVx1_ASAP7_75t_L g1278 ( .A(n_690), .Y(n_1278) );
INVx1_ASAP7_75t_L g717 ( .A(n_692), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_692), .A2(n_694), .B1(n_697), .B2(n_982), .C(n_983), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g1046 ( .A1(n_692), .A2(n_697), .B(n_1022), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_692), .A2(n_694), .B1(n_697), .B2(n_1116), .C(n_1117), .Y(n_1115) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_692), .A2(n_1170), .B1(n_1172), .B2(n_1173), .C(n_1174), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_693), .B(n_885), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_694), .Y(n_714) );
INVx1_ASAP7_75t_L g1171 ( .A(n_694), .Y(n_1171) );
AND2x4_ASAP7_75t_L g1597 ( .A(n_695), .B(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_697), .A2(n_714), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_713) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_697), .Y(n_1174) );
INVx1_ASAP7_75t_L g1129 ( .A(n_698), .Y(n_1129) );
XNOR2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_831), .Y(n_707) );
AO22x2_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_781), .B1(n_829), .B2(n_830), .Y(n_708) );
INVx1_ASAP7_75t_L g830 ( .A(n_709), .Y(n_830) );
XNOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
AND2x4_ASAP7_75t_L g711 ( .A(n_712), .B(n_744), .Y(n_711) );
AND4x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_719), .C(n_722), .D(n_726), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_721), .A2(n_723), .B1(n_757), .B2(n_758), .C(n_760), .Y(n_756) );
BUFx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g1184 ( .A(n_728), .Y(n_1184) );
NAND3xp33_ASAP7_75t_L g1640 ( .A(n_728), .B(n_1641), .C(n_1644), .Y(n_1640) );
INVx2_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_731), .A2(n_997), .B1(n_998), .B2(n_999), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1551 ( .A1(n_731), .A2(n_1011), .B1(n_1552), .B2(n_1553), .Y(n_1551) );
INVx4_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx3_ASAP7_75t_L g740 ( .A(n_732), .Y(n_740) );
INVx2_ASAP7_75t_SL g944 ( .A(n_732), .Y(n_944) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_732), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1191 ( .A(n_732), .Y(n_1191) );
INVx2_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g743 ( .A(n_734), .Y(n_743) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g1097 ( .A(n_740), .Y(n_1097) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_754), .B(n_916), .Y(n_1290) );
OAI221xp5_ASAP7_75t_L g1562 ( .A1(n_757), .A2(n_760), .B1(n_899), .B2(n_1531), .C(n_1533), .Y(n_1562) );
OAI221xp5_ASAP7_75t_L g1203 ( .A1(n_758), .A2(n_1178), .B1(n_1180), .B2(n_1204), .C(n_1206), .Y(n_1203) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_764), .B2(n_769), .C(n_774), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_762), .A2(n_774), .B1(n_1151), .B2(n_1152), .C(n_1156), .Y(n_1150) );
AOI221xp5_ASAP7_75t_L g1207 ( .A1(n_762), .A2(n_774), .B1(n_1208), .B2(n_1211), .C(n_1213), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1563 ( .A1(n_762), .A2(n_774), .B1(n_1550), .B2(n_1564), .C(n_1567), .Y(n_1563) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
BUFx2_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
BUFx6f_ASAP7_75t_L g1662 ( .A(n_772), .Y(n_1662) );
AND2x4_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_776), .B(n_894), .Y(n_1201) );
BUFx6f_ASAP7_75t_L g1655 ( .A(n_777), .Y(n_1655) );
INVx3_ASAP7_75t_L g829 ( .A(n_781), .Y(n_829) );
INVx1_ASAP7_75t_L g827 ( .A(n_782), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_806), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_794), .C(n_802), .Y(n_784) );
INVx2_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1037 ( .A(n_799), .Y(n_1037) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
BUFx2_ASAP7_75t_L g1568 ( .A(n_800), .Y(n_1568) );
NOR3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_815), .C(n_816), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_811), .Y(n_807) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_986), .B1(n_987), .B2(n_1107), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1108 ( .A(n_833), .Y(n_1108) );
XNOR2x1_ASAP7_75t_L g833 ( .A(n_834), .B(n_926), .Y(n_833) );
INVx1_ASAP7_75t_L g924 ( .A(n_835), .Y(n_924) );
NAND4xp25_ASAP7_75t_L g835 ( .A(n_836), .B(n_880), .C(n_887), .D(n_911), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_861), .B(n_878), .Y(n_836) );
INVx8_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_842) );
INVx3_ASAP7_75t_L g1258 ( .A(n_844), .Y(n_1258) );
INVx3_ASAP7_75t_L g1259 ( .A(n_846), .Y(n_1259) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_852), .B(n_855), .Y(n_847) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_849), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1545 ( .A(n_850), .Y(n_1545) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx3_ASAP7_75t_L g1103 ( .A(n_851), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_853), .Y(n_1127) );
INVx1_ASAP7_75t_L g1137 ( .A(n_853), .Y(n_1137) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g885 ( .A(n_858), .Y(n_885) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
CKINVDCx11_ASAP7_75t_R g1283 ( .A(n_860), .Y(n_1283) );
CKINVDCx6p67_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_865), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
BUFx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g1006 ( .A(n_866), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_873), .B2(n_875), .C(n_876), .Y(n_870) );
BUFx2_ASAP7_75t_L g1262 ( .A(n_871), .Y(n_1262) );
INVx1_ASAP7_75t_L g1540 ( .A(n_871), .Y(n_1540) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_873), .A2(n_1233), .B1(n_1237), .B2(n_1262), .C(n_1263), .Y(n_1261) );
INVx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx8_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g1050 ( .A(n_879), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_882), .B(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
BUFx2_ASAP7_75t_L g1650 ( .A(n_886), .Y(n_1650) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_895), .C(n_907), .Y(n_887) );
INVx2_ASAP7_75t_L g1254 ( .A(n_889), .Y(n_1254) );
NAND2x1p5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
INVx2_ASAP7_75t_SL g891 ( .A(n_892), .Y(n_891) );
OR2x6_ASAP7_75t_L g893 ( .A(n_892), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g910 ( .A(n_892), .Y(n_910) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_892), .B(n_894), .Y(n_1255) );
OAI22xp5_ASAP7_75t_SL g895 ( .A1(n_896), .A2(n_898), .B1(n_901), .B2(n_903), .Y(n_895) );
OAI22xp33_ASAP7_75t_L g1227 ( .A1(n_901), .A2(n_1228), .B1(n_1231), .B2(n_1243), .Y(n_1227) );
INVx4_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
BUFx4f_ASAP7_75t_L g1664 ( .A(n_902), .Y(n_1664) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_907), .Y(n_1251) );
AND2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_910), .Y(n_907) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_908), .Y(n_1155) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_917), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_913), .B(n_915), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g1209 ( .A(n_914), .Y(n_1209) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
OR2x6_ASAP7_75t_L g922 ( .A(n_916), .B(n_923), .Y(n_922) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_916), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1247 ( .A(n_923), .Y(n_1247) );
INVx1_ASAP7_75t_SL g985 ( .A(n_927), .Y(n_985) );
NAND4xp75_ASAP7_75t_L g927 ( .A(n_928), .B(n_948), .C(n_953), .D(n_981), .Y(n_927) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
OAI211xp5_ASAP7_75t_L g969 ( .A1(n_936), .A2(n_970), .B(n_971), .C(n_973), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_938), .A2(n_943), .B1(n_956), .B2(n_957), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B1(n_943), .B2(n_944), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g1274 ( .A1(n_944), .A2(n_1095), .B1(n_1275), .B2(n_1276), .C(n_1277), .Y(n_1274) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NOR2x1_ASAP7_75t_L g948 ( .A(n_949), .B(n_952), .Y(n_948) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_956), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_969), .Y(n_960) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_963), .B(n_966), .C(n_967), .Y(n_961) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_972), .Y(n_1212) );
INVx3_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1337 ( .A1(n_984), .A2(n_1302), .B1(n_1311), .B2(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
XNOR2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_1047), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
AND2x2_ASAP7_75t_L g990 ( .A(n_991), .B(n_1014), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_995), .Y(n_991) );
OAI221xp5_ASAP7_75t_SL g1029 ( .A1(n_999), .A2(n_1002), .B1(n_1026), .B2(n_1030), .C(n_1031), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1007), .B2(n_1008), .Y(n_1003) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1007), .Y(n_1270) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1012), .Y(n_1091) );
NAND4xp25_ASAP7_75t_SL g1015 ( .A(n_1016), .B(n_1024), .C(n_1029), .D(n_1032), .Y(n_1015) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1028), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1035), .B1(n_1036), .B2(n_1038), .C(n_1039), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1041), .Y(n_1210) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
XNOR2x1_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1106), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1076), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1051), .B1(n_1074), .B2(n_1075), .Y(n_1049) );
NAND3xp33_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1062), .C(n_1071), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_1059), .A2(n_1073), .B1(n_1099), .B2(n_1102), .Y(n_1098) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
NOR3xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1086), .C(n_1088), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1082), .Y(n_1077) );
OAI22xp5_ASAP7_75t_SL g1093 ( .A1(n_1094), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1542 ( .A1(n_1095), .A2(n_1543), .B1(n_1544), .B2(n_1546), .Y(n_1542) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1537 ( .A1(n_1105), .A2(n_1538), .B1(n_1539), .B2(n_1541), .Y(n_1537) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
XOR2xp5_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1219), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1163), .B1(n_1164), .B2(n_1218), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1218 ( .A(n_1112), .Y(n_1218) );
XNOR2x1_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1162), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1138), .Y(n_1113) );
AND4x1_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1118), .C(n_1122), .D(n_1125), .Y(n_1114) );
OAI211xp5_ASAP7_75t_L g1144 ( .A1(n_1121), .A2(n_1145), .B(n_1146), .C(n_1147), .Y(n_1144) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
AOI31xp33_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1150), .A3(n_1158), .B(n_1161), .Y(n_1140) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1148), .Y(n_1654) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1149), .Y(n_1206) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx2_ASAP7_75t_SL g1561 ( .A(n_1154), .Y(n_1561) );
AOI31xp33_ASAP7_75t_L g1197 ( .A1(n_1161), .A2(n_1198), .A3(n_1207), .B(n_1214), .Y(n_1197) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1194), .Y(n_1167) );
AND4x1_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1175), .C(n_1179), .D(n_1182), .Y(n_1168) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
AOI21xp33_ASAP7_75t_SL g1194 ( .A1(n_1195), .A2(n_1196), .B(n_1197), .Y(n_1194) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
XNOR2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
AND4x1_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1226), .C(n_1256), .D(n_1285), .Y(n_1223) );
NOR3xp33_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1251), .C(n_1252), .Y(n_1226) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
CKINVDCx5p33_ASAP7_75t_R g1659 ( .A(n_1230), .Y(n_1659) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_1232), .A2(n_1233), .B1(n_1234), .B2(n_1237), .C(n_1238), .Y(n_1231) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1240), .Y(n_1565) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1245), .B1(n_1246), .B2(n_1248), .C(n_1249), .Y(n_1243) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_1262), .A2(n_1548), .B1(n_1549), .B2(n_1550), .Y(n_1547) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1268), .B1(n_1269), .B2(n_1271), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_1270), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_1280), .A2(n_1282), .B1(n_1283), .B2(n_1284), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
NOR2xp33_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_1292), .A2(n_1523), .B1(n_1525), .B2(n_1570), .C(n_1574), .Y(n_1291) );
AND3x1_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1481), .C(n_1511), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_1294), .A2(n_1381), .B1(n_1389), .B2(n_1432), .C(n_1459), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1366), .Y(n_1294) );
O2A1O1Ixp33_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1347), .B(n_1350), .C(n_1355), .Y(n_1295) );
AOI21xp5_ASAP7_75t_L g1493 ( .A1(n_1296), .A2(n_1494), .B(n_1496), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1324), .Y(n_1296) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1297), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1297), .B(n_1379), .Y(n_1480) );
INVx2_ASAP7_75t_L g1496 ( .A(n_1297), .Y(n_1496) );
INVx2_ASAP7_75t_SL g1297 ( .A(n_1298), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1298), .B(n_1369), .Y(n_1372) );
AND2x4_ASAP7_75t_L g1380 ( .A(n_1298), .B(n_1351), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1298), .B(n_1352), .Y(n_1394) );
HB1xp67_ASAP7_75t_L g1410 ( .A(n_1298), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1298), .B(n_1382), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g1298 ( .A(n_1299), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1299), .B(n_1351), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1299), .B(n_1352), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1314), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1308), .B1(n_1309), .B2(n_1313), .Y(n_1300) );
BUFx3_ASAP7_75t_L g1426 ( .A(n_1301), .Y(n_1426) );
BUFx6f_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1304), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_1303), .B(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1303), .Y(n_1331) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1304), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1307), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1307), .Y(n_1318) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_1309), .Y(n_1428) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1312), .Y(n_1333) );
OAI22xp5_ASAP7_75t_L g1314 ( .A1(n_1315), .A2(n_1320), .B1(n_1321), .B2(n_1323), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
BUFx3_ASAP7_75t_L g1424 ( .A(n_1316), .Y(n_1424) );
AND2x4_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1319), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1317), .B(n_1319), .Y(n_1335) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
AND2x4_ASAP7_75t_L g1322 ( .A(n_1318), .B(n_1319), .Y(n_1322) );
INVx2_ASAP7_75t_L g1388 ( .A(n_1321), .Y(n_1388) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1325), .B(n_1339), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1325), .B(n_1379), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1325), .B(n_1344), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1325), .B(n_1358), .Y(n_1477) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
NOR2xp33_ASAP7_75t_L g1445 ( .A(n_1326), .B(n_1379), .Y(n_1445) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1326), .B(n_1483), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1522 ( .A(n_1326), .B(n_1422), .Y(n_1522) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1336), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1327), .B(n_1336), .Y(n_1349) );
INVx2_ASAP7_75t_L g1363 ( .A(n_1327), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1327), .B(n_1377), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1327), .B(n_1376), .Y(n_1442) );
NOR2xp33_ASAP7_75t_L g1474 ( .A(n_1327), .B(n_1377), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1334), .Y(n_1327) );
AND2x4_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
AND2x4_ASAP7_75t_L g1332 ( .A(n_1331), .B(n_1333), .Y(n_1332) );
BUFx2_ASAP7_75t_L g1386 ( .A(n_1332), .Y(n_1386) );
HB1xp67_ASAP7_75t_L g1669 ( .A(n_1333), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1336), .B(n_1363), .Y(n_1362) );
INVx2_ASAP7_75t_SL g1376 ( .A(n_1336), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1336), .B(n_1344), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1336), .B(n_1377), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1339), .B(n_1349), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1339), .B(n_1362), .Y(n_1393) );
INVxp67_ASAP7_75t_SL g1443 ( .A(n_1339), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1343), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1340), .B(n_1349), .Y(n_1359) );
INVx2_ASAP7_75t_L g1369 ( .A(n_1340), .Y(n_1369) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1340), .Y(n_1379) );
BUFx2_ASAP7_75t_L g1398 ( .A(n_1340), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1422 ( .A(n_1340), .B(n_1377), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1340), .B(n_1404), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1343), .B(n_1362), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1343), .B(n_1349), .Y(n_1406) );
NOR2x1_ASAP7_75t_L g1453 ( .A(n_1343), .B(n_1376), .Y(n_1453) );
NOR2xp33_ASAP7_75t_L g1506 ( .A(n_1343), .B(n_1363), .Y(n_1506) );
BUFx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVxp67_ASAP7_75t_L g1358 ( .A(n_1344), .Y(n_1358) );
BUFx3_ASAP7_75t_L g1377 ( .A(n_1344), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1346), .Y(n_1344) );
AOI21xp5_ASAP7_75t_L g1516 ( .A1(n_1347), .A2(n_1496), .B(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1349), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1349), .B(n_1421), .Y(n_1420) );
OAI221xp5_ASAP7_75t_L g1439 ( .A1(n_1349), .A2(n_1440), .B1(n_1441), .B2(n_1443), .C(n_1444), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1349), .B(n_1379), .Y(n_1502) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1350), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1514 ( .A(n_1350), .B(n_1398), .Y(n_1514) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1351), .B(n_1384), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1465 ( .A(n_1351), .B(n_1466), .Y(n_1465) );
A2O1A1Ixp33_ASAP7_75t_SL g1511 ( .A1(n_1351), .A2(n_1429), .B(n_1512), .C(n_1513), .Y(n_1511) );
INVx3_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1352), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1438 ( .A(n_1352), .B(n_1384), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1352), .B(n_1383), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1354), .Y(n_1352) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1360), .B(n_1364), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
AOI22xp5_ASAP7_75t_L g1498 ( .A1(n_1357), .A2(n_1413), .B1(n_1499), .B2(n_1501), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1359), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1358), .B(n_1362), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1358), .B(n_1442), .Y(n_1492) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1362), .B(n_1379), .Y(n_1488) );
A2O1A1Ixp33_ASAP7_75t_L g1447 ( .A1(n_1363), .A2(n_1448), .B(n_1451), .C(n_1454), .Y(n_1447) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
O2A1O1Ixp33_ASAP7_75t_L g1419 ( .A1(n_1365), .A2(n_1420), .B(n_1423), .C(n_1429), .Y(n_1419) );
OAI21xp5_ASAP7_75t_L g1460 ( .A1(n_1365), .A2(n_1368), .B(n_1461), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1365), .B(n_1369), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1365), .B(n_1519), .Y(n_1518) );
AOI211xp5_ASAP7_75t_SL g1366 ( .A1(n_1367), .A2(n_1368), .B(n_1371), .C(n_1373), .Y(n_1366) );
A2O1A1Ixp33_ASAP7_75t_SL g1490 ( .A1(n_1367), .A2(n_1489), .B(n_1491), .C(n_1493), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1370), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1369), .B(n_1506), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1370), .B(n_1372), .Y(n_1371) );
NOR2xp33_ASAP7_75t_L g1515 ( .A(n_1370), .B(n_1408), .Y(n_1515) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1372), .Y(n_1440) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1378), .Y(n_1373) );
OAI221xp5_ASAP7_75t_L g1389 ( .A1(n_1374), .A2(n_1390), .B1(n_1411), .B2(n_1412), .C(n_1414), .Y(n_1389) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1377), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1377), .B(n_1392), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1377), .B(n_1502), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1380), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1379), .B(n_1404), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1379), .B(n_1408), .Y(n_1407) );
OAI21xp33_ASAP7_75t_L g1475 ( .A1(n_1379), .A2(n_1402), .B(n_1476), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1380), .B(n_1382), .Y(n_1413) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_1380), .A2(n_1415), .B1(n_1472), .B2(n_1475), .C(n_1478), .Y(n_1471) );
AOI21xp5_ASAP7_75t_L g1487 ( .A1(n_1380), .A2(n_1488), .B(n_1489), .Y(n_1487) );
INVx2_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1382), .B(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1383), .Y(n_1431) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1384), .Y(n_1411) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1384), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1387), .Y(n_1384) );
AOI22xp5_ASAP7_75t_L g1432 ( .A1(n_1390), .A2(n_1433), .B1(n_1436), .B2(n_1447), .Y(n_1432) );
AND3x1_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1395), .C(n_1405), .Y(n_1390) );
OAI21xp5_ASAP7_75t_L g1391 ( .A1(n_1392), .A2(n_1393), .B(n_1394), .Y(n_1391) );
AOI221xp5_ASAP7_75t_L g1414 ( .A1(n_1393), .A2(n_1415), .B1(n_1417), .B2(n_1418), .C(n_1419), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1394), .B(n_1450), .Y(n_1449) );
A2O1A1Ixp33_ASAP7_75t_L g1503 ( .A1(n_1394), .A2(n_1423), .B(n_1504), .C(n_1507), .Y(n_1503) );
AOI22xp5_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1399), .B1(n_1400), .B2(n_1403), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
AOI21xp5_ASAP7_75t_L g1507 ( .A1(n_1397), .A2(n_1401), .B(n_1476), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1399), .Y(n_1397) );
INVx2_ASAP7_75t_L g1450 ( .A(n_1398), .Y(n_1450) );
NAND2xp5_ASAP7_75t_SL g1473 ( .A(n_1398), .B(n_1474), .Y(n_1473) );
CKINVDCx5p33_ASAP7_75t_R g1470 ( .A(n_1399), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1402), .Y(n_1400) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1403), .Y(n_1486) );
OAI21xp33_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1407), .B(n_1409), .Y(n_1405) );
AOI221xp5_ASAP7_75t_L g1463 ( .A1(n_1406), .A2(n_1407), .B1(n_1418), .B2(n_1464), .C(n_1467), .Y(n_1463) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1407), .Y(n_1485) );
INVxp67_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_1410), .B(n_1522), .Y(n_1521) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1411), .B(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1413), .B(n_1417), .Y(n_1510) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1418), .Y(n_1500) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1423), .B(n_1430), .Y(n_1429) );
INVx3_ASAP7_75t_L g1435 ( .A(n_1423), .Y(n_1435) );
AOI31xp33_ASAP7_75t_L g1459 ( .A1(n_1423), .A2(n_1460), .A3(n_1463), .B(n_1471), .Y(n_1459) );
INVx3_ASAP7_75t_L g1489 ( .A(n_1423), .Y(n_1489) );
BUFx2_ASAP7_75t_SL g1524 ( .A(n_1428), .Y(n_1524) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
AOI211xp5_ASAP7_75t_L g1436 ( .A1(n_1431), .A2(n_1437), .B(n_1439), .C(n_1446), .Y(n_1436) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1431), .Y(n_1469) );
NAND3xp33_ASAP7_75t_SL g1479 ( .A(n_1431), .B(n_1442), .C(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1467 ( .A(n_1441), .B(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
AOI21xp33_ASAP7_75t_L g1508 ( .A1(n_1446), .A2(n_1509), .B(n_1510), .Y(n_1508) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1450), .B(n_1453), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1491 ( .A(n_1450), .B(n_1492), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1450), .B(n_1474), .Y(n_1495) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1457), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1458), .B(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1470), .Y(n_1468) );
A2O1A1Ixp33_ASAP7_75t_L g1484 ( .A1(n_1470), .A2(n_1485), .B(n_1486), .C(n_1487), .Y(n_1484) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
O2A1O1Ixp33_ASAP7_75t_L g1481 ( .A1(n_1482), .A2(n_1484), .B(n_1490), .C(n_1497), .Y(n_1481) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1491), .Y(n_1512) );
INVx2_ASAP7_75t_L g1519 ( .A(n_1492), .Y(n_1519) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
NAND3xp33_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1503), .C(n_1508), .Y(n_1497) );
INVxp67_ASAP7_75t_SL g1504 ( .A(n_1505), .Y(n_1504) );
OAI211xp5_ASAP7_75t_L g1513 ( .A1(n_1514), .A2(n_1515), .B(n_1516), .C(n_1520), .Y(n_1513) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
HB1xp67_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1554), .Y(n_1526) );
NOR3xp33_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1535), .C(n_1536), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1532), .Y(n_1528) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
CKINVDCx5p33_ASAP7_75t_R g1570 ( .A(n_1571), .Y(n_1570) );
BUFx2_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
OAI21xp5_ASAP7_75t_L g1668 ( .A1(n_1573), .A2(n_1669), .B(n_1670), .Y(n_1668) );
BUFx3_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
BUFx2_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
HB1xp67_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1581), .Y(n_1666) );
AOI221xp5_ASAP7_75t_L g1581 ( .A1(n_1582), .A2(n_1609), .B1(n_1611), .B2(n_1637), .C(n_1639), .Y(n_1581) );
NAND4xp25_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1591), .C(n_1600), .D(n_1606), .Y(n_1582) );
AOI22xp33_ASAP7_75t_L g1583 ( .A1(n_1584), .A2(n_1585), .B1(n_1587), .B2(n_1588), .Y(n_1583) );
AND2x4_ASAP7_75t_L g1588 ( .A(n_1586), .B(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
AOI222xp33_ASAP7_75t_L g1591 ( .A1(n_1592), .A2(n_1593), .B1(n_1594), .B2(n_1595), .C1(n_1596), .C2(n_1597), .Y(n_1591) );
INVxp67_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1599), .Y(n_1608) );
AOI22xp33_ASAP7_75t_L g1600 ( .A1(n_1601), .A2(n_1602), .B1(n_1603), .B2(n_1604), .Y(n_1600) );
AOI22xp33_ASAP7_75t_L g1622 ( .A1(n_1603), .A2(n_1623), .B1(n_1626), .B2(n_1627), .Y(n_1622) );
INVx4_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
CKINVDCx11_ASAP7_75t_R g1606 ( .A(n_1607), .Y(n_1606) );
CKINVDCx16_ASAP7_75t_R g1609 ( .A(n_1610), .Y(n_1609) );
NAND4xp25_ASAP7_75t_SL g1611 ( .A(n_1612), .B(n_1622), .C(n_1628), .D(n_1634), .Y(n_1611) );
AOI22xp33_ASAP7_75t_L g1612 ( .A1(n_1613), .A2(n_1614), .B1(n_1618), .B2(n_1619), .Y(n_1612) );
AND2x4_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1617), .Y(n_1614) );
INVx1_ASAP7_75t_SL g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1620), .Y(n_1636) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
AND2x2_ASAP7_75t_SL g1630 ( .A(n_1624), .B(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
CKINVDCx8_ASAP7_75t_R g1634 ( .A(n_1635), .Y(n_1634) );
NAND4xp25_ASAP7_75t_SL g1639 ( .A(n_1640), .B(n_1646), .C(n_1651), .D(n_1660), .Y(n_1639) );
NAND3xp33_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1656), .C(n_1659), .Y(n_1651) );
INVx2_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
NAND3xp33_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1663), .C(n_1664), .Y(n_1660) );
HB1xp67_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
endmodule