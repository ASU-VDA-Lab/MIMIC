module fake_jpeg_17115_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_56),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_47),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_62),
.B(n_68),
.C(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_42),
.B1(n_45),
.B2(n_44),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_79),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_1),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_18),
.B1(n_35),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_82),
.B1(n_3),
.B2(n_4),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_3),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_0),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_4),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_13),
.B(n_14),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_9),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_78),
.B1(n_75),
.B2(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_20),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_15),
.C(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_21),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_104),
.B(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_105),
.B(n_103),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_108),
.B(n_90),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_108),
.B(n_101),
.C(n_25),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_22),
.C(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_26),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_30),
.Y(n_116)
);


endmodule