module real_jpeg_20183_n_11 (n_5, n_4, n_8, n_0, n_245, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_245;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_0),
.A2(n_2),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_6),
.B1(n_21),
.B2(n_40),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_0),
.A2(n_5),
.B1(n_40),
.B2(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_0),
.A2(n_4),
.B1(n_26),
.B2(n_40),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_6),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_4),
.B1(n_20),
.B2(n_26),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_5),
.B1(n_20),
.B2(n_52),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_10),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_36),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_32),
.B(n_36),
.C(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_4),
.A2(n_7),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_4),
.A2(n_9),
.B1(n_26),
.B2(n_53),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_10),
.B1(n_26),
.B2(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_32),
.B(n_53),
.C(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_9),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_5),
.B(n_91),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_10),
.B1(n_32),
.B2(n_52),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_5),
.A2(n_9),
.B(n_10),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_7),
.B1(n_21),
.B2(n_25),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_8),
.B1(n_21),
.B2(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_10),
.B1(n_21),
.B2(n_32),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_10),
.B(n_104),
.Y(n_103)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_7),
.A2(n_10),
.B(n_21),
.C(n_149),
.Y(n_148)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_10),
.B(n_41),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_24),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_71),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_70),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_58),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_15),
.B(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_29),
.B2(n_30),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_24),
.B1(n_27),
.B2(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_23),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_24),
.A2(n_27),
.B1(n_47),
.B2(n_68),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_25),
.A2(n_26),
.B(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_32),
.B(n_51),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_32),
.B(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.C(n_48),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_83),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_61),
.B1(n_83),
.B2(n_84),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_44),
.A2(n_61),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_44),
.A2(n_83),
.B(n_100),
.C(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_44),
.A2(n_61),
.B1(n_200),
.B2(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_44),
.A2(n_61),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_44),
.A2(n_201),
.B(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_44),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_48),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_48),
.A2(n_65),
.B1(n_67),
.B2(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_56),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_51),
.A2(n_54),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OA22x2_ASAP7_75t_SL g216 ( 
.A1(n_51),
.A2(n_54),
.B1(n_56),
.B2(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_52),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_66),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_65),
.C(n_67),
.Y(n_66)
);

AOI211xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_80),
.B(n_82),
.C(n_86),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_61),
.B(n_84),
.Y(n_208)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_66),
.B(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_225),
.A3(n_236),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_210),
.B(n_224),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_192),
.B(n_209),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_119),
.B(n_174),
.C(n_191),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_108),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_76),
.B(n_108),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_97),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_88),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_78),
.B(n_88),
.C(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_85),
.B1(n_89),
.B2(n_96),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_85),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_85),
.B1(n_126),
.B2(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_105),
.C(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_80),
.A2(n_85),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_80),
.B(n_157),
.C(n_163),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_80),
.A2(n_85),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_80),
.B(n_89),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_80),
.B(n_181),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_82),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_83),
.A2(n_85),
.B(n_151),
.C(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_83),
.A2(n_84),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_83),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_83),
.B(n_216),
.Y(n_217)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_105),
.C(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_86),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_107),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_98),
.A2(n_99),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_98),
.A2(n_99),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_115),
.B1(n_129),
.B2(n_132),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_115),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_160)
);

NAND2x1_ASAP7_75t_SL g164 ( 
.A(n_105),
.B(n_148),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_116),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_110),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_147),
.B2(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_116),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_173),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_166),
.B(n_172),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_153),
.B(n_165),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_144),
.B(n_152),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_133),
.B(n_143),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_128),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_129),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_146),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_148),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_156),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_176),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_188),
.B2(n_190),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_187),
.C(n_190),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_189),
.B(n_208),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_188),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_197),
.B(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_194),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_211),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.CI(n_207),
.CON(n_195),
.SN(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_197),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_206),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_203),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_222),
.B2(n_223),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_219),
.C(n_223),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_227),
.B1(n_231),
.B2(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.C(n_232),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);


endmodule