module fake_jpeg_27809_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_0),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_79),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_66),
.B1(n_63),
.B2(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_91),
.B1(n_48),
.B2(n_71),
.Y(n_104)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_51),
.B1(n_64),
.B2(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_59),
.B1(n_61),
.B2(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_64),
.B1(n_51),
.B2(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_92),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_62),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_57),
.CI(n_61),
.CON(n_97),
.SN(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_87),
.B(n_86),
.Y(n_114)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_104),
.B1(n_109),
.B2(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_86),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_106),
.B(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_97),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_120),
.B(n_123),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_100),
.B1(n_99),
.B2(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_1),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_119),
.B1(n_115),
.B2(n_68),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_115),
.B1(n_47),
.B2(n_56),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_20),
.B1(n_43),
.B2(n_42),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_4),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_14),
.B(n_40),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_15),
.B(n_31),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_13),
.B1(n_37),
.B2(n_33),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_10),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_152),
.C(n_137),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_2),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_147),
.C(n_151),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_145),
.B(n_148),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_134),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_153),
.C(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_150),
.C(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_45),
.B1(n_30),
.B2(n_29),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_27),
.B(n_26),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_24),
.B(n_5),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_8),
.Y(n_165)
);


endmodule