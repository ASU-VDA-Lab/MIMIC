module fake_jpeg_27615_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_39),
.Y(n_41)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_15),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_40),
.A2(n_50),
.B1(n_33),
.B2(n_36),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_52),
.B1(n_33),
.B2(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_46),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_15),
.B1(n_31),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_15),
.B1(n_31),
.B2(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_54),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_33),
.B1(n_36),
.B2(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_62),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_53),
.B1(n_32),
.B2(n_31),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_70),
.B1(n_42),
.B2(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_35),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_76),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_32),
.B1(n_0),
.B2(n_2),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_16),
.C(n_29),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_18),
.B(n_22),
.C(n_17),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_22),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_32),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_101),
.B1(n_0),
.B2(n_1),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_50),
.B(n_40),
.C(n_52),
.Y(n_87)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_56),
.B(n_74),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_50),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_45),
.B1(n_32),
.B2(n_16),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_96),
.B1(n_74),
.B2(n_56),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_47),
.B1(n_45),
.B2(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_25),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_61),
.B1(n_78),
.B2(n_77),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_57),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_105),
.B(n_94),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_128),
.B1(n_131),
.B2(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_111),
.B(n_114),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_72),
.C(n_60),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_90),
.C(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_68),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_122),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_60),
.B(n_58),
.C(n_79),
.D(n_64),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_65),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_65),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_9),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_9),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_10),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_104),
.B(n_94),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_74),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_86),
.B(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_85),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_141),
.C(n_124),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_84),
.B(n_93),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_118),
.B1(n_110),
.B2(n_127),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_94),
.B(n_93),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_147),
.B(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_156),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_109),
.B(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_158),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_94),
.B(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_169),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_112),
.C(n_124),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_141),
.C(n_154),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_177),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_153),
.B1(n_138),
.B2(n_132),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_131),
.B1(n_128),
.B2(n_126),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_107),
.C(n_1),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_86),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_126),
.B1(n_108),
.B2(n_119),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_119),
.B1(n_91),
.B2(n_4),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_135),
.B1(n_134),
.B2(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_137),
.B(n_133),
.Y(n_189)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_8),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_177),
.B1(n_163),
.B2(n_164),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_139),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_172),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_133),
.B1(n_142),
.B2(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_197),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_199),
.C(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_146),
.B1(n_147),
.B2(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_171),
.B1(n_167),
.B2(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_144),
.C(n_158),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_206),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_8),
.B1(n_1),
.B2(n_4),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_159),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_190),
.B1(n_168),
.B2(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_189),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_212),
.C(n_186),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_181),
.C(n_161),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_187),
.C(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_214),
.B1(n_10),
.B2(n_4),
.Y(n_226)
);

AOI22x1_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_170),
.B1(n_180),
.B2(n_174),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_197),
.B1(n_191),
.B2(n_190),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_226),
.B1(n_203),
.B2(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_225),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_156),
.C(n_178),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_219),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_229),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_5),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_202),
.B1(n_200),
.B2(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_234),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_5),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_240),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_220),
.B(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_233),
.B1(n_232),
.B2(n_234),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_240),
.B(n_230),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_12),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_242),
.A2(n_229),
.B1(n_6),
.B2(n_10),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_239),
.B(n_6),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_0),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_228),
.C2(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_13),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_13),
.Y(n_256)
);


endmodule