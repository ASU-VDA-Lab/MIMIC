module fake_jpeg_15276_n_298 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_64),
.Y(n_88)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_4),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_68),
.Y(n_117)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_34),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_24),
.A2(n_9),
.B(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_13),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_29),
.B1(n_23),
.B2(n_20),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_102),
.B1(n_106),
.B2(n_99),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_77),
.B1(n_97),
.B2(n_115),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_39),
.B1(n_24),
.B2(n_38),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_39),
.B1(n_25),
.B2(n_15),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_79),
.A2(n_82),
.B1(n_101),
.B2(n_85),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_25),
.B1(n_15),
.B2(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_83),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_108),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_43),
.A2(n_35),
.B1(n_29),
.B2(n_27),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_46),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_10),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_18),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_60),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_65),
.B1(n_30),
.B2(n_2),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_119),
.A2(n_145),
.B1(n_137),
.B2(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_0),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_10),
.B(n_0),
.C(n_1),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_127),
.Y(n_168)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_78),
.Y(n_130)
);

BUFx2_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_84),
.B1(n_100),
.B2(n_107),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_73),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_110),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_84),
.A2(n_100),
.B1(n_81),
.B2(n_115),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_73),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_75),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_98),
.B(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_155),
.Y(n_173)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_79),
.B(n_75),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_119),
.Y(n_165)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_86),
.B(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_37),
.B1(n_33),
.B2(n_16),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_159),
.B(n_120),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_92),
.A2(n_37),
.B1(n_33),
.B2(n_16),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_92),
.B(n_104),
.C(n_125),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_167),
.B(n_156),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_157),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_122),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_139),
.C(n_147),
.Y(n_208)
);

NOR2x1_ASAP7_75t_R g167 ( 
.A(n_121),
.B(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_175),
.B1(n_151),
.B2(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_143),
.B1(n_127),
.B2(n_124),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_177),
.B(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_185),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_168),
.B(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_148),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_131),
.B(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_136),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g190 ( 
.A(n_160),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_195),
.B(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_217),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_146),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_198),
.B(n_199),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_160),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_200),
.B(n_209),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_158),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_212),
.C(n_216),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_128),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_168),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_215),
.A2(n_165),
.B(n_187),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_154),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_181),
.B(n_161),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_161),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_233),
.B(n_217),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_227),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_204),
.A3(n_217),
.B1(n_203),
.B2(n_212),
.C1(n_213),
.C2(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_234),
.C(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_170),
.B1(n_201),
.B2(n_187),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_243),
.B1(n_192),
.B2(n_179),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_175),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_173),
.A3(n_194),
.B1(n_184),
.B2(n_186),
.C1(n_193),
.C2(n_177),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_178),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_173),
.C(n_172),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_196),
.A2(n_193),
.B1(n_186),
.B2(n_179),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_203),
.B(n_216),
.C(n_221),
.D(n_214),
.Y(n_244)
);

OA21x2_ASAP7_75t_SL g267 ( 
.A1(n_244),
.A2(n_245),
.B(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_198),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_260),
.Y(n_266)
);

AO221x1_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_220),
.B1(n_211),
.B2(n_172),
.C(n_207),
.Y(n_254)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_254),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_205),
.C(n_191),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_256),
.C(n_253),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_209),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_257),
.A2(n_258),
.B1(n_228),
.B2(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_233),
.B1(n_232),
.B2(n_234),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_240),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_192),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_268),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_224),
.B1(n_225),
.B2(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_260),
.B1(n_257),
.B2(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_247),
.B(n_244),
.Y(n_274)
);

AOI211xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_279),
.B(n_268),
.C(n_263),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_255),
.B(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_223),
.B(n_252),
.Y(n_279)
);

NOR2x1_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_279),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_282),
.A2(n_283),
.B1(n_266),
.B2(n_265),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_272),
.B1(n_266),
.B2(n_236),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_243),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_286),
.A2(n_273),
.B(n_264),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_290),
.B(n_282),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_284),
.A2(n_225),
.B(n_235),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_291),
.B(n_283),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_293),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_295),
.B(n_292),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_296),
.Y(n_298)
);


endmodule