module fake_netlist_6_199_n_1707 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1707);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1707;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_23),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_54),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_104),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_46),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_66),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_68),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_71),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_95),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_72),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_42),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

BUFx8_ASAP7_75t_SL g170 ( 
.A(n_61),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_59),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_82),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_1),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_87),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_74),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_42),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_38),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_108),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_115),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_29),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_10),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_62),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_23),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_15),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_75),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_49),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_84),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_131),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_51),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_101),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_30),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_73),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_130),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_144),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_37),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_27),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_53),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_110),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_96),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_43),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_122),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_90),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_32),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_83),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_5),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_28),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_140),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_142),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_25),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_147),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_18),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_148),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_0),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_4),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_126),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_97),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_127),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_100),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_77),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_34),
.Y(n_251)
);

BUFx8_ASAP7_75t_SL g252 ( 
.A(n_91),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_3),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_120),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_43),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_47),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_123),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_47),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_36),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_17),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_134),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_44),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_117),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_113),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_58),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_26),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_76),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_57),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_24),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_18),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_48),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_69),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_41),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_124),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_141),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_99),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_33),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_49),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_50),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_153),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_60),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_28),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_93),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_20),
.Y(n_297)
);

BUFx2_ASAP7_75t_SL g298 ( 
.A(n_70),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_13),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_40),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_136),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_2),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_94),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_182),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_182),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_185),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_170),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_210),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_196),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_193),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_186),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_252),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_196),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_189),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_154),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_227),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_227),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_216),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_194),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_232),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_232),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_168),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_201),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_202),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_225),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_242),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_231),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_208),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_218),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_215),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_234),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_221),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_245),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_228),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_216),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_238),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_240),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_264),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_230),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_269),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_236),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_278),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_250),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_237),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_249),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_233),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_233),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_155),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_158),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_239),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_220),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_247),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_165),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_171),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_175),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_255),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_180),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_205),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_373),
.B(n_205),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_200),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_308),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_209),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_335),
.B(n_209),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_327),
.B(n_295),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_332),
.A2(n_281),
.B1(n_303),
.B2(n_173),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_313),
.B(n_220),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_307),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_322),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_310),
.B(n_160),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_348),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_181),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_156),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_312),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_187),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_190),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_156),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_318),
.B(n_177),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_195),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_346),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_197),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_367),
.B(n_220),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_323),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_371),
.A2(n_324),
.B(n_323),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_336),
.B(n_159),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_353),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_329),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_326),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_374),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_334),
.Y(n_446)
);

BUFx8_ASAP7_75t_SL g447 ( 
.A(n_378),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_375),
.A2(n_314),
.B1(n_298),
.B2(n_340),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_375),
.B(n_338),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_374),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_420),
.B(n_342),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_419),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_395),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_388),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_410),
.B(n_330),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_405),
.B(n_345),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_381),
.B(n_350),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_374),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_414),
.A2(n_337),
.B1(n_325),
.B2(n_200),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_387),
.B(n_352),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

NOR2x1p5_ASAP7_75t_L g486 ( 
.A(n_399),
.B(n_309),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_384),
.B(n_198),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_381),
.B(n_359),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

NOR2x1p5_ASAP7_75t_L g490 ( 
.A(n_404),
.B(n_315),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_381),
.B(n_366),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_374),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_381),
.B(n_368),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_379),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_379),
.B(n_200),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_379),
.B(n_372),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_376),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g504 ( 
.A(n_387),
.B(n_154),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_L g510 ( 
.A1(n_385),
.A2(n_263),
.B1(n_207),
.B2(n_266),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_414),
.A2(n_213),
.B1(n_200),
.B2(n_355),
.Y(n_512)
);

INVx4_ASAP7_75t_SL g513 ( 
.A(n_376),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_414),
.A2(n_200),
.B1(n_213),
.B2(n_282),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_402),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_381),
.B(n_354),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_402),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_379),
.B(n_259),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_402),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_410),
.B(n_358),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_379),
.B(n_288),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_403),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_384),
.B(n_265),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_427),
.B(n_432),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_406),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_427),
.B(n_199),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_412),
.B(n_361),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_421),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_410),
.B(n_270),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_421),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

AND3x2_ASAP7_75t_L g547 ( 
.A(n_396),
.B(n_290),
.C(n_294),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_415),
.B(n_274),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_415),
.B(n_358),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_409),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_396),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_378),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_415),
.A2(n_213),
.B1(n_203),
.B2(n_204),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_412),
.A2(n_417),
.B1(n_432),
.B2(n_271),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_417),
.B(n_206),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_425),
.B(n_226),
.C(n_279),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_425),
.B(n_377),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_418),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_425),
.B(n_213),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_377),
.B(n_275),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_428),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_376),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_413),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_381),
.B(n_292),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_428),
.Y(n_570)
);

BUFx4f_ASAP7_75t_L g571 ( 
.A(n_376),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_428),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_428),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_428),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_428),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_431),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_411),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_431),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_R g580 ( 
.A(n_416),
.B(n_159),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_422),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_431),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_442),
.B(n_381),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_484),
.B(n_381),
.Y(n_585)
);

INVxp33_ASAP7_75t_L g586 ( 
.A(n_441),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_474),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_442),
.B(n_389),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_473),
.B(n_389),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_446),
.B(n_422),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_473),
.B(n_494),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_494),
.B(n_389),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_581),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_479),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_480),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_440),
.B(n_191),
.C(n_188),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_497),
.B(n_389),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_480),
.Y(n_599)
);

BUFx6f_ASAP7_75t_SL g600 ( 
.A(n_535),
.Y(n_600)
);

AO22x2_ASAP7_75t_L g601 ( 
.A1(n_452),
.A2(n_219),
.B1(n_211),
.B2(n_212),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_483),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_328),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_497),
.B(n_389),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_443),
.B(n_398),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_564),
.B(n_213),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_443),
.B(n_398),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_526),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_506),
.B(n_386),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_449),
.B(n_398),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_450),
.B(n_386),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_455),
.B(n_161),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_485),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_449),
.B(n_398),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_555),
.B(n_161),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_555),
.B(n_465),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_529),
.B(n_162),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

AND2x2_ASAP7_75t_SL g621 ( 
.A(n_564),
.B(n_571),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_530),
.A2(n_331),
.B1(n_333),
.B2(n_344),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_453),
.B(n_398),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_539),
.B(n_162),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_511),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_539),
.B(n_163),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_499),
.B(n_163),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_507),
.B(n_285),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_509),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_L g631 ( 
.A(n_504),
.B(n_217),
.C(n_257),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_448),
.B(n_164),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_530),
.A2(n_183),
.B1(n_303),
.B2(n_173),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_SL g635 ( 
.A(n_466),
.B(n_214),
.Y(n_635)
);

AOI221xp5_ASAP7_75t_L g636 ( 
.A1(n_510),
.A2(n_183),
.B1(n_157),
.B2(n_281),
.C(n_283),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_521),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_447),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_454),
.B(n_408),
.Y(n_639)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_530),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_507),
.Y(n_641)
);

AO221x1_ASAP7_75t_L g642 ( 
.A1(n_578),
.A2(n_223),
.B1(n_241),
.B2(n_248),
.C(n_268),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_530),
.B(n_164),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_511),
.B(n_429),
.Y(n_645)
);

BUFx5_ASAP7_75t_L g646 ( 
.A(n_457),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_530),
.A2(n_360),
.B1(n_166),
.B2(n_167),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_538),
.B(n_285),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_558),
.B(n_167),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_522),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_528),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_457),
.A2(n_235),
.B(n_437),
.C(n_433),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_528),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_456),
.B(n_172),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_561),
.B(n_285),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_552),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_558),
.B(n_172),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_540),
.B(n_383),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_526),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_523),
.B(n_174),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_527),
.B(n_174),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_383),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_532),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_460),
.B(n_383),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_556),
.B(n_176),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_538),
.A2(n_176),
.B1(n_305),
.B2(n_178),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_460),
.B(n_463),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_463),
.A2(n_437),
.B(n_434),
.C(n_433),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_542),
.B(n_178),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_467),
.B(n_431),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_467),
.B(n_431),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_469),
.B(n_431),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_561),
.B(n_469),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_548),
.A2(n_380),
.B(n_436),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_566),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_557),
.A2(n_361),
.B1(n_434),
.B2(n_380),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_550),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_550),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_535),
.A2(n_157),
.B1(n_283),
.B2(n_286),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_554),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_554),
.B(n_431),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_560),
.Y(n_684)
);

INVx8_ASAP7_75t_L g685 ( 
.A(n_556),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_557),
.B(n_179),
.C(n_184),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_560),
.Y(n_687)
);

CKINVDCx16_ASAP7_75t_R g688 ( 
.A(n_551),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_565),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_556),
.B(n_179),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_468),
.B(n_488),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_565),
.B(n_431),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_567),
.B(n_569),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_464),
.B(n_390),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_567),
.B(n_435),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_556),
.B(n_184),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_556),
.B(n_284),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_464),
.B(n_390),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_549),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_538),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_487),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_SL g702 ( 
.A(n_466),
.B(n_284),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_569),
.B(n_435),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_572),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_487),
.A2(n_376),
.B1(n_285),
.B2(n_287),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_487),
.A2(n_305),
.B1(n_293),
.B2(n_302),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_572),
.B(n_562),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_487),
.B(n_293),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_439),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_487),
.B(n_435),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_535),
.B(n_302),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_553),
.B(n_435),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_514),
.B(n_435),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_439),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_512),
.B(n_435),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_551),
.B(n_390),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_476),
.B(n_292),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_535),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_535),
.B(n_439),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_491),
.A2(n_376),
.B1(n_285),
.B2(n_292),
.Y(n_720)
);

OAI22x1_ASAP7_75t_SL g721 ( 
.A1(n_580),
.A2(n_300),
.B1(n_299),
.B2(n_297),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_444),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_486),
.B(n_392),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_517),
.B(n_192),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_564),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_439),
.B(n_435),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_477),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_477),
.B(n_438),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_492),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_568),
.B(n_495),
.C(n_243),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_477),
.B(n_438),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_498),
.A2(n_376),
.B1(n_285),
.B2(n_287),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_571),
.A2(n_286),
.B1(n_289),
.B2(n_297),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_561),
.B(n_285),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_478),
.B(n_438),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_486),
.B(n_392),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_498),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_704),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_611),
.B(n_547),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_625),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_662),
.B(n_608),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_704),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_660),
.B(n_500),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_700),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_625),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_611),
.A2(n_498),
.B1(n_561),
.B2(n_299),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_716),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_694),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_694),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_707),
.B(n_478),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_698),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_619),
.B(n_478),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_669),
.A2(n_500),
.B(n_481),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_594),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_656),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_699),
.B(n_500),
.Y(n_757)
);

BUFx12f_ASAP7_75t_L g758 ( 
.A(n_620),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_SL g759 ( 
.A(n_633),
.B(n_300),
.C(n_289),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_700),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_698),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_587),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_618),
.A2(n_490),
.B1(n_498),
.B2(n_561),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_595),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_700),
.B(n_500),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_609),
.B(n_229),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_725),
.B(n_466),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_619),
.A2(n_490),
.B1(n_498),
.B2(n_561),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_614),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_646),
.B(n_482),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_590),
.B(n_244),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_723),
.B(n_513),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_SL g773 ( 
.A(n_612),
.B(n_246),
.C(n_251),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_591),
.A2(n_489),
.B(n_445),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_700),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_725),
.B(n_466),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_601),
.A2(n_705),
.B1(n_633),
.B2(n_606),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_630),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_725),
.B(n_466),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_634),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_646),
.B(n_482),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_653),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_646),
.B(n_482),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_646),
.B(n_482),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_659),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_620),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_665),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_645),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_592),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_646),
.B(n_496),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_646),
.B(n_496),
.Y(n_791)
);

AOI22x1_ASAP7_75t_L g792 ( 
.A1(n_729),
.A2(n_445),
.B1(n_458),
.B2(n_489),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_592),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_641),
.A2(n_459),
.B1(n_481),
.B2(n_475),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_672),
.A2(n_458),
.B(n_459),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_603),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_584),
.B(n_496),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_641),
.A2(n_472),
.B1(n_475),
.B2(n_577),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_586),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_640),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_SL g801 ( 
.A1(n_600),
.A2(n_276),
.B1(n_253),
.B2(n_254),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_644),
.A2(n_498),
.B1(n_561),
.B2(n_472),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_612),
.B(n_466),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_621),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_679),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_601),
.A2(n_498),
.B1(n_376),
.B2(n_256),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_688),
.B(n_258),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_687),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_689),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_736),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_644),
.B(n_513),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_601),
.A2(n_376),
.B1(n_260),
.B2(n_261),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_640),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_673),
.A2(n_519),
.B(n_493),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_711),
.B(n_513),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_621),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_711),
.B(n_513),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_624),
.B(n_262),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_640),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_596),
.B(n_513),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_705),
.A2(n_273),
.B1(n_280),
.B2(n_272),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_599),
.B(n_501),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_626),
.B(n_392),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_602),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_661),
.A2(n_543),
.B1(n_519),
.B2(n_577),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_677),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_649),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_701),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_718),
.B(n_444),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_613),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_617),
.B(n_501),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_628),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_657),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_637),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_643),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_661),
.A2(n_543),
.B1(n_516),
.B2(n_525),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_622),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_650),
.Y(n_838)
);

OR2x2_ASAP7_75t_SL g839 ( 
.A(n_597),
.B(n_401),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_701),
.Y(n_840)
);

AND2x4_ASAP7_75t_SL g841 ( 
.A(n_730),
.B(n_518),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_651),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_680),
.B(n_682),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_684),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_667),
.A2(n_518),
.B(n_534),
.C(n_536),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_R g846 ( 
.A(n_701),
.B(n_52),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_693),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_685),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_733),
.B(n_501),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_471),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_606),
.B(n_444),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_678),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_674),
.A2(n_563),
.B(n_536),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_708),
.B(n_401),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_690),
.A2(n_534),
.B1(n_537),
.B2(n_545),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_709),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_714),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_678),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_722),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_654),
.Y(n_860)
);

NAND2x2_ASAP7_75t_L g861 ( 
.A(n_721),
.B(n_636),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_631),
.B(n_537),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_631),
.B(n_546),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_600),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_727),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_605),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_690),
.A2(n_573),
.B(n_546),
.C(n_563),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_607),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_678),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_654),
.B(n_505),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_610),
.Y(n_871)
);

BUFx2_ASAP7_75t_R g872 ( 
.A(n_616),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_615),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_708),
.B(n_401),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_691),
.B(n_570),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_733),
.B(n_505),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_647),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_666),
.A2(n_570),
.B(n_573),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_658),
.B(n_515),
.Y(n_880)
);

AOI21xp33_ASAP7_75t_L g881 ( 
.A1(n_696),
.A2(n_575),
.B(n_582),
.Y(n_881)
);

CKINVDCx8_ASAP7_75t_R g882 ( 
.A(n_685),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_697),
.A2(n_730),
.B1(n_629),
.B2(n_648),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_681),
.A2(n_575),
.B1(n_579),
.B2(n_471),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_719),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_664),
.B(n_670),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_652),
.A2(n_582),
.B(n_579),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_681),
.B(n_697),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_663),
.B(n_407),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_676),
.B(n_508),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_706),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_686),
.B(n_671),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_627),
.B(n_686),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_623),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_724),
.B(n_582),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_732),
.A2(n_579),
.B1(n_471),
.B2(n_502),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_629),
.B(n_502),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_710),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_639),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_648),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_588),
.B(n_576),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_642),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_589),
.B(n_593),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_732),
.A2(n_502),
.B1(n_531),
.B2(n_533),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_683),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_692),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_598),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_888),
.A2(n_632),
.B1(n_717),
.B2(n_585),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_749),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_834),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_745),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_R g912 ( 
.A(n_756),
.B(n_675),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_860),
.B(n_668),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_795),
.A2(n_728),
.B(n_735),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_859),
.A2(n_583),
.B(n_604),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_828),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_888),
.A2(n_712),
.B(n_713),
.C(n_715),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_847),
.B(n_695),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_860),
.B(n_638),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_766),
.A2(n_703),
.B(n_720),
.C(n_737),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_907),
.B(n_726),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_826),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_766),
.B(n_737),
.Y(n_923)
);

CKINVDCx6p67_ASAP7_75t_R g924 ( 
.A(n_758),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_828),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_800),
.B(n_524),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_903),
.A2(n_731),
.B(n_734),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_753),
.A2(n_655),
.B(n_533),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_773),
.A2(n_893),
.B1(n_739),
.B2(n_892),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_750),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_907),
.B(n_533),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_795),
.A2(n_531),
.B(n_515),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_859),
.B(n_461),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_883),
.A2(n_702),
.B(n_531),
.C(n_576),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_828),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_752),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_747),
.B(n_574),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_747),
.B(n_574),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_859),
.A2(n_470),
.B(n_462),
.Y(n_939)
);

AND2x2_ASAP7_75t_SL g940 ( 
.A(n_777),
.B(n_407),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_SL g941 ( 
.A1(n_849),
.A2(n_635),
.B(n_574),
.C(n_515),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_744),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_748),
.B(n_541),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_866),
.B(n_520),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_868),
.B(n_520),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_740),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_837),
.B(n_112),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_748),
.B(n_541),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_761),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_828),
.Y(n_950)
);

INVx3_ASAP7_75t_SL g951 ( 
.A(n_864),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_744),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_877),
.A2(n_470),
.B(n_461),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_871),
.B(n_541),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_R g955 ( 
.A(n_773),
.B(n_121),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_848),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_834),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_902),
.A2(n_436),
.B(n_426),
.C(n_407),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_877),
.A2(n_470),
.B(n_461),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_755),
.B(n_541),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_771),
.A2(n_524),
.B(n_520),
.C(n_426),
.Y(n_961)
);

BUFx8_ASAP7_75t_SL g962 ( 
.A(n_786),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_838),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_755),
.B(n_740),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_835),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_877),
.A2(n_559),
.B(n_470),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_L g967 ( 
.A(n_771),
.B(n_426),
.C(n_436),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_848),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_838),
.Y(n_969)
);

AOI21xp33_ASAP7_75t_L g970 ( 
.A1(n_777),
.A2(n_524),
.B(n_520),
.Y(n_970)
);

OAI21x1_ASAP7_75t_SL g971 ( 
.A1(n_858),
.A2(n_150),
.B(n_146),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_877),
.B(n_559),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_739),
.A2(n_833),
.B(n_827),
.C(n_849),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_873),
.B(n_559),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_869),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_848),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_744),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_810),
.B(n_559),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_SL g979 ( 
.A1(n_876),
.A2(n_470),
.B(n_462),
.C(n_461),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_814),
.A2(n_462),
.B(n_461),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_824),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_830),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_840),
.B(n_86),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_832),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_6),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_770),
.A2(n_783),
.B(n_781),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_905),
.B(n_462),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_741),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_746),
.A2(n_462),
.B1(n_451),
.B2(n_438),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_906),
.B(n_451),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_754),
.A2(n_451),
.B(n_438),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_894),
.B(n_451),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_SL g993 ( 
.A1(n_878),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_788),
.B(n_796),
.Y(n_994)
);

OAI21xp33_ASAP7_75t_SL g995 ( 
.A1(n_851),
.A2(n_12),
.B(n_13),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_842),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_886),
.A2(n_451),
.B(n_438),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_784),
.A2(n_438),
.B(n_133),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_876),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_746),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_799),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_846),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_SL g1003 ( 
.A1(n_891),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_788),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_852),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_843),
.B(n_89),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_846),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_840),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_843),
.A2(n_80),
.B1(n_78),
.B2(n_65),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_885),
.B(n_56),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_899),
.B(n_854),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_759),
.B(n_21),
.C(n_22),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_807),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_818),
.B(n_25),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_840),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_823),
.B(n_26),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_738),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_790),
.A2(n_48),
.B(n_30),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_759),
.A2(n_29),
.B(n_31),
.C(n_34),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_839),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_742),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_844),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_885),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_874),
.B(n_31),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_882),
.B(n_35),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_744),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_769),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_848),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_856),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_791),
.A2(n_46),
.B(n_39),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_751),
.A2(n_36),
.B(n_40),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_898),
.B(n_45),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_819),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_813),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_813),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_SL g1036 ( 
.A(n_861),
.B(n_45),
.C(n_778),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_787),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_808),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_813),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_845),
.A2(n_867),
.B(n_809),
.C(n_889),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_885),
.B(n_804),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_760),
.B(n_775),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_857),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_884),
.A2(n_816),
.B1(n_804),
.B2(n_812),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_900),
.B(n_804),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_865),
.Y(n_1046)
);

AOI33xp33_ASAP7_75t_L g1047 ( 
.A1(n_821),
.A2(n_801),
.A3(n_812),
.B1(n_806),
.B2(n_884),
.B3(n_762),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_1004),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_994),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_932),
.A2(n_774),
.B(n_887),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_1039),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1011),
.B(n_900),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1005),
.B(n_1014),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_1044),
.A2(n_798),
.A3(n_794),
.B(n_870),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_R g1055 ( 
.A(n_912),
.B(n_1002),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1011),
.B(n_804),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_980),
.A2(n_879),
.B(n_853),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_929),
.A2(n_768),
.B(n_763),
.C(n_841),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_980),
.A2(n_881),
.B(n_774),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_986),
.A2(n_803),
.B(n_793),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_946),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_1000),
.B(n_872),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_981),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_914),
.A2(n_792),
.B(n_890),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_923),
.B(n_816),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_997),
.A2(n_754),
.B(n_901),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_982),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1047),
.A2(n_862),
.B(n_863),
.C(n_780),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_1015),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_918),
.B(n_816),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1020),
.B(n_801),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_991),
.A2(n_811),
.B(n_880),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_964),
.A2(n_821),
.B(n_985),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_984),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1001),
.B(n_1007),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_918),
.B(n_816),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_991),
.A2(n_793),
.B(n_815),
.Y(n_1077)
);

AOI211x1_ASAP7_75t_L g1078 ( 
.A1(n_1000),
.A2(n_829),
.B(n_817),
.C(n_831),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_1034),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_973),
.A2(n_862),
.B(n_863),
.C(n_782),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_928),
.A2(n_797),
.B(n_822),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_1044),
.A2(n_805),
.A3(n_785),
.B(n_764),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_919),
.B(n_775),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_915),
.A2(n_917),
.B(n_1040),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1045),
.B(n_760),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_911),
.B(n_789),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_1013),
.B(n_789),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_910),
.B(n_800),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_920),
.A2(n_836),
.B(n_825),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_913),
.A2(n_776),
.B(n_779),
.C(n_765),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_922),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_934),
.A2(n_855),
.B(n_904),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1032),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_908),
.A2(n_802),
.B(n_895),
.C(n_806),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_979),
.A2(n_875),
.B(n_757),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1016),
.A2(n_895),
.B(n_875),
.C(n_897),
.Y(n_1096)
);

BUFx10_ASAP7_75t_L g1097 ( 
.A(n_983),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_957),
.B(n_850),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1024),
.A2(n_743),
.B(n_850),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_963),
.B(n_800),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1039),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1035),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_989),
.A2(n_897),
.B(n_896),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_SL g1104 ( 
.A1(n_1024),
.A2(n_772),
.B(n_820),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_1039),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_961),
.A2(n_904),
.A3(n_896),
.B(n_850),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_989),
.A2(n_800),
.A3(n_767),
.B(n_819),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_939),
.A2(n_767),
.B(n_819),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1023),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_970),
.A2(n_772),
.B(n_820),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_916),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_969),
.B(n_819),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1045),
.B(n_921),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_921),
.B(n_931),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1019),
.A2(n_995),
.B(n_958),
.C(n_988),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1008),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1031),
.A2(n_999),
.B(n_1030),
.C(n_1018),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_965),
.B(n_996),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_916),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_953),
.A2(n_959),
.B(n_966),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_916),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_931),
.B(n_940),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_925),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_925),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1022),
.B(n_937),
.Y(n_1125)
);

OA21x2_ASAP7_75t_L g1126 ( 
.A1(n_970),
.A2(n_967),
.B(n_998),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1027),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_1036),
.B(n_1003),
.C(n_1012),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_925),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_938),
.B(n_974),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_974),
.B(n_960),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_943),
.B(n_948),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_947),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_944),
.B(n_954),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_945),
.A2(n_990),
.B(n_987),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_935),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_941),
.A2(n_971),
.B(n_1041),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_933),
.A2(n_972),
.B(n_978),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_987),
.A2(n_990),
.B(n_992),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_993),
.A2(n_1037),
.B1(n_1038),
.B2(n_936),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_909),
.B(n_949),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_992),
.A2(n_1010),
.B(n_1021),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1006),
.A2(n_926),
.B(n_930),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1017),
.A2(n_1046),
.B(n_1043),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_983),
.A2(n_1009),
.B1(n_951),
.B2(n_1029),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_926),
.A2(n_1026),
.B(n_942),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_975),
.A2(n_955),
.B1(n_1025),
.B2(n_1028),
.C(n_1042),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_935),
.A2(n_968),
.B1(n_976),
.B2(n_950),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_942),
.A2(n_1026),
.B(n_977),
.C(n_950),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_977),
.A2(n_952),
.B(n_1033),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_L g1151 ( 
.A(n_924),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_935),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_950),
.B(n_956),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_956),
.A2(n_968),
.B1(n_976),
.B2(n_962),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_968),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_976),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_927),
.A2(n_877),
.B(n_859),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_927),
.A2(n_877),
.B(n_859),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_929),
.A2(n_888),
.B(n_611),
.C(n_484),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_927),
.A2(n_877),
.B(n_859),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_929),
.A2(n_888),
.B(n_611),
.C(n_484),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_994),
.B(n_716),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1000),
.B(n_888),
.Y(n_1163)
);

CKINVDCx14_ASAP7_75t_R g1164 ( 
.A(n_922),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_913),
.A2(n_888),
.B(n_618),
.C(n_484),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_932),
.A2(n_914),
.B(n_795),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_932),
.A2(n_914),
.B(n_795),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1000),
.A2(n_618),
.B(n_920),
.C(n_1006),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_916),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1015),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_981),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_927),
.A2(n_877),
.B(n_859),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_927),
.A2(n_877),
.B(n_859),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_916),
.Y(n_1174)
);

AND2x6_ASAP7_75t_L g1175 ( 
.A(n_983),
.B(n_804),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_SL g1176 ( 
.A1(n_971),
.A2(n_869),
.B(n_858),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1039),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_932),
.A2(n_914),
.B(n_795),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_981),
.Y(n_1179)
);

BUFx4f_ASAP7_75t_SL g1180 ( 
.A(n_1069),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1159),
.B(n_1161),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1064),
.A2(n_1167),
.B(n_1166),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1109),
.Y(n_1183)
);

BUFx4_ASAP7_75t_SL g1184 ( 
.A(n_1091),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1084),
.A2(n_1060),
.B(n_1103),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1162),
.B(n_1053),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1178),
.A2(n_1120),
.B(n_1050),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1067),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1165),
.A2(n_1117),
.B(n_1163),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1085),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1066),
.A2(n_1158),
.B(n_1157),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1171),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1116),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1164),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_SL g1195 ( 
.A1(n_1176),
.A2(n_1143),
.B(n_1125),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1163),
.A2(n_1062),
.B1(n_1073),
.B2(n_1128),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1074),
.Y(n_1197)
);

AOI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1145),
.A2(n_1143),
.B1(n_1095),
.B2(n_1127),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1157),
.A2(n_1158),
.B(n_1081),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1062),
.A2(n_1140),
.B1(n_1071),
.B2(n_1093),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_SL g1201 ( 
.A1(n_1125),
.A2(n_1130),
.B(n_1144),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1085),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1082),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_1103),
.A2(n_1131),
.B(n_1092),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1140),
.A2(n_1147),
.B1(n_1133),
.B2(n_1083),
.Y(n_1205)
);

AND2x6_ASAP7_75t_L g1206 ( 
.A(n_1070),
.B(n_1076),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1049),
.B(n_1097),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1049),
.B(n_1065),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1147),
.A2(n_1075),
.B1(n_1175),
.B2(n_1055),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1092),
.A2(n_1173),
.B(n_1172),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1088),
.B(n_1100),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1097),
.B(n_1112),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1078),
.B(n_1070),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1048),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1051),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1089),
.A2(n_1072),
.B(n_1057),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1118),
.B(n_1056),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1079),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1104),
.A2(n_1135),
.B(n_1139),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1058),
.A2(n_1077),
.B(n_1115),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1057),
.A2(n_1168),
.B(n_1094),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1113),
.A2(n_1122),
.B1(n_1114),
.B2(n_1076),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1080),
.A2(n_1068),
.A3(n_1096),
.B(n_1130),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1056),
.B(n_1113),
.Y(n_1224)
);

OAI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1052),
.A2(n_1065),
.B1(n_1122),
.B2(n_1061),
.C(n_1110),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1099),
.A2(n_1108),
.B(n_1138),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1052),
.B(n_1179),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1098),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1141),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1102),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1151),
.B(n_1170),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1132),
.A2(n_1114),
.B1(n_1131),
.B2(n_1134),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_SL g1233 ( 
.A(n_1154),
.B(n_1087),
.C(n_1086),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1151),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1156),
.B(n_1105),
.Y(n_1236)
);

OR3x4_ASAP7_75t_SL g1237 ( 
.A(n_1105),
.B(n_1175),
.C(n_1177),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1090),
.A2(n_1110),
.B(n_1126),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1082),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1051),
.Y(n_1240)
);

AOI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1059),
.A2(n_1126),
.B(n_1142),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1149),
.A2(n_1059),
.A3(n_1148),
.B(n_1054),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1153),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1051),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1148),
.A2(n_1054),
.A3(n_1106),
.B(n_1137),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1150),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1146),
.A2(n_1054),
.B(n_1137),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1106),
.A2(n_1107),
.B(n_1152),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1175),
.A2(n_1129),
.B(n_1174),
.C(n_1169),
.Y(n_1249)
);

NOR2x1_ASAP7_75t_SL g1250 ( 
.A(n_1111),
.B(n_1136),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1107),
.A2(n_1124),
.B(n_1155),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1121),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1119),
.B(n_1155),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1101),
.A2(n_1177),
.B1(n_1119),
.B2(n_1124),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1101),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1177),
.A2(n_1111),
.B1(n_1123),
.B2(n_1136),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1136),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1123),
.B(n_1162),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1162),
.B(n_1053),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1159),
.A2(n_1161),
.B(n_1165),
.Y(n_1260)
);

NAND2x1p5_ASAP7_75t_L g1261 ( 
.A(n_1088),
.B(n_800),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1163),
.A2(n_1062),
.B1(n_888),
.B2(n_1000),
.Y(n_1262)
);

OR2x6_ASAP7_75t_L g1263 ( 
.A(n_1103),
.B(n_1145),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1159),
.A2(n_1161),
.B(n_888),
.C(n_1165),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1162),
.B(n_1053),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1116),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1163),
.A2(n_888),
.B1(n_1062),
.B2(n_1073),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_1159),
.B(n_1161),
.C(n_440),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1069),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1112),
.B(n_1008),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1159),
.A2(n_1161),
.B1(n_777),
.B2(n_888),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1159),
.A2(n_1161),
.B1(n_777),
.B2(n_888),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1084),
.A2(n_1089),
.B(n_1092),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1085),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1069),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1084),
.A2(n_1060),
.B(n_1103),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1063),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1063),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1159),
.A2(n_1161),
.B1(n_777),
.B2(n_888),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1175),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1164),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1166),
.A2(n_1178),
.B(n_1167),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1063),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1049),
.B(n_1162),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1069),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1158),
.B(n_1160),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1064),
.A2(n_1167),
.B(n_1166),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1049),
.B(n_1162),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1166),
.A2(n_1178),
.B(n_1167),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1088),
.B(n_800),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1159),
.B(n_1161),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1063),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1166),
.A2(n_1178),
.B(n_1167),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1103),
.B(n_1145),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1162),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1159),
.A2(n_1161),
.B(n_1165),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1239),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1186),
.B(n_1259),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1197),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1217),
.B(n_1224),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1185),
.A2(n_1276),
.B(n_1273),
.Y(n_1301)
);

NOR2x1_ASAP7_75t_SL g1302 ( 
.A(n_1263),
.B(n_1294),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1208),
.B(n_1235),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1185),
.A2(n_1276),
.B(n_1273),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1208),
.B(n_1235),
.Y(n_1305)
);

NOR2xp67_ASAP7_75t_L g1306 ( 
.A(n_1295),
.B(n_1193),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1265),
.B(n_1284),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1207),
.B(n_1212),
.Y(n_1308)
);

O2A1O1Ixp5_ASAP7_75t_L g1309 ( 
.A1(n_1181),
.A2(n_1291),
.B(n_1189),
.C(n_1279),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1184),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1295),
.B(n_1258),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1200),
.B(n_1288),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1200),
.B(n_1196),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1248),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1267),
.A2(n_1196),
.B1(n_1205),
.B2(n_1209),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1248),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1280),
.B(n_1228),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1210),
.A2(n_1191),
.B(n_1199),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1214),
.Y(n_1319)
);

INVx5_ASAP7_75t_L g1320 ( 
.A(n_1263),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1268),
.A2(n_1279),
.B(n_1272),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1210),
.A2(n_1189),
.B(n_1271),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1222),
.B(n_1267),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1270),
.B(n_1188),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1271),
.A2(n_1272),
.B(n_1264),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1192),
.B(n_1292),
.Y(n_1326)
);

O2A1O1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1262),
.A2(n_1264),
.B(n_1181),
.C(n_1291),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1229),
.B(n_1277),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1262),
.A2(n_1296),
.B(n_1260),
.C(n_1232),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1227),
.B(n_1190),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_R g1331 ( 
.A(n_1218),
.B(n_1234),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1260),
.A2(n_1296),
.B(n_1221),
.C(n_1216),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1229),
.B(n_1278),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1242),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1190),
.B(n_1202),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1183),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1242),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1220),
.B(n_1198),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_SL g1339 ( 
.A(n_1281),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1202),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1233),
.A2(n_1294),
.B1(n_1211),
.B2(n_1225),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1221),
.A2(n_1216),
.B1(n_1204),
.B2(n_1238),
.C(n_1201),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1249),
.A2(n_1220),
.B(n_1250),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1213),
.A2(n_1266),
.B1(n_1249),
.B2(n_1261),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1242),
.Y(n_1345)
);

NOR2xp67_ASAP7_75t_L g1346 ( 
.A(n_1283),
.B(n_1252),
.Y(n_1346)
);

OR2x6_ASAP7_75t_L g1347 ( 
.A(n_1213),
.B(n_1195),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1255),
.B(n_1243),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1274),
.B(n_1223),
.Y(n_1349)
);

AND2x6_ASAP7_75t_L g1350 ( 
.A(n_1280),
.B(n_1246),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1203),
.A2(n_1236),
.B(n_1237),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1184),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1223),
.B(n_1257),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1261),
.A2(n_1290),
.B1(n_1285),
.B2(n_1256),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1238),
.A2(n_1290),
.B(n_1231),
.C(n_1240),
.Y(n_1355)
);

INVxp33_ASAP7_75t_L g1356 ( 
.A(n_1236),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1206),
.B(n_1223),
.Y(n_1357)
);

BUFx2_ASAP7_75t_SL g1358 ( 
.A(n_1269),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_SL g1359 ( 
.A1(n_1245),
.A2(n_1223),
.B(n_1251),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1215),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1206),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1206),
.B(n_1194),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1245),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1253),
.A2(n_1275),
.B(n_1254),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1206),
.Y(n_1365)
);

INVxp33_ASAP7_75t_SL g1366 ( 
.A(n_1230),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1285),
.A2(n_1180),
.B1(n_1253),
.B2(n_1244),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_1244),
.B(n_1241),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1219),
.A2(n_1187),
.B(n_1293),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1206),
.B(n_1244),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_SL g1371 ( 
.A1(n_1245),
.A2(n_1286),
.B(n_1247),
.Y(n_1371)
);

AOI21x1_ASAP7_75t_SL g1372 ( 
.A1(n_1245),
.A2(n_1247),
.B(n_1226),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1180),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1182),
.B(n_1287),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1282),
.B(n_1289),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1186),
.B(n_1259),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1200),
.A2(n_993),
.B1(n_1196),
.B2(n_1267),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1217),
.B(n_1224),
.Y(n_1378)
);

O2A1O1Ixp5_ASAP7_75t_L g1379 ( 
.A1(n_1181),
.A2(n_1161),
.B(n_1159),
.C(n_1291),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1197),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1217),
.B(n_1224),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1210),
.A2(n_1191),
.B(n_1199),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1186),
.B(n_1259),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1207),
.B(n_1212),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1237),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1217),
.B(n_1224),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1284),
.B(n_1288),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1267),
.A2(n_1196),
.B1(n_1200),
.B2(n_1161),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1322),
.B(n_1321),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1330),
.B(n_1340),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1361),
.B(n_1365),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1314),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1297),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1297),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_1316),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1334),
.B(n_1345),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1377),
.A2(n_1315),
.B1(n_1388),
.B2(n_1313),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1320),
.B(n_1302),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1299),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1335),
.B(n_1303),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1301),
.A2(n_1304),
.B(n_1332),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1349),
.B(n_1380),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1320),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1316),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1374),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1319),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1305),
.B(n_1323),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1369),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1347),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1375),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1353),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1357),
.B(n_1320),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1369),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1311),
.B(n_1337),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1332),
.B(n_1312),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1375),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1342),
.A2(n_1309),
.B(n_1379),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1363),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1318),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_SL g1421 ( 
.A1(n_1327),
.A2(n_1355),
.B(n_1341),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1347),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1318),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1368),
.A2(n_1362),
.B(n_1344),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1350),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1300),
.B(n_1378),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1382),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_L g1428 ( 
.A(n_1343),
.B(n_1370),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1381),
.B(n_1386),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1336),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1338),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1364),
.B(n_1385),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1309),
.B(n_1328),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1333),
.B(n_1387),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1307),
.B(n_1384),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1350),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1379),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1406),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1396),
.B(n_1410),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1393),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1408),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1396),
.B(n_1298),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1433),
.B(n_1326),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1396),
.B(n_1383),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1433),
.B(n_1348),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1392),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1404),
.B(n_1308),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1400),
.B(n_1376),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1410),
.B(n_1308),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1389),
.A2(n_1306),
.B(n_1346),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1394),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1397),
.A2(n_1385),
.B1(n_1339),
.B2(n_1324),
.Y(n_1452)
);

AND2x2_ASAP7_75t_SL g1453 ( 
.A(n_1418),
.B(n_1385),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1400),
.B(n_1350),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1398),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1430),
.Y(n_1456)
);

NOR4xp25_ASAP7_75t_SL g1457 ( 
.A(n_1436),
.B(n_1310),
.C(n_1360),
.D(n_1351),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1417),
.B(n_1372),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1417),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1404),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1405),
.B(n_1317),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1395),
.B(n_1371),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1395),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1412),
.B(n_1359),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1405),
.B(n_1356),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1399),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1441),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1450),
.A2(n_1389),
.B1(n_1411),
.B2(n_1432),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1449),
.B(n_1413),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1450),
.B(n_1389),
.C(n_1411),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1452),
.A2(n_1389),
.B1(n_1421),
.B2(n_1418),
.Y(n_1472)
);

OAI33xp33_ASAP7_75t_L g1473 ( 
.A1(n_1464),
.A2(n_1407),
.A3(n_1390),
.B1(n_1412),
.B2(n_1419),
.B3(n_1434),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1449),
.B(n_1413),
.Y(n_1474)
);

AO221x2_ASAP7_75t_L g1475 ( 
.A1(n_1454),
.A2(n_1407),
.B1(n_1437),
.B2(n_1389),
.C(n_1367),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1466),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1452),
.A2(n_1432),
.B1(n_1428),
.B2(n_1418),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_R g1478 ( 
.A(n_1456),
.B(n_1339),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1456),
.A2(n_1432),
.B1(n_1428),
.B2(n_1418),
.Y(n_1479)
);

OAI211xp5_ASAP7_75t_L g1480 ( 
.A1(n_1438),
.A2(n_1401),
.B(n_1418),
.C(n_1416),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1453),
.A2(n_1421),
.B(n_1432),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1453),
.A2(n_1432),
.B1(n_1435),
.B2(n_1430),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1453),
.A2(n_1416),
.B1(n_1422),
.B2(n_1409),
.Y(n_1483)
);

OAI211xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1438),
.A2(n_1406),
.B(n_1390),
.C(n_1434),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1448),
.A2(n_1435),
.B1(n_1354),
.B2(n_1422),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1443),
.B(n_1426),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1441),
.A2(n_1414),
.B(n_1423),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1460),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1460),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_SL g1490 ( 
.A(n_1455),
.B(n_1447),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1455),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1445),
.A2(n_1429),
.B1(n_1448),
.B2(n_1443),
.C(n_1437),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1440),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1449),
.B(n_1415),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1455),
.A2(n_1352),
.B1(n_1366),
.B2(n_1358),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1454),
.A2(n_1424),
.B(n_1399),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1455),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1445),
.A2(n_1437),
.B1(n_1426),
.B2(n_1409),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1447),
.A2(n_1425),
.B1(n_1436),
.B2(n_1403),
.Y(n_1499)
);

OAI211xp5_ASAP7_75t_L g1500 ( 
.A1(n_1465),
.A2(n_1461),
.B(n_1457),
.C(n_1462),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1461),
.B(n_1402),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1447),
.A2(n_1425),
.B1(n_1403),
.B2(n_1356),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1440),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1440),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1464),
.B(n_1391),
.C(n_1431),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1451),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1496),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1493),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1487),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1492),
.B(n_1398),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1503),
.Y(n_1511)
);

OAI21xp33_ASAP7_75t_L g1512 ( 
.A1(n_1480),
.A2(n_1465),
.B(n_1462),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1467),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1504),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1506),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1469),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1476),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1497),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1479),
.B(n_1462),
.C(n_1457),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1471),
.B(n_1481),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1486),
.B(n_1373),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1505),
.A2(n_1427),
.B(n_1420),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1458),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1478),
.B(n_1398),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1497),
.Y(n_1525)
);

NAND2x1_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1459),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1488),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1489),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1478),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1475),
.Y(n_1530)
);

NOR3xp33_ASAP7_75t_SL g1531 ( 
.A(n_1495),
.B(n_1500),
.C(n_1484),
.Y(n_1531)
);

INVx4_ASAP7_75t_SL g1532 ( 
.A(n_1475),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1470),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1494),
.B(n_1439),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1474),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1512),
.B(n_1485),
.Y(n_1536)
);

NAND4xp25_ASAP7_75t_L g1537 ( 
.A(n_1519),
.B(n_1472),
.C(n_1468),
.D(n_1477),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1512),
.B(n_1498),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1509),
.Y(n_1539)
);

NAND4xp25_ASAP7_75t_L g1540 ( 
.A(n_1519),
.B(n_1472),
.C(n_1529),
.D(n_1507),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1523),
.B(n_1475),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1509),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1508),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1527),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1509),
.Y(n_1545)
);

BUFx2_ASAP7_75t_SL g1546 ( 
.A(n_1529),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1527),
.B(n_1501),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1531),
.B(n_1482),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1523),
.B(n_1498),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1511),
.Y(n_1552)
);

AND3x2_ASAP7_75t_L g1553 ( 
.A(n_1507),
.B(n_1463),
.C(n_1459),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1511),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1530),
.B(n_1531),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1524),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1528),
.Y(n_1557)
);

AND2x4_ASAP7_75t_SL g1558 ( 
.A(n_1523),
.B(n_1398),
.Y(n_1558)
);

NOR2x1_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1530),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1532),
.B(n_1442),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1514),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1514),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1515),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1515),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1526),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1528),
.B(n_1446),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1530),
.B(n_1510),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1516),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1521),
.B(n_1442),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1532),
.B(n_1442),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1532),
.B(n_1444),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1517),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1444),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1517),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1550),
.B(n_1331),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1539),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1569),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1569),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1546),
.B(n_1520),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1573),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1546),
.B(n_1533),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1532),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1555),
.A2(n_1520),
.B(n_1518),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1539),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1536),
.B(n_1532),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1568),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1574),
.B(n_1520),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1541),
.B(n_1520),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1540),
.B(n_1520),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1573),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1520),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1557),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1575),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1556),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1533),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1575),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_L g1599 ( 
.A(n_1559),
.B(n_1525),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1538),
.B(n_1535),
.Y(n_1600)
);

INVxp33_ASAP7_75t_L g1601 ( 
.A(n_1537),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1570),
.B(n_1535),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1549),
.B(n_1513),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1559),
.A2(n_1499),
.B1(n_1502),
.B2(n_1518),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1566),
.B(n_1522),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1549),
.B(n_1513),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1542),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1566),
.B(n_1571),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1560),
.B(n_1534),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1518),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1579),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1608),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1597),
.B(n_1548),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1596),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1580),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1608),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1601),
.A2(n_1537),
.B1(n_1551),
.B2(n_1548),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1601),
.B(n_1551),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1584),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1597),
.B(n_1558),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1599),
.B(n_1566),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1605),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1583),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1610),
.B(n_1584),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1608),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1610),
.B(n_1558),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1592),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1591),
.A2(n_1572),
.B1(n_1502),
.B2(n_1525),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1588),
.B(n_1572),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1595),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1581),
.A2(n_1525),
.B1(n_1567),
.B2(n_1554),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1598),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1543),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1617),
.A2(n_1585),
.B1(n_1587),
.B2(n_1604),
.C(n_1590),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1625),
.B(n_1590),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1622),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1614),
.B(n_1619),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1618),
.A2(n_1629),
.B1(n_1625),
.B2(n_1613),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1616),
.Y(n_1641)
);

INVx2_ASAP7_75t_R g1642 ( 
.A(n_1611),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1611),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1615),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1624),
.A2(n_1576),
.B(n_1594),
.C(n_1578),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1613),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1615),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1624),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1622),
.A2(n_1633),
.B(n_1630),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1620),
.A2(n_1578),
.B1(n_1594),
.B2(n_1593),
.C(n_1609),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1622),
.A2(n_1593),
.B(n_1602),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1612),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1635),
.A2(n_1589),
.B1(n_1473),
.B2(n_1553),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1620),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_1635),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_R g1656 ( 
.A(n_1648),
.B(n_1639),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1638),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1641),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1641),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1645),
.B(n_1626),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1637),
.B(n_1621),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1642),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1638),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1642),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1640),
.B(n_1589),
.Y(n_1665)
);

OAI32xp33_ASAP7_75t_L g1666 ( 
.A1(n_1662),
.A2(n_1653),
.A3(n_1626),
.B1(n_1612),
.B2(n_1649),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1660),
.A2(n_1636),
.B1(n_1650),
.B2(n_1653),
.C(n_1664),
.Y(n_1667)
);

OAI21xp33_ASAP7_75t_L g1668 ( 
.A1(n_1656),
.A2(n_1651),
.B(n_1621),
.Y(n_1668)
);

NOR3xp33_ASAP7_75t_SL g1669 ( 
.A(n_1660),
.B(n_1659),
.C(n_1658),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1657),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1661),
.B(n_1652),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_SL g1672 ( 
.A1(n_1665),
.A2(n_1654),
.B1(n_1647),
.B2(n_1644),
.C(n_1643),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1655),
.A2(n_1622),
.B(n_1616),
.C(n_1612),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1663),
.A2(n_1627),
.B1(n_1626),
.B2(n_1612),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1670),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1671),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_SL g1677 ( 
.A(n_1669),
.B(n_1657),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_SL g1678 ( 
.A(n_1668),
.B(n_1626),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1667),
.A2(n_1627),
.B1(n_1657),
.B2(n_1632),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1677),
.B(n_1673),
.C(n_1666),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1675),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1678),
.B(n_1672),
.C(n_1674),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1676),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1679),
.B(n_1628),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1675),
.Y(n_1685)
);

AOI211x1_ASAP7_75t_SL g1686 ( 
.A1(n_1682),
.A2(n_1632),
.B(n_1623),
.C(n_1577),
.Y(n_1686)
);

AOI321xp33_ASAP7_75t_L g1687 ( 
.A1(n_1680),
.A2(n_1632),
.A3(n_1623),
.B1(n_1631),
.B2(n_1628),
.C(n_1634),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1681),
.B(n_1623),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1685),
.B(n_1631),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1684),
.B(n_1634),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1686),
.B(n_1683),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1688),
.B(n_1577),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1689),
.Y(n_1693)
);

XNOR2xp5_ASAP7_75t_L g1694 ( 
.A(n_1691),
.B(n_1690),
.Y(n_1694)
);

OAI322xp33_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1693),
.A3(n_1692),
.B1(n_1687),
.B2(n_1605),
.C1(n_1586),
.C2(n_1607),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1695),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1696),
.B(n_1586),
.Y(n_1697)
);

OAI22x1_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1607),
.B1(n_1542),
.B2(n_1545),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1545),
.B1(n_1606),
.B2(n_1603),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1698),
.A2(n_1606),
.B1(n_1603),
.B2(n_1564),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1543),
.B(n_1562),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1699),
.B(n_1547),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1701),
.B(n_1702),
.Y(n_1703)
);

AOI22x1_ASAP7_75t_L g1704 ( 
.A1(n_1701),
.A2(n_1552),
.B1(n_1562),
.B2(n_1554),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1703),
.A2(n_1547),
.B1(n_1552),
.B2(n_1564),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1705),
.A2(n_1704),
.B1(n_1563),
.B2(n_1565),
.C(n_1509),
.Y(n_1706)
);

AOI211xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1563),
.B(n_1565),
.C(n_1567),
.Y(n_1707)
);


endmodule