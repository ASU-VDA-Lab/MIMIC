module fake_netlist_6_2969_n_1205 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1205);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1205;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_208;
wire n_1033;
wire n_1052;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_1101;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_718;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_923;
wire n_504;
wire n_1078;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_174;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_886;
wire n_343;
wire n_953;
wire n_448;
wire n_1094;
wire n_1017;
wire n_1106;
wire n_1004;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_228;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_811;
wire n_312;
wire n_394;
wire n_630;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_880;
wire n_792;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_1198;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_201;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_221;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_1154;
wire n_437;
wire n_1082;
wire n_259;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1177;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

INVx1_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_47),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_18),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_39),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_56),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_69),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_57),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_38),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_76),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_61),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_9),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_6),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_38),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_136),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_35),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_25),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_67),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_23),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_7),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_5),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_79),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_65),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_149),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_43),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_98),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_82),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_152),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_30),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_160),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_145),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_44),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_117),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_171),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_55),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_42),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_27),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_184),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_187),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_188),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_190),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_191),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_192),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_196),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_202),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_205),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_174),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_200),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_214),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_215),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_234),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_240),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_242),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_246),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_249),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_253),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_254),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_258),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_233),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_243),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_247),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_247),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_230),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_230),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_259),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_259),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_265),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_265),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_266),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_274),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_262),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_274),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_284),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_275),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_270),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_305),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_311),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_267),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_284),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_289),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_271),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_272),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_291),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_273),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_270),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_270),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_292),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_292),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_260),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_356),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_293),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_318),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_314),
.B(n_300),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_314),
.B(n_300),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_347),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_293),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_312),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_319),
.B(n_294),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_315),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_321),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_301),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_324),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_323),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_294),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_327),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_325),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_344),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_334),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

OAI22x1_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_307),
.B1(n_310),
.B2(n_260),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_320),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_320),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_333),
.B(n_322),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_322),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_333),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_361),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_377),
.A2(n_307),
.B1(n_310),
.B2(n_336),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_338),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_372),
.A2(n_341),
.B(n_338),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_385),
.A2(n_290),
.B1(n_342),
.B2(n_341),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_395),
.A2(n_339),
.B1(n_331),
.B2(n_358),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_342),
.B1(n_337),
.B2(n_340),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_375),
.A2(n_348),
.B(n_328),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

NOR2x1_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_303),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_376),
.B(n_346),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_369),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_377),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_329),
.Y(n_449)
);

BUFx12f_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_386),
.A2(n_339),
.B1(n_331),
.B2(n_354),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_304),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_382),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_403),
.B(n_299),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_399),
.Y(n_458)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_399),
.B(n_213),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_403),
.B(n_179),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_373),
.B(n_352),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_373),
.A2(n_301),
.B1(n_296),
.B2(n_217),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_361),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_394),
.B(n_180),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_385),
.A2(n_296),
.B1(n_224),
.B2(n_302),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_363),
.B(n_329),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_385),
.A2(n_198),
.B1(n_182),
.B2(n_185),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_363),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_361),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_385),
.A2(n_201),
.B1(n_195),
.B2(n_197),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_363),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_363),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_377),
.Y(n_475)
);

CKINVDCx6p67_ASAP7_75t_R g476 ( 
.A(n_384),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_385),
.B(n_176),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_361),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_361),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_383),
.A2(n_199),
.B(n_286),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_361),
.Y(n_482)
);

CKINVDCx6p67_ASAP7_75t_R g483 ( 
.A(n_384),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_363),
.B(n_288),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_411),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_431),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_446),
.B(n_288),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_431),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_349),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_464),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_438),
.A2(n_295),
.B(n_349),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_419),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_424),
.B(n_418),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_416),
.Y(n_499)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_464),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_288),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_469),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_424),
.B(n_349),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_476),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_193),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_418),
.B(n_439),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_418),
.B(n_45),
.Y(n_509)
);

INVxp33_ASAP7_75t_SL g510 ( 
.A(n_422),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_450),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_444),
.B(n_445),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_467),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_481),
.A2(n_219),
.B(n_218),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_471),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_467),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_426),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_427),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_437),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_437),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_175),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_432),
.B(n_175),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_439),
.B(n_225),
.Y(n_528)
);

AND3x2_ASAP7_75t_L g529 ( 
.A(n_441),
.B(n_178),
.C(n_177),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_418),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_501),
.A2(n_459),
.B1(n_449),
.B2(n_453),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_498),
.A2(n_459),
.B1(n_449),
.B2(n_453),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_498),
.A2(n_475),
.B1(n_448),
.B2(n_455),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_498),
.A2(n_475),
.B1(n_448),
.B2(n_455),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_520),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g536 ( 
.A(n_514),
.B(n_509),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_L g537 ( 
.A1(n_516),
.A2(n_458),
.B1(n_436),
.B2(n_457),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_SL g538 ( 
.A1(n_527),
.A2(n_456),
.B1(n_458),
.B2(n_466),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_498),
.A2(n_484),
.B1(n_461),
.B2(n_433),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_515),
.B(n_484),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_514),
.B(n_450),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_510),
.A2(n_487),
.B1(n_528),
.B2(n_458),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_519),
.A2(n_405),
.B1(n_439),
.B2(n_461),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_504),
.A2(n_451),
.B1(n_405),
.B2(n_435),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_506),
.B(n_454),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_490),
.B(n_447),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_505),
.A2(n_439),
.B1(n_447),
.B2(n_468),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_515),
.A2(n_462),
.B1(n_415),
.B2(n_420),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_489),
.A2(n_471),
.B1(n_423),
.B2(n_434),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_485),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

AO22x2_ASAP7_75t_L g552 ( 
.A1(n_485),
.A2(n_470),
.B1(n_478),
.B2(n_463),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_488),
.A2(n_407),
.B1(n_410),
.B2(n_406),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_492),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_506),
.B(n_435),
.Y(n_555)
);

OA22x2_ASAP7_75t_L g556 ( 
.A1(n_486),
.A2(n_491),
.B1(n_502),
.B2(n_529),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_509),
.A2(n_454),
.B1(n_452),
.B2(n_483),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_443),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_526),
.B(n_454),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_442),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_511),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_493),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_490),
.B(n_471),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_511),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_493),
.A2(n_482),
.B1(n_480),
.B2(n_479),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_511),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_511),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_495),
.A2(n_428),
.B1(n_460),
.B2(n_472),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_495),
.A2(n_483),
.B1(n_476),
.B2(n_430),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_535),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_555),
.B(n_496),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_551),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_531),
.A2(n_452),
.B1(n_460),
.B2(n_440),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_550),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_563),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_554),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_566),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_552),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_562),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_561),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_545),
.B(n_412),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_565),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_565),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_548),
.A2(n_494),
.B(n_517),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_460),
.C(n_477),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

INVx4_ASAP7_75t_SL g590 ( 
.A(n_563),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_558),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_561),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_L g593 ( 
.A(n_543),
.B(n_477),
.C(n_452),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_569),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_532),
.B(n_412),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_540),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_549),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_559),
.A2(n_465),
.B1(n_423),
.B2(n_434),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_560),
.B(n_409),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_538),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_546),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_557),
.B(n_508),
.Y(n_603)
);

AO21x2_ASAP7_75t_L g604 ( 
.A1(n_553),
.A2(n_494),
.B(n_438),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_537),
.B(n_423),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_546),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_536),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_539),
.B(n_409),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

INVxp67_ASAP7_75t_SL g611 ( 
.A(n_547),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_570),
.Y(n_612)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_533),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_567),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_534),
.B(n_509),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_550),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_536),
.B(n_496),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_555),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_531),
.B(n_423),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_550),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_550),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_531),
.B(n_430),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_535),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_545),
.B(n_412),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_545),
.B(n_409),
.Y(n_634)
);

OAI22xp33_ASAP7_75t_SL g635 ( 
.A1(n_531),
.A2(n_178),
.B1(n_204),
.B2(n_177),
.Y(n_635)
);

AND3x1_ASAP7_75t_L g636 ( 
.A(n_541),
.B(n_474),
.C(n_421),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_563),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_536),
.B(n_497),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_535),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_544),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_535),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_563),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_L g643 ( 
.A(n_549),
.B(n_508),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_558),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_535),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_531),
.B(n_430),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_531),
.B(n_430),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_536),
.B(n_497),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_617),
.B(n_509),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_621),
.B(n_507),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_573),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_619),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_625),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_619),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_591),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_600),
.B(n_507),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_623),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_623),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_626),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_626),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_628),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_581),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_592),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_530),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_628),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_588),
.B(n_434),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_610),
.Y(n_672)
);

INVx4_ASAP7_75t_SL g673 ( 
.A(n_625),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_592),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_632),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_632),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_572),
.B(n_465),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_572),
.B(n_512),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_592),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_618),
.A2(n_434),
.B1(n_229),
.B2(n_204),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_620),
.B(n_465),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_592),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_512),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_633),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_580),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_593),
.B(n_530),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_633),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_591),
.B(n_530),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_576),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_581),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_571),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_521),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_638),
.B(n_521),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_580),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_638),
.B(n_522),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_522),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_584),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_592),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_652),
.B(n_523),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_571),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_590),
.B(n_490),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_590),
.B(n_607),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_649),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_625),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_625),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_586),
.Y(n_707)
);

AND3x4_ASAP7_75t_L g708 ( 
.A(n_607),
.B(n_474),
.C(n_421),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_591),
.B(n_530),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_608),
.B(n_523),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_585),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_649),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_601),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_583),
.B(n_421),
.Y(n_714)
);

BUFx4f_ASAP7_75t_L g715 ( 
.A(n_625),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_637),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_586),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_601),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_645),
.B(n_530),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_637),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_585),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_574),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_637),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_617),
.B(n_499),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_645),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_594),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_596),
.B(n_524),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_594),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_637),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_596),
.B(n_524),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_645),
.B(n_413),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_637),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_608),
.B(n_525),
.Y(n_733)
);

OAI221xp5_ASAP7_75t_L g734 ( 
.A1(n_575),
.A2(n_229),
.B1(n_203),
.B2(n_206),
.C(n_207),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_613),
.B(n_609),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_574),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_578),
.Y(n_737)
);

CKINVDCx6p67_ASAP7_75t_R g738 ( 
.A(n_610),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_649),
.B(n_474),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_725),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_735),
.B(n_610),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_735),
.B(n_618),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_713),
.B(n_589),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_726),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_728),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_658),
.Y(n_746)
);

AND2x6_ASAP7_75t_L g747 ( 
.A(n_702),
.B(n_612),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_712),
.B(n_618),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_692),
.B(n_602),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_712),
.B(n_612),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_715),
.A2(n_643),
.B(n_603),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_660),
.B(n_640),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_667),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_672),
.A2(n_627),
.B1(n_647),
.B2(n_622),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_689),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_685),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_689),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_654),
.Y(n_758)
);

XOR2xp5_ASAP7_75t_L g759 ( 
.A(n_681),
.B(n_636),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_674),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_685),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_694),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_714),
.B(n_635),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_696),
.B(n_602),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_738),
.B(n_672),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_697),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_704),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_693),
.B(n_615),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_704),
.B(n_640),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_690),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_714),
.B(n_648),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_695),
.B(n_615),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_658),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_700),
.Y(n_774)
);

INVxp33_ASAP7_75t_L g775 ( 
.A(n_708),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_683),
.B(n_631),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_691),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_699),
.B(n_615),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_658),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_734),
.A2(n_650),
.B1(n_589),
.B2(n_595),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_658),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_678),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_713),
.B(n_598),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_718),
.B(n_598),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_718),
.B(n_614),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_655),
.B(n_614),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_691),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_737),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_739),
.B(n_634),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_653),
.B(n_669),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_661),
.B(n_616),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_705),
.B(n_616),
.Y(n_792)
);

BUFx6f_ASAP7_75t_SL g793 ( 
.A(n_668),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_703),
.B(n_648),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_677),
.B(n_577),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_655),
.B(n_614),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_703),
.B(n_715),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_710),
.B(n_614),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_668),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_671),
.B(n_606),
.C(n_599),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_708),
.B(n_577),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_733),
.B(n_614),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_680),
.B(n_702),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_680),
.B(n_648),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_705),
.B(n_651),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_673),
.B(n_590),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_653),
.A2(n_671),
.B1(n_686),
.B2(n_724),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_707),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_717),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_662),
.B(n_578),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_716),
.B(n_577),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_737),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_782),
.B(n_721),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_790),
.B(n_711),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_758),
.B(n_711),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_781),
.B(n_669),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_768),
.B(n_656),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_767),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_776),
.B(n_686),
.C(n_688),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_783),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_740),
.B(n_724),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_755),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_748),
.A2(n_603),
.B1(n_653),
.B2(n_724),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_772),
.B(n_657),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_744),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_745),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_762),
.Y(n_827)
);

OAI221xp5_ASAP7_75t_L g828 ( 
.A1(n_763),
.A2(n_210),
.B1(n_208),
.B2(n_220),
.C(n_688),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_799),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_742),
.A2(n_724),
.B1(n_176),
.B2(n_669),
.Y(n_830)
);

AND2x2_ASAP7_75t_SL g831 ( 
.A(n_806),
.B(n_705),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_741),
.B(n_709),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_778),
.B(n_659),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_757),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_756),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_790),
.B(n_716),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_750),
.B(n_709),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_746),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_746),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_749),
.B(n_663),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_770),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_766),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_753),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_748),
.A2(n_724),
.B1(n_624),
.B2(n_642),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_764),
.B(n_664),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_774),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_798),
.B(n_665),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_743),
.B(n_719),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_743),
.B(n_719),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_780),
.A2(n_176),
.B1(n_642),
.B2(n_624),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_746),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_802),
.B(n_666),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_808),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_791),
.B(n_731),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_773),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_761),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_803),
.A2(n_624),
.B1(n_642),
.B2(n_651),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_754),
.B(n_751),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_747),
.B(n_705),
.Y(n_859)
);

AOI221xp5_ASAP7_75t_L g860 ( 
.A1(n_804),
.A2(n_176),
.B1(n_225),
.B2(n_226),
.C(n_227),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_795),
.B(n_731),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_785),
.B(n_684),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_765),
.B(n_706),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_801),
.B(n_706),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_800),
.A2(n_730),
.B(n_727),
.C(n_643),
.Y(n_866)
);

AND2x6_ASAP7_75t_SL g867 ( 
.A(n_752),
.B(n_736),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_789),
.B(n_651),
.C(n_720),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_809),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_786),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_785),
.B(n_687),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_SL g872 ( 
.A(n_775),
.B(n_706),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_783),
.B(n_784),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_806),
.B(n_706),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_777),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_796),
.B(n_670),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_787),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_771),
.B(n_723),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_788),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_807),
.B(n_723),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_790),
.B(n_796),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_784),
.B(n_675),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_812),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_810),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_810),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_811),
.B(n_723),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_825),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_870),
.Y(n_888)
);

AO22x2_ASAP7_75t_L g889 ( 
.A1(n_880),
.A2(n_805),
.B1(n_759),
.B2(n_676),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_873),
.B(n_676),
.Y(n_890)
);

OAI221xp5_ASAP7_75t_L g891 ( 
.A1(n_858),
.A2(n_769),
.B1(n_794),
.B2(n_792),
.C(n_797),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_858),
.A2(n_747),
.B1(n_793),
.B2(n_720),
.Y(n_892)
);

BUFx8_ASAP7_75t_L g893 ( 
.A(n_829),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_880),
.A2(n_747),
.B1(n_732),
.B2(n_723),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_826),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_827),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_839),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_820),
.A2(n_673),
.B1(n_760),
.B2(n_732),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_881),
.B(n_779),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_842),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_848),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_848),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_849),
.B(n_701),
.Y(n_903)
);

AO22x2_ASAP7_75t_L g904 ( 
.A1(n_820),
.A2(n_673),
.B1(n_682),
.B2(n_722),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_L g905 ( 
.A(n_819),
.B(n_747),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_849),
.B(n_779),
.Y(n_906)
);

AO22x2_ASAP7_75t_L g907 ( 
.A1(n_846),
.A2(n_682),
.B1(n_698),
.B2(n_679),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_836),
.B(n_679),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_854),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_839),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_853),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_831),
.B(n_729),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_823),
.B(n_729),
.Y(n_913)
);

AO22x2_ASAP7_75t_L g914 ( 
.A1(n_869),
.A2(n_698),
.B1(n_590),
.B2(n_582),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_854),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_835),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_835),
.Y(n_917)
);

AO22x2_ASAP7_75t_L g918 ( 
.A1(n_868),
.A2(n_582),
.B1(n_605),
.B2(n_597),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_828),
.A2(n_729),
.B1(n_226),
.B2(n_227),
.C(n_228),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_885),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_815),
.B(n_729),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_850),
.A2(n_228),
.B1(n_605),
.B2(n_597),
.C(n_176),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_884),
.B(n_604),
.Y(n_923)
);

AO22x2_ASAP7_75t_L g924 ( 
.A1(n_868),
.A2(n_605),
.B1(n_597),
.B2(n_579),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_816),
.B(n_674),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_841),
.Y(n_926)
);

AO22x2_ASAP7_75t_L g927 ( 
.A1(n_856),
.A2(n_579),
.B1(n_630),
.B2(n_629),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_856),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_839),
.Y(n_929)
);

AO22x2_ASAP7_75t_L g930 ( 
.A1(n_813),
.A2(n_630),
.B1(n_646),
.B2(n_644),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_843),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_822),
.Y(n_932)
);

BUFx8_ASAP7_75t_L g933 ( 
.A(n_855),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_847),
.B(n_604),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_860),
.A2(n_850),
.B(n_857),
.C(n_866),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_832),
.B(n_837),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_837),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_892),
.B(n_832),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_937),
.B(n_861),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_909),
.B(n_861),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_893),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_936),
.B(n_915),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_935),
.A2(n_821),
.B(n_859),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_907),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_908),
.B(n_865),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_901),
.B(n_818),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_907),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_902),
.B(n_863),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_920),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_887),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_905),
.A2(n_830),
.B(n_878),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_L g952 ( 
.A1(n_889),
.A2(n_830),
.B(n_824),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_893),
.B(n_831),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_910),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_894),
.B(n_844),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_922),
.A2(n_872),
.B(n_864),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_919),
.A2(n_886),
.B(n_874),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_891),
.B(n_867),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_913),
.A2(n_833),
.B(n_817),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_889),
.A2(n_882),
.B(n_871),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_910),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_934),
.A2(n_916),
.B(n_928),
.C(n_917),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_887),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_908),
.B(n_814),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_903),
.A2(n_852),
.B(n_845),
.C(n_840),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_930),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_913),
.A2(n_814),
.B1(n_793),
.B2(n_838),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_918),
.A2(n_876),
.B(n_834),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_933),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_895),
.Y(n_970)
);

INVx5_ASAP7_75t_L g971 ( 
.A(n_913),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_918),
.A2(n_877),
.B(n_875),
.Y(n_972)
);

AOI21xp33_ASAP7_75t_L g973 ( 
.A1(n_924),
.A2(n_883),
.B(n_879),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_906),
.A2(n_923),
.B(n_921),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_890),
.B(n_851),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_896),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_899),
.B(n_862),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_925),
.B(n_838),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_888),
.B(n_862),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_900),
.B(n_911),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_912),
.A2(n_587),
.B(n_629),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_924),
.A2(n_855),
.B(n_517),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_914),
.A2(n_500),
.B1(n_855),
.B2(n_517),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_933),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_930),
.A2(n_855),
.B(n_517),
.Y(n_985)
);

NOR2x1_ASAP7_75t_L g986 ( 
.A(n_929),
.B(n_604),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_932),
.B(n_587),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_926),
.B(n_931),
.Y(n_988)
);

NAND2x1_ASAP7_75t_L g989 ( 
.A(n_898),
.B(n_904),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_927),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_927),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_910),
.B(n_500),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_897),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_892),
.B(n_500),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_907),
.Y(n_995)
);

BUFx4f_ASAP7_75t_L g996 ( 
.A(n_941),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_971),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_954),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_990),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_SL g1000 ( 
.A(n_958),
.B(n_222),
.C(n_221),
.Y(n_1000)
);

OR2x6_ASAP7_75t_SL g1001 ( 
.A(n_944),
.B(n_639),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_R g1002 ( 
.A(n_984),
.B(n_0),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_964),
.B(n_641),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_942),
.B(n_0),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_950),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_963),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_971),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_940),
.B(n_1),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_SL g1009 ( 
.A1(n_969),
.A2(n_500),
.B1(n_641),
.B2(n_3),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_939),
.B(n_1),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_938),
.Y(n_1011)
);

CKINVDCx6p67_ASAP7_75t_R g1012 ( 
.A(n_971),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_948),
.B(n_2),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_999),
.A2(n_989),
.B(n_943),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1011),
.B(n_960),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1013),
.B(n_962),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1002),
.A2(n_952),
.B1(n_1009),
.B2(n_955),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_996),
.B(n_946),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_1004),
.A2(n_953),
.B(n_951),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_996),
.A2(n_959),
.B(n_994),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1006),
.B(n_991),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1008),
.B(n_968),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1010),
.A2(n_966),
.B(n_959),
.C(n_947),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_996),
.A2(n_971),
.B1(n_967),
.B2(n_1012),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_997),
.A2(n_957),
.B(n_956),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_997),
.A2(n_995),
.B(n_972),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_1012),
.B(n_945),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_998),
.B(n_965),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1002),
.A2(n_978),
.B1(n_992),
.B2(n_974),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_997),
.A2(n_974),
.B(n_973),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_L g1031 ( 
.A(n_1007),
.B(n_982),
.C(n_985),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1007),
.A2(n_983),
.B1(n_993),
.B2(n_975),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_998),
.B(n_954),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_998),
.B(n_954),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1007),
.A2(n_973),
.B(n_980),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1005),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_1000),
.A2(n_981),
.B(n_986),
.C(n_998),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_1005),
.A2(n_988),
.B(n_987),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_1017),
.A2(n_1023),
.B(n_1025),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1016),
.B(n_1003),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_1014),
.A2(n_979),
.B(n_981),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1027),
.B(n_1033),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_1018),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1021),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_1001),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_1043),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_1043),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_1040),
.B(n_1015),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1047),
.A2(n_1039),
.B(n_1028),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_1048),
.A2(n_1026),
.B(n_1030),
.C(n_1044),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1046),
.B(n_1044),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_1049),
.A2(n_1041),
.B(n_1042),
.Y(n_1052)
);

AO21x2_ASAP7_75t_L g1053 ( 
.A1(n_1051),
.A2(n_1041),
.B(n_1019),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_1053),
.Y(n_1054)
);

INVx8_ASAP7_75t_L g1055 ( 
.A(n_1052),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1055),
.A2(n_1053),
.B1(n_1046),
.B2(n_1042),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_1054),
.A2(n_1052),
.B(n_1036),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1056),
.B(n_1055),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1057),
.B(n_1045),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_1022),
.B1(n_1029),
.B2(n_1024),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_1059),
.A2(n_1053),
.B1(n_1045),
.B2(n_1031),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_1061),
.B(n_1035),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_1060),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1063),
.B(n_1020),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1062),
.B(n_1031),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_SL g1066 ( 
.A(n_1063),
.B(n_1050),
.C(n_1037),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1064),
.B(n_1032),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1065),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1066),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1067),
.B(n_1038),
.Y(n_1070)
);

AND2x4_ASAP7_75t_SL g1071 ( 
.A(n_1068),
.B(n_961),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1071),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1070),
.A2(n_1069),
.B1(n_961),
.B2(n_970),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1072),
.A2(n_961),
.B1(n_976),
.B2(n_949),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1073),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_977),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_1076),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_2),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1078),
.B(n_1001),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1079),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1081),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1080),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_1081),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1084),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1082),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1083),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1087),
.B(n_3),
.Y(n_1088)
);

AOI221xp5_ASAP7_75t_L g1089 ( 
.A1(n_1086),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1089),
.B(n_1085),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1088),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1090),
.B(n_4),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1091),
.B(n_8),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1092),
.A2(n_1093),
.B1(n_9),
.B2(n_10),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1095),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1094),
.A2(n_277),
.B(n_270),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_8),
.Y(n_1098)
);

AOI222xp33_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1099),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1098),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1100),
.A2(n_1102),
.B1(n_1101),
.B2(n_13),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1102),
.B(n_11),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1102),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1105),
.B(n_12),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1103),
.Y(n_1107)
);

XOR2xp5_ASAP7_75t_L g1108 ( 
.A(n_1107),
.B(n_1104),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1106),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1109)
);

NOR4xp75_ASAP7_75t_L g1110 ( 
.A(n_1108),
.B(n_1109),
.C(n_16),
.D(n_17),
.Y(n_1110)
);

NAND4xp25_ASAP7_75t_L g1111 ( 
.A(n_1108),
.B(n_15),
.C(n_17),
.D(n_18),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1110),
.A2(n_19),
.B(n_20),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1113),
.B(n_19),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1112),
.B(n_20),
.Y(n_1115)
);

OR3x1_ASAP7_75t_L g1116 ( 
.A(n_1115),
.B(n_21),
.C(n_22),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_L g1117 ( 
.A(n_1114),
.B(n_22),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1117),
.Y(n_1118)
);

AOI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1116),
.A2(n_277),
.B(n_24),
.C(n_26),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_277),
.B(n_23),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1118),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1120),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1119),
.A2(n_277),
.B1(n_26),
.B2(n_27),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_1121),
.B(n_24),
.C(n_28),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_SL g1125 ( 
.A(n_1122),
.B(n_28),
.C(n_29),
.Y(n_1125)
);

NAND4xp25_ASAP7_75t_SL g1126 ( 
.A(n_1124),
.B(n_1123),
.C(n_1125),
.D(n_31),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1125),
.A2(n_277),
.B1(n_30),
.B2(n_31),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1127),
.B(n_29),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1126),
.B(n_32),
.Y(n_1129)
);

AOI31xp33_ASAP7_75t_L g1130 ( 
.A1(n_1128),
.A2(n_32),
.A3(n_33),
.B(n_34),
.Y(n_1130)
);

OA22x2_ASAP7_75t_L g1131 ( 
.A1(n_1129),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1131),
.B(n_1130),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_1131),
.Y(n_1133)
);

AOI322xp5_ASAP7_75t_L g1134 ( 
.A1(n_1133),
.A2(n_36),
.A3(n_37),
.B1(n_39),
.B2(n_40),
.C1(n_41),
.C2(n_46),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1132),
.Y(n_1135)
);

OA22x2_ASAP7_75t_L g1136 ( 
.A1(n_1135),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1134),
.B(n_41),
.C(n_48),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_49),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1137),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

OAI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1136),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_1141)
);

AOI322xp5_ASAP7_75t_L g1142 ( 
.A1(n_1140),
.A2(n_53),
.A3(n_54),
.B1(n_58),
.B2(n_59),
.C1(n_60),
.C2(n_62),
.Y(n_1142)
);

OAI322xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1139),
.A2(n_64),
.A3(n_66),
.B1(n_68),
.B2(n_70),
.C1(n_72),
.C2(n_73),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1143),
.Y(n_1144)
);

AO22x1_ASAP7_75t_L g1145 ( 
.A1(n_1142),
.A2(n_1141),
.B1(n_75),
.B2(n_77),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1144),
.A2(n_503),
.B1(n_489),
.B2(n_413),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1145),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1147),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1146),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1148),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1149),
.Y(n_1151)
);

XNOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1150),
.B(n_74),
.Y(n_1152)
);

OR3x1_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_78),
.C(n_80),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_81),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1153),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1152),
.B(n_84),
.Y(n_1156)
);

OAI22x1_ASAP7_75t_L g1157 ( 
.A1(n_1153),
.A2(n_503),
.B1(n_489),
.B2(n_87),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1155),
.A2(n_503),
.B(n_489),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1154),
.A2(n_503),
.B(n_429),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1157),
.A2(n_85),
.B(n_86),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1156),
.A2(n_429),
.B(n_408),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1160),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1159),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1158),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1163),
.A2(n_1161),
.B(n_92),
.Y(n_1165)
);

AOI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1164),
.A2(n_91),
.B(n_93),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1162),
.A2(n_94),
.B(n_95),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1164),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1162),
.A2(n_518),
.B1(n_97),
.B2(n_99),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1164),
.A2(n_518),
.B1(n_413),
.B2(n_101),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1164),
.A2(n_518),
.B1(n_413),
.B2(n_102),
.Y(n_1171)
);

AOI22x1_ASAP7_75t_L g1172 ( 
.A1(n_1162),
.A2(n_96),
.B1(n_100),
.B2(n_104),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1164),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_1173)
);

INVx3_ASAP7_75t_SL g1174 ( 
.A(n_1164),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1164),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1164),
.A2(n_110),
.B(n_111),
.Y(n_1176)
);

OR5x1_ASAP7_75t_L g1177 ( 
.A(n_1174),
.B(n_112),
.C(n_114),
.D(n_115),
.E(n_116),
.Y(n_1177)
);

OAI322xp33_ASAP7_75t_L g1178 ( 
.A1(n_1175),
.A2(n_1168),
.A3(n_1165),
.B1(n_1169),
.B2(n_1171),
.C1(n_1170),
.C2(n_1172),
.Y(n_1178)
);

NOR3xp33_ASAP7_75t_SL g1179 ( 
.A(n_1176),
.B(n_1167),
.C(n_1173),
.Y(n_1179)
);

XOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1166),
.B(n_119),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1175),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_1175),
.B(n_120),
.C(n_121),
.Y(n_1182)
);

XNOR2xp5_ASAP7_75t_L g1183 ( 
.A(n_1175),
.B(n_122),
.Y(n_1183)
);

XNOR2xp5_ASAP7_75t_L g1184 ( 
.A(n_1175),
.B(n_125),
.Y(n_1184)
);

XNOR2xp5_ASAP7_75t_L g1185 ( 
.A(n_1175),
.B(n_126),
.Y(n_1185)
);

OAI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1181),
.A2(n_127),
.B(n_128),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1179),
.A2(n_1178),
.B1(n_1180),
.B2(n_1177),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1182),
.A2(n_129),
.B(n_131),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1183),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1184),
.B(n_135),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1185),
.A2(n_137),
.B(n_138),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1181),
.B(n_142),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1187),
.A2(n_143),
.B(n_144),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1190),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1188),
.A2(n_146),
.B(n_147),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1194),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1196),
.A2(n_1195),
.B(n_1192),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1197),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1198),
.A2(n_1191),
.B1(n_1189),
.B2(n_1193),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1199),
.A2(n_1186),
.B(n_150),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1200),
.A2(n_148),
.B1(n_154),
.B2(n_155),
.C(n_156),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1201),
.A2(n_157),
.B(n_158),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1202),
.A2(n_159),
.B1(n_162),
.B2(n_164),
.Y(n_1203)
);

AOI211xp5_ASAP7_75t_L g1204 ( 
.A1(n_1203),
.A2(n_165),
.B(n_166),
.C(n_167),
.Y(n_1204)
);

AOI211xp5_ASAP7_75t_L g1205 ( 
.A1(n_1204),
.A2(n_168),
.B(n_169),
.C(n_170),
.Y(n_1205)
);


endmodule