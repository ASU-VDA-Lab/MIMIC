module fake_aes_3995_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
OR2x6_ASAP7_75t_L g11 ( .A(n_10), .B(n_3), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_9), .B(n_4), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_7), .B1(n_2), .B2(n_6), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
BUFx12f_ASAP7_75t_SL g16 ( .A(n_11), .Y(n_16) );
A2O1A1Ixp33_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_0), .B(n_1), .C(n_2), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
OAI21xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_12), .B(n_15), .Y(n_19) );
OAI22xp5_ASAP7_75t_SL g20 ( .A1(n_18), .A2(n_13), .B1(n_11), .B2(n_14), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_19), .B(n_17), .Y(n_21) );
NAND3xp33_ASAP7_75t_L g22 ( .A(n_20), .B(n_11), .C(n_14), .Y(n_22) );
AO22x1_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_16), .B1(n_11), .B2(n_14), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OAI211xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_14), .B(n_16), .C(n_0), .Y(n_25) );
OAI221xp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_14), .B1(n_0), .B2(n_4), .C(n_5), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
OAI21xp33_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_1), .B(n_5), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_27), .B(n_6), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_27), .B(n_7), .Y(n_32) );
CKINVDCx16_ASAP7_75t_R g33 ( .A(n_31), .Y(n_33) );
OAI21xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_28), .B(n_8), .Y(n_34) );
BUFx2_ASAP7_75t_SL g35 ( .A(n_33), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_34), .B1(n_30), .B2(n_9), .Y(n_36) );
endmodule