module real_aes_18416_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_0), .A2(n_72), .B1(n_807), .B2(n_813), .Y(n_812) );
INVxp33_ASAP7_75t_SL g853 ( .A(n_0), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_1), .A2(n_5), .B1(n_1187), .B2(n_1190), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_2), .A2(n_83), .B1(n_685), .B2(n_711), .Y(n_1025) );
OAI22xp33_ASAP7_75t_SL g1045 ( .A1(n_2), .A2(n_244), .B1(n_662), .B2(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g909 ( .A(n_3), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g1413 ( .A1(n_4), .A2(n_191), .B1(n_783), .B2(n_831), .C(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1440 ( .A(n_4), .Y(n_1440) );
INVx1_ASAP7_75t_L g1415 ( .A(n_6), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g1442 ( .A1(n_6), .A2(n_140), .B1(n_498), .B2(n_1043), .C(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1128 ( .A(n_7), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_7), .A2(n_111), .B1(n_491), .B2(n_674), .Y(n_1149) );
INVx1_ASAP7_75t_L g1367 ( .A(n_8), .Y(n_1367) );
OAI22xp33_ASAP7_75t_L g1397 ( .A1(n_8), .A2(n_121), .B1(n_1020), .B2(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g1017 ( .A(n_9), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_10), .A2(n_204), .B1(n_277), .B2(n_457), .C(n_707), .Y(n_1119) );
OA222x2_ASAP7_75t_L g1151 ( .A1(n_10), .A2(n_49), .B1(n_208), .B2(n_838), .C1(n_841), .C2(n_1083), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_11), .A2(n_20), .B1(n_585), .B2(n_589), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_11), .A2(n_20), .B1(n_622), .B2(n_625), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_12), .A2(n_178), .B1(n_783), .B2(n_966), .C(n_967), .Y(n_965) );
INVx1_ASAP7_75t_L g992 ( .A(n_12), .Y(n_992) );
AND2x2_ASAP7_75t_L g357 ( .A(n_13), .B(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_13), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g402 ( .A(n_13), .Y(n_402) );
AND2x2_ASAP7_75t_L g410 ( .A(n_13), .B(n_210), .Y(n_410) );
INVx1_ASAP7_75t_L g540 ( .A(n_14), .Y(n_540) );
INVx1_ASAP7_75t_L g460 ( .A(n_15), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_15), .A2(n_32), .B1(n_489), .B2(n_490), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g1369 ( .A1(n_16), .A2(n_235), .B1(n_1028), .B2(n_1370), .C(n_1372), .Y(n_1369) );
INVx1_ASAP7_75t_L g1395 ( .A(n_16), .Y(n_1395) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_17), .A2(n_118), .B1(n_328), .B2(n_447), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_17), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_18), .B(n_106), .Y(n_1174) );
INVx2_ASAP7_75t_L g1185 ( .A(n_18), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_18), .B(n_1189), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1381 ( .A1(n_19), .A2(n_199), .B1(n_685), .B2(n_711), .Y(n_1381) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_21), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_21), .A2(n_157), .B1(n_726), .B2(n_727), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_22), .A2(n_215), .B1(n_1187), .B2(n_1190), .Y(n_1193) );
INVx1_ASAP7_75t_L g1069 ( .A(n_23), .Y(n_1069) );
INVx1_ASAP7_75t_L g335 ( .A(n_24), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_25), .A2(n_81), .B1(n_299), .B2(n_816), .C(n_817), .Y(n_815) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_25), .A2(n_26), .B1(n_494), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_26), .A2(n_128), .B1(n_804), .B2(n_807), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g1076 ( .A1(n_27), .A2(n_163), .B1(n_200), .B2(n_305), .C1(n_325), .C2(n_466), .Y(n_1076) );
INVx1_ASAP7_75t_L g1103 ( .A(n_27), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_28), .Y(n_756) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_29), .B(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_30), .A2(n_241), .B1(n_1183), .B2(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g820 ( .A(n_31), .Y(n_820) );
OA222x2_ASAP7_75t_L g837 ( .A1(n_31), .A2(n_153), .B1(n_246), .B2(n_838), .C1(n_840), .C2(n_841), .Y(n_837) );
INVx1_ASAP7_75t_L g476 ( .A(n_32), .Y(n_476) );
OAI22xp5_ASAP7_75t_SL g993 ( .A1(n_33), .A2(n_994), .B1(n_995), .B2(n_1048), .Y(n_993) );
INVx1_ASAP7_75t_L g1048 ( .A(n_33), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_33), .A2(n_994), .B1(n_995), .B2(n_1048), .Y(n_1050) );
INVx1_ASAP7_75t_L g472 ( .A(n_34), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_34), .A2(n_161), .B1(n_489), .B2(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g1416 ( .A(n_35), .Y(n_1416) );
AOI221xp5_ASAP7_75t_L g1436 ( .A1(n_35), .A2(n_80), .B1(n_1376), .B2(n_1437), .C(n_1439), .Y(n_1436) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_36), .A2(n_190), .B1(n_321), .B2(n_809), .C(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g858 ( .A(n_36), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_37), .A2(n_239), .B1(n_886), .B2(n_887), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_37), .A2(n_239), .B1(n_937), .B2(n_939), .Y(n_936) );
AOI211xp5_ASAP7_75t_L g957 ( .A1(n_38), .A2(n_816), .B(n_958), .C(n_960), .Y(n_957) );
INVx1_ASAP7_75t_L g988 ( .A(n_38), .Y(n_988) );
INVx1_ASAP7_75t_L g507 ( .A(n_39), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g1425 ( .A1(n_40), .A2(n_66), .B1(n_274), .B2(n_279), .C(n_285), .Y(n_1425) );
INVxp67_ASAP7_75t_SL g1432 ( .A(n_40), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_41), .A2(n_222), .B1(n_1187), .B2(n_1190), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1363 ( .A1(n_42), .A2(n_129), .B1(n_668), .B2(n_848), .C(n_1364), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_42), .A2(n_90), .B1(n_806), .B2(n_1393), .Y(n_1392) );
AO22x1_ASAP7_75t_L g1182 ( .A1(n_43), .A2(n_61), .B1(n_1172), .B2(n_1183), .Y(n_1182) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_44), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_44), .A2(n_48), .B1(n_297), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_45), .A2(n_155), .B1(n_430), .B2(n_674), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_45), .A2(n_107), .B1(n_720), .B2(n_783), .Y(n_1389) );
INVx1_ASAP7_75t_L g912 ( .A(n_46), .Y(n_912) );
INVx1_ASAP7_75t_L g267 ( .A(n_47), .Y(n_267) );
INVx1_ASAP7_75t_L g284 ( .A(n_47), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_48), .A2(n_157), .B1(n_667), .B2(n_668), .C(n_672), .Y(n_666) );
INVx1_ASAP7_75t_L g1118 ( .A(n_49), .Y(n_1118) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_50), .A2(n_227), .B1(n_274), .B2(n_279), .C(n_285), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_50), .A2(n_123), .B1(n_407), .B2(n_486), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_51), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_52), .Y(n_761) );
INVx1_ASAP7_75t_L g314 ( .A(n_53), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g1000 ( .A1(n_54), .A2(n_156), .B1(n_728), .B2(n_1001), .C(n_1003), .Y(n_1000) );
OAI211xp5_ASAP7_75t_L g1027 ( .A1(n_54), .A2(n_1028), .B(n_1029), .C(n_1034), .Y(n_1027) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_55), .A2(n_108), .B1(n_328), .B2(n_447), .C(n_448), .Y(n_446) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_55), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_56), .A2(n_148), .B1(n_1062), .B2(n_1064), .C(n_1066), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_56), .A2(n_206), .B1(n_1099), .B2(n_1101), .C(n_1102), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1405 ( .A1(n_57), .A2(n_1406), .B1(n_1407), .B2(n_1408), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1406 ( .A(n_57), .Y(n_1406) );
INVx1_ASAP7_75t_L g577 ( .A(n_58), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g1058 ( .A1(n_59), .A2(n_226), .B1(n_274), .B2(n_279), .C(n_285), .Y(n_1058) );
OAI21xp33_ASAP7_75t_SL g1089 ( .A1(n_59), .A2(n_418), .B(n_841), .Y(n_1089) );
INVx1_ASAP7_75t_L g1163 ( .A(n_60), .Y(n_1163) );
INVx2_ASAP7_75t_L g270 ( .A(n_62), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g1424 ( .A1(n_63), .A2(n_197), .B1(n_328), .B2(n_447), .Y(n_1424) );
INVx1_ASAP7_75t_L g1435 ( .A(n_63), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_64), .A2(n_173), .B1(n_337), .B2(n_340), .Y(n_1412) );
INVx1_ASAP7_75t_L g1433 ( .A(n_64), .Y(n_1433) );
INVx1_ASAP7_75t_L g904 ( .A(n_65), .Y(n_904) );
INVx1_ASAP7_75t_L g1449 ( .A(n_66), .Y(n_1449) );
INVx1_ASAP7_75t_L g522 ( .A(n_67), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g319 ( .A1(n_68), .A2(n_320), .B(n_321), .Y(n_319) );
INVxp67_ASAP7_75t_L g384 ( .A(n_68), .Y(n_384) );
INVx1_ASAP7_75t_L g518 ( .A(n_69), .Y(n_518) );
INVx1_ASAP7_75t_L g531 ( .A(n_70), .Y(n_531) );
INVx1_ASAP7_75t_L g766 ( .A(n_71), .Y(n_766) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_72), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g1070 ( .A1(n_73), .A2(n_74), .B1(n_337), .B2(n_340), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1081 ( .A(n_73), .Y(n_1081) );
INVx1_ASAP7_75t_L g1087 ( .A(n_74), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_75), .A2(n_165), .B1(n_1172), .B2(n_1183), .Y(n_1204) );
AO221x2_ASAP7_75t_L g1230 ( .A1(n_76), .A2(n_202), .B1(n_1187), .B2(n_1190), .C(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1380 ( .A(n_77), .Y(n_1380) );
OAI211xp5_ASAP7_75t_L g571 ( .A1(n_78), .A2(n_393), .B(n_572), .C(n_576), .Y(n_571) );
INVx1_ASAP7_75t_L g620 ( .A(n_78), .Y(n_620) );
INVx1_ASAP7_75t_L g1057 ( .A(n_79), .Y(n_1057) );
OAI21xp33_ASAP7_75t_L g1082 ( .A1(n_79), .A2(n_1083), .B(n_1084), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1417 ( .A1(n_80), .A2(n_192), .B1(n_783), .B2(n_1418), .C(n_1419), .Y(n_1417) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_81), .A2(n_190), .B1(n_847), .B2(n_848), .C(n_849), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g1123 ( .A(n_82), .Y(n_1123) );
INVx1_ASAP7_75t_L g1130 ( .A(n_84), .Y(n_1130) );
AOI221x1_ASAP7_75t_SL g1144 ( .A1(n_84), .A2(n_101), .B1(n_430), .B2(n_668), .C(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g905 ( .A(n_85), .Y(n_905) );
OAI222xp33_ASAP7_75t_L g772 ( .A1(n_86), .A2(n_122), .B1(n_220), .B2(n_332), .C1(n_773), .C2(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g795 ( .A(n_86), .Y(n_795) );
INVx1_ASAP7_75t_L g524 ( .A(n_87), .Y(n_524) );
INVx1_ASAP7_75t_L g830 ( .A(n_88), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_88), .B(n_350), .Y(n_835) );
INVx1_ASAP7_75t_L g474 ( .A(n_89), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_89), .A2(n_211), .B1(n_430), .B2(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_SL g1374 ( .A(n_90), .Y(n_1374) );
XOR2x2_ASAP7_75t_L g949 ( .A(n_91), .B(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g897 ( .A(n_92), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_93), .Y(n_454) );
INVx1_ASAP7_75t_L g682 ( .A(n_94), .Y(n_682) );
INVx1_ASAP7_75t_L g1115 ( .A(n_95), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_95), .A2(n_204), .B1(n_405), .B2(n_414), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_96), .A2(n_168), .B1(n_337), .B2(n_340), .Y(n_336) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_96), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_97), .A2(n_123), .B1(n_337), .B2(n_340), .Y(n_964) );
OAI211xp5_ASAP7_75t_L g971 ( .A1(n_97), .A2(n_350), .B(n_972), .C(n_975), .Y(n_971) );
INVx1_ASAP7_75t_L g760 ( .A(n_98), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_98), .A2(n_139), .B1(n_781), .B2(n_783), .C(n_784), .Y(n_780) );
INVx1_ASAP7_75t_L g832 ( .A(n_99), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_99), .A2(n_169), .B1(n_407), .B2(n_486), .Y(n_865) );
INVx1_ASAP7_75t_L g963 ( .A(n_100), .Y(n_963) );
INVx1_ASAP7_75t_L g1139 ( .A(n_101), .Y(n_1139) );
INVx1_ASAP7_75t_L g533 ( .A(n_102), .Y(n_533) );
OA22x2_ASAP7_75t_L g869 ( .A1(n_103), .A2(n_870), .B1(n_943), .B2(n_944), .Y(n_869) );
INVxp67_ASAP7_75t_L g944 ( .A(n_103), .Y(n_944) );
INVx1_ASAP7_75t_L g969 ( .A(n_104), .Y(n_969) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_105), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_105), .B(n_1163), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_106), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1189 ( .A(n_106), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_107), .A2(n_146), .B1(n_670), .B2(n_1044), .C(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g506 ( .A(n_108), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_109), .Y(n_698) );
INVx1_ASAP7_75t_L g968 ( .A(n_110), .Y(n_968) );
INVx1_ASAP7_75t_L g1134 ( .A(n_111), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_112), .A2(n_240), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_112), .A2(n_144), .B1(n_720), .B2(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g892 ( .A(n_113), .Y(n_892) );
INVx2_ASAP7_75t_L g272 ( .A(n_114), .Y(n_272) );
INVx1_ASAP7_75t_L g302 ( .A(n_114), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_114), .B(n_270), .Y(n_331) );
INVx1_ASAP7_75t_L g316 ( .A(n_115), .Y(n_316) );
INVx1_ASAP7_75t_L g767 ( .A(n_116), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_116), .A2(n_145), .B1(n_274), .B2(n_279), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g874 ( .A1(n_117), .A2(n_171), .B1(n_875), .B2(n_877), .Y(n_874) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_117), .A2(n_171), .B1(n_595), .B2(n_942), .Y(n_941) );
INVxp67_ASAP7_75t_SL g1078 ( .A(n_118), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_119), .A2(n_198), .B1(n_1172), .B2(n_1183), .Y(n_1228) );
XOR2xp5_ASAP7_75t_L g1106 ( .A(n_120), .B(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1368 ( .A(n_121), .Y(n_1368) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_122), .A2(n_145), .B1(n_405), .B2(n_414), .C(n_418), .Y(n_763) );
INVx1_ASAP7_75t_L g736 ( .A(n_124), .Y(n_736) );
INVx1_ASAP7_75t_L g477 ( .A(n_125), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_125), .A2(n_172), .B1(n_503), .B2(n_505), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g1132 ( .A(n_126), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_127), .A2(n_164), .B1(n_593), .B2(n_597), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_127), .A2(n_164), .B1(n_605), .B2(n_606), .Y(n_604) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_128), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_129), .A2(n_158), .B1(n_804), .B2(n_809), .Y(n_1385) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_130), .A2(n_136), .B1(n_473), .B2(n_811), .Y(n_1116) );
INVx1_ASAP7_75t_L g1154 ( .A(n_130), .Y(n_1154) );
INVx1_ASAP7_75t_L g1423 ( .A(n_131), .Y(n_1423) );
INVx1_ASAP7_75t_L g527 ( .A(n_132), .Y(n_527) );
INVx1_ASAP7_75t_L g902 ( .A(n_133), .Y(n_902) );
XOR2x2_ASAP7_75t_L g255 ( .A(n_134), .B(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_135), .A2(n_138), .B1(n_328), .B2(n_447), .Y(n_955) );
INVxp67_ASAP7_75t_SL g976 ( .A(n_135), .Y(n_976) );
INVx1_ASAP7_75t_L g1153 ( .A(n_136), .Y(n_1153) );
AO22x1_ASAP7_75t_L g1186 ( .A1(n_137), .A2(n_213), .B1(n_1187), .B2(n_1190), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g973 ( .A(n_138), .Y(n_973) );
INVx1_ASAP7_75t_L g742 ( .A(n_139), .Y(n_742) );
INVx1_ASAP7_75t_L g1420 ( .A(n_140), .Y(n_1420) );
INVx1_ASAP7_75t_L g645 ( .A(n_141), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_141), .A2(n_240), .B1(n_722), .B2(n_724), .Y(n_723) );
BUFx3_ASAP7_75t_L g264 ( .A(n_142), .Y(n_264) );
INVx1_ASAP7_75t_L g1011 ( .A(n_143), .Y(n_1011) );
INVx1_ASAP7_75t_L g647 ( .A(n_144), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_146), .A2(n_155), .B1(n_1387), .B2(n_1388), .Y(n_1386) );
INVx1_ASAP7_75t_L g259 ( .A(n_147), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_148), .B(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g959 ( .A(n_149), .Y(n_959) );
INVx1_ASAP7_75t_L g1068 ( .A(n_150), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_151), .A2(n_160), .B1(n_1187), .B2(n_1190), .Y(n_1209) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_152), .Y(n_363) );
INVx1_ASAP7_75t_L g834 ( .A(n_153), .Y(n_834) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_154), .A2(n_685), .B(n_688), .Y(n_684) );
OAI221xp5_ASAP7_75t_SL g1035 ( .A1(n_156), .A2(n_183), .B1(n_657), .B2(n_1036), .C(n_1038), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g1373 ( .A(n_158), .Y(n_1373) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_159), .A2(n_297), .B(n_299), .Y(n_296) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_159), .Y(n_378) );
INVx1_ASAP7_75t_L g458 ( .A(n_161), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_162), .A2(n_230), .B1(n_831), .B2(n_1019), .Y(n_1018) );
INVxp67_ASAP7_75t_SL g1041 ( .A(n_162), .Y(n_1041) );
INVx1_ASAP7_75t_L g1095 ( .A(n_163), .Y(n_1095) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_166), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_167), .A2(n_223), .B1(n_1172), .B2(n_1183), .Y(n_1194) );
AOI222xp33_ASAP7_75t_L g1355 ( .A1(n_167), .A2(n_1356), .B1(n_1401), .B2(n_1404), .C1(n_1450), .C2(n_1452), .Y(n_1355) );
XOR2x2_ASAP7_75t_L g1357 ( .A(n_167), .B(n_1358), .Y(n_1357) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_168), .A2(n_193), .B1(n_405), .B2(n_414), .C(n_418), .Y(n_404) );
INVx1_ASAP7_75t_L g819 ( .A(n_169), .Y(n_819) );
OAI211xp5_ASAP7_75t_SL g878 ( .A1(n_170), .A2(n_610), .B(n_879), .C(n_881), .Y(n_878) );
INVx1_ASAP7_75t_L g933 ( .A(n_170), .Y(n_933) );
INVx1_ASAP7_75t_L g468 ( .A(n_172), .Y(n_468) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_173), .Y(n_1447) );
INVx1_ASAP7_75t_L g883 ( .A(n_174), .Y(n_883) );
INVx1_ASAP7_75t_L g333 ( .A(n_175), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_176), .A2(n_219), .B1(n_1172), .B2(n_1183), .Y(n_1208) );
INVxp67_ASAP7_75t_SL g1006 ( .A(n_177), .Y(n_1006) );
AOI221xp5_ASAP7_75t_L g1042 ( .A1(n_177), .A2(n_218), .B1(n_1031), .B2(n_1043), .C(n_1044), .Y(n_1042) );
INVx1_ASAP7_75t_L g983 ( .A(n_178), .Y(n_983) );
INVx1_ASAP7_75t_L g308 ( .A(n_179), .Y(n_308) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_180), .Y(n_361) );
OAI222xp33_ASAP7_75t_L g637 ( .A1(n_181), .A2(n_238), .B1(n_638), .B2(n_642), .C1(n_651), .C2(n_657), .Y(n_637) );
INVx1_ASAP7_75t_L g701 ( .A(n_181), .Y(n_701) );
INVx1_ASAP7_75t_L g450 ( .A(n_182), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_182), .A2(n_184), .B1(n_407), .B2(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_SL g997 ( .A(n_183), .Y(n_997) );
INVx1_ASAP7_75t_L g453 ( .A(n_184), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g1126 ( .A(n_185), .Y(n_1126) );
INVx1_ASAP7_75t_L g961 ( .A(n_186), .Y(n_961) );
INVx1_ASAP7_75t_L g884 ( .A(n_187), .Y(n_884) );
OAI211xp5_ASAP7_75t_SL g929 ( .A1(n_187), .A2(n_572), .B(n_930), .C(n_931), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_188), .Y(n_751) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_189), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_189), .A2(n_447), .B1(n_788), .B2(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g1444 ( .A(n_191), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_192), .Y(n_1445) );
OAI221xp5_ASAP7_75t_L g273 ( .A1(n_193), .A2(n_216), .B1(n_274), .B2(n_279), .C(n_285), .Y(n_273) );
AO22x1_ASAP7_75t_L g1224 ( .A1(n_194), .A2(n_214), .B1(n_1183), .B2(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g679 ( .A(n_195), .Y(n_679) );
CKINVDCx16_ASAP7_75t_R g1232 ( .A(n_196), .Y(n_1232) );
INVxp67_ASAP7_75t_SL g1427 ( .A(n_197), .Y(n_1427) );
OAI211xp5_ASAP7_75t_L g1360 ( .A1(n_199), .A2(n_1361), .B(n_1362), .C(n_1366), .Y(n_1360) );
AOI21xp33_ASAP7_75t_L g1096 ( .A1(n_200), .A2(n_545), .B(n_667), .Y(n_1096) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_201), .A2(n_261), .B(n_285), .C(n_452), .Y(n_451) );
INVxp33_ASAP7_75t_SL g484 ( .A(n_201), .Y(n_484) );
INVx1_ASAP7_75t_L g953 ( .A(n_203), .Y(n_953) );
INVx1_ASAP7_75t_L g1012 ( .A(n_205), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_205), .A2(n_230), .B1(n_489), .B2(n_1031), .C(n_1033), .Y(n_1030) );
AOI21xp33_ASAP7_75t_L g1071 ( .A1(n_206), .A2(n_1072), .B(n_1075), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_207), .Y(n_744) );
INVx1_ASAP7_75t_L g1112 ( .A(n_208), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_209), .A2(n_229), .B1(n_1187), .B2(n_1190), .Y(n_1198) );
INVx1_ASAP7_75t_L g358 ( .A(n_210), .Y(n_358) );
BUFx3_ASAP7_75t_L g371 ( .A(n_210), .Y(n_371) );
INVx1_ASAP7_75t_L g464 ( .A(n_211), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g1234 ( .A(n_212), .Y(n_1234) );
INVx1_ASAP7_75t_L g866 ( .A(n_213), .Y(n_866) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_216), .Y(n_435) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_217), .A2(n_662), .B(n_665), .C(n_677), .Y(n_661) );
INVx1_ASAP7_75t_L g709 ( .A(n_217), .Y(n_709) );
INVx1_ASAP7_75t_L g1014 ( .A(n_218), .Y(n_1014) );
INVx1_ASAP7_75t_L g769 ( .A(n_220), .Y(n_769) );
INVx2_ASAP7_75t_L g346 ( .A(n_221), .Y(n_346) );
INVx1_ASAP7_75t_L g355 ( .A(n_221), .Y(n_355) );
INVx1_ASAP7_75t_L g424 ( .A(n_221), .Y(n_424) );
XOR2x2_ASAP7_75t_L g511 ( .A(n_222), .B(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_224), .A2(n_233), .B1(n_324), .B2(n_325), .Y(n_323) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_224), .Y(n_398) );
INVx1_ASAP7_75t_L g1421 ( .A(n_225), .Y(n_1421) );
INVx1_ASAP7_75t_L g1085 ( .A(n_226), .Y(n_1085) );
INVxp67_ASAP7_75t_SL g974 ( .A(n_227), .Y(n_974) );
AO22x1_ASAP7_75t_L g1226 ( .A1(n_228), .A2(n_242), .B1(n_1187), .B2(n_1190), .Y(n_1226) );
XOR2x2_ASAP7_75t_L g1053 ( .A(n_229), .B(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1024 ( .A(n_231), .Y(n_1024) );
INVx1_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_233), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g1136 ( .A(n_234), .Y(n_1136) );
INVx1_ASAP7_75t_L g1396 ( .A(n_235), .Y(n_1396) );
OAI21xp33_ASAP7_75t_SL g444 ( .A1(n_236), .A2(n_350), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g449 ( .A(n_236), .Y(n_449) );
INVx1_ASAP7_75t_L g543 ( .A(n_237), .Y(n_543) );
INVx1_ASAP7_75t_L g704 ( .A(n_238), .Y(n_704) );
INVx1_ASAP7_75t_L g1009 ( .A(n_243), .Y(n_1009) );
OAI322xp33_ASAP7_75t_SL g1004 ( .A1(n_244), .A2(n_534), .A3(n_914), .B1(n_1005), .B2(n_1010), .C1(n_1013), .C2(n_1020), .Y(n_1004) );
INVx1_ASAP7_75t_L g580 ( .A(n_245), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g609 ( .A1(n_245), .A2(n_541), .B(n_610), .C(n_612), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g824 ( .A1(n_246), .A2(n_248), .B1(n_825), .B2(n_826), .C(n_829), .Y(n_824) );
INVx1_ASAP7_75t_L g900 ( .A(n_247), .Y(n_900) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_248), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_1157), .B(n_1169), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_731), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g1157 ( .A1(n_252), .A2(n_1158), .B(n_1159), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_508), .B1(n_509), .B2(n_730), .Y(n_252) );
INVx1_ASAP7_75t_L g730 ( .A(n_253), .Y(n_730) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_442), .Y(n_254) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_364), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_326), .B(n_343), .C(n_347), .Y(n_257) );
AOI211xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_273), .C(n_290), .Y(n_258) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_259), .A2(n_335), .B1(n_421), .B2(n_427), .C1(n_433), .C2(n_435), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_260), .A2(n_766), .B1(n_772), .B2(n_775), .C(n_777), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_260), .A2(n_822), .B1(n_824), .B2(n_834), .Y(n_821) );
AOI211xp5_ASAP7_75t_L g952 ( .A1(n_260), .A2(n_953), .B(n_954), .C(n_955), .Y(n_952) );
AOI211xp5_ASAP7_75t_SL g1056 ( .A1(n_260), .A2(n_1057), .B(n_1058), .C(n_1059), .Y(n_1056) );
AOI211xp5_ASAP7_75t_SL g1422 ( .A1(n_260), .A2(n_1423), .B(n_1424), .C(n_1425), .Y(n_1422) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g711 ( .A(n_261), .B(n_712), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_262), .B(n_268), .Y(n_261) );
INVx8_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
BUFx3_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
AND2x2_ASAP7_75t_L g338 ( .A(n_262), .B(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g806 ( .A(n_262), .Y(n_806) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
AND2x4_ASAP7_75t_L g306 ( .A(n_263), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_264), .B(n_284), .Y(n_313) );
AND2x4_ASAP7_75t_L g342 ( .A(n_264), .B(n_283), .Y(n_342) );
OR2x2_ASAP7_75t_L g467 ( .A(n_264), .B(n_266), .Y(n_467) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_L g307 ( .A(n_267), .Y(n_307) );
AND2x6_ASAP7_75t_L g275 ( .A(n_268), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g280 ( .A(n_268), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
AND2x4_ASAP7_75t_L g703 ( .A(n_268), .B(n_423), .Y(n_703) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_269), .B(n_302), .Y(n_301) );
NAND3x1_ASAP7_75t_L g537 ( .A(n_269), .B(n_302), .C(n_538), .Y(n_537) );
OR2x4_ASAP7_75t_L g605 ( .A(n_269), .B(n_467), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_269), .Y(n_608) );
AND2x4_ASAP7_75t_L g611 ( .A(n_269), .B(n_342), .Y(n_611) );
OR2x6_ASAP7_75t_L g626 ( .A(n_269), .B(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp33_ASAP7_75t_SL g322 ( .A(n_270), .B(n_272), .Y(n_322) );
BUFx3_ASAP7_75t_L g462 ( .A(n_270), .Y(n_462) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g461 ( .A(n_272), .B(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_272), .Y(n_631) );
AND3x4_ASAP7_75t_L g715 ( .A(n_272), .B(n_345), .C(n_462), .Y(n_715) );
INVx4_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_275), .A2(n_280), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_275), .A2(n_280), .B1(n_779), .B2(n_819), .C(n_820), .Y(n_818) );
AND2x2_ASAP7_75t_L g702 ( .A(n_276), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_276), .B(n_703), .Y(n_1002) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_278), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g325 ( .A(n_278), .B(n_282), .Y(n_325) );
BUFx2_ASAP7_75t_L g616 ( .A(n_278), .Y(n_616) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g707 ( .A(n_281), .Y(n_707) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g288 ( .A(n_284), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_285), .Y(n_779) );
OR2x6_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx1_ASAP7_75t_L g880 ( .A(n_286), .Y(n_880) );
INVx1_ASAP7_75t_L g1074 ( .A(n_286), .Y(n_1074) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_287), .Y(n_295) );
BUFx3_ASAP7_75t_L g542 ( .A(n_287), .Y(n_542) );
BUFx2_ASAP7_75t_L g619 ( .A(n_288), .Y(n_619) );
INVx1_ASAP7_75t_L g1120 ( .A(n_289), .Y(n_1120) );
OAI21xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_303), .B(n_315), .Y(n_290) );
OAI21xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_296), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_292), .A2(n_316), .B1(n_392), .B2(n_393), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_293), .A2(n_300), .B1(n_472), .B2(n_473), .C(n_474), .Y(n_471) );
OAI221xp5_ASAP7_75t_L g1135 ( .A1(n_293), .A2(n_461), .B1(n_1136), .B2(n_1137), .C(n_1139), .Y(n_1135) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g1065 ( .A(n_294), .Y(n_1065) );
INVx1_ASAP7_75t_L g1129 ( .A(n_294), .Y(n_1129) );
INVx4_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx3_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_295), .Y(n_457) );
OR2x2_ASAP7_75t_L g686 ( .A(n_295), .B(n_687), .Y(n_686) );
INVx8_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g690 ( .A(n_298), .Y(n_690) );
INVx3_ASAP7_75t_L g726 ( .A(n_298), .Y(n_726) );
INVx2_ASAP7_75t_L g831 ( .A(n_298), .Y(n_831) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_300), .A2(n_473), .B1(n_542), .B2(n_744), .C(n_756), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_300), .A2(n_473), .B1(n_542), .B2(n_968), .C(n_969), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_300), .B(n_1076), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_300), .A2(n_773), .B1(n_1128), .B2(n_1129), .C(n_1130), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1419 ( .A1(n_300), .A2(n_521), .B1(n_542), .B2(n_1420), .C(n_1421), .Y(n_1419) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x6_ASAP7_75t_L g1391 ( .A(n_301), .B(n_369), .Y(n_1391) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_308), .B1(n_309), .B2(n_314), .Y(n_303) );
INVx1_ASAP7_75t_L g1418 ( .A(n_304), .Y(n_1418) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g459 ( .A(n_305), .Y(n_459) );
AND2x4_ASAP7_75t_L g692 ( .A(n_305), .B(n_691), .Y(n_692) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_305), .Y(n_724) );
INVx3_ASAP7_75t_L g790 ( .A(n_305), .Y(n_790) );
BUFx8_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_306), .Y(n_320) );
INVx2_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_306), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_308), .A2(n_384), .B1(n_385), .B2(n_388), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_309), .A2(n_459), .B1(n_476), .B2(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g532 ( .A(n_311), .Y(n_532) );
OR2x2_ASAP7_75t_L g696 ( .A(n_311), .B(n_687), .Y(n_696) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_312), .Y(n_470) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g627 ( .A(n_313), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_314), .A2(n_379), .B1(n_396), .B2(n_398), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_319), .C(n_323), .Y(n_315) );
INVx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g774 ( .A(n_318), .Y(n_774) );
INVx5_ASAP7_75t_L g721 ( .A(n_320), .Y(n_721) );
INVx2_ASAP7_75t_SL g811 ( .A(n_320), .Y(n_811) );
INVx2_ASAP7_75t_SL g814 ( .A(n_320), .Y(n_814) );
INVx3_ASAP7_75t_L g825 ( .A(n_320), .Y(n_825) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_320), .Y(n_1125) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g516 ( .A(n_322), .B(n_403), .Y(n_516) );
INVx1_ASAP7_75t_L g782 ( .A(n_324), .Y(n_782) );
BUFx2_ASAP7_75t_L g817 ( .A(n_324), .Y(n_817) );
AND2x4_ASAP7_75t_L g334 ( .A(n_325), .B(n_330), .Y(n_334) );
BUFx3_ASAP7_75t_L g722 ( .A(n_325), .Y(n_722) );
BUFx3_ASAP7_75t_L g783 ( .A(n_325), .Y(n_783) );
BUFx2_ASAP7_75t_L g807 ( .A(n_325), .Y(n_807) );
INVx5_ASAP7_75t_L g1067 ( .A(n_325), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_333), .B1(n_334), .B2(n_335), .C(n_336), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_328), .Y(n_327) );
OR2x6_ASAP7_75t_SL g328 ( .A(n_329), .B(n_332), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_330), .Y(n_776) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g339 ( .A(n_331), .Y(n_339) );
OR2x2_ASAP7_75t_L g687 ( .A(n_331), .B(n_403), .Y(n_687) );
BUFx2_ASAP7_75t_L g530 ( .A(n_332), .Y(n_530) );
INVx3_ASAP7_75t_L g786 ( .A(n_332), .Y(n_786) );
INVx1_ASAP7_75t_L g1008 ( .A(n_332), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_333), .B(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g447 ( .A(n_334), .Y(n_447) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_338), .A2(n_341), .B1(n_449), .B2(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g341 ( .A(n_339), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g718 ( .A(n_342), .Y(n_718) );
BUFx2_ASAP7_75t_L g727 ( .A(n_342), .Y(n_727) );
BUFx2_ASAP7_75t_L g809 ( .A(n_342), .Y(n_809) );
BUFx3_ASAP7_75t_L g816 ( .A(n_342), .Y(n_816) );
BUFx2_ASAP7_75t_L g833 ( .A(n_342), .Y(n_833) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_342), .Y(n_1019) );
INVx2_ASAP7_75t_L g1114 ( .A(n_342), .Y(n_1114) );
INVx1_ASAP7_75t_L g1378 ( .A(n_343), .Y(n_1378) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI31xp33_ASAP7_75t_SL g445 ( .A1(n_345), .A2(n_446), .A3(n_451), .B(n_455), .Y(n_445) );
INVx2_ASAP7_75t_SL g683 ( .A(n_345), .Y(n_683) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g369 ( .A(n_346), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_346), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_351), .B(n_769), .Y(n_768) );
AOI211xp5_ASAP7_75t_L g1080 ( .A1(n_351), .A2(n_1081), .B(n_1082), .C(n_1089), .Y(n_1080) );
AOI22xp33_ASAP7_75t_SL g1152 ( .A1(n_351), .A2(n_437), .B1(n_1153), .B2(n_1154), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_351), .B(n_1447), .Y(n_1446) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .Y(n_351) );
AND2x4_ASAP7_75t_L g437 ( .A(n_352), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g414 ( .A(n_353), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g486 ( .A(n_353), .B(n_415), .Y(n_486) );
INVx1_ASAP7_75t_L g602 ( .A(n_353), .Y(n_602) );
INVxp67_ASAP7_75t_L g712 ( .A(n_353), .Y(n_712) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_356), .Y(n_678) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_357), .B(n_424), .Y(n_429) );
AND2x2_ASAP7_75t_L g438 ( .A(n_357), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_SL g641 ( .A(n_357), .B(n_491), .Y(n_641) );
AND2x4_ASAP7_75t_L g663 ( .A(n_357), .B(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g681 ( .A(n_357), .B(n_439), .Y(n_681) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_358), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_359), .B(n_410), .Y(n_426) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_359), .Y(n_494) );
INVx3_ASAP7_75t_L g504 ( .A(n_359), .Y(n_504) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
OR2x2_ASAP7_75t_L g387 ( .A(n_360), .B(n_363), .Y(n_387) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g377 ( .A(n_361), .B(n_363), .Y(n_377) );
INVx2_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
NAND2x1_ASAP7_75t_L g390 ( .A(n_361), .B(n_363), .Y(n_390) );
INVx1_ASAP7_75t_L g417 ( .A(n_361), .Y(n_417) );
AND2x2_ASAP7_75t_L g440 ( .A(n_361), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g492 ( .A(n_361), .B(n_363), .Y(n_492) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_363), .B(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g413 ( .A(n_363), .Y(n_413) );
AND2x2_ASAP7_75t_L g432 ( .A(n_363), .B(n_382), .Y(n_432) );
INVx2_ASAP7_75t_L g441 ( .A(n_363), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_420), .C(n_436), .Y(n_364) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_404), .Y(n_365) );
OAI33xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_372), .A3(n_383), .B1(n_391), .B2(n_395), .B3(n_399), .Y(n_366) );
OAI33xp33_ASAP7_75t_L g740 ( .A1(n_367), .A2(n_741), .A3(n_746), .B1(n_752), .B2(n_757), .B3(n_762), .Y(n_740) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g496 ( .A(n_368), .Y(n_496) );
INVx2_ASAP7_75t_L g545 ( .A(n_368), .Y(n_545) );
INVx2_ASAP7_75t_L g864 ( .A(n_368), .Y(n_864) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_368), .Y(n_1143) );
AOI222xp33_ASAP7_75t_L g1434 ( .A1(n_368), .A2(n_421), .B1(n_499), .B2(n_1435), .C1(n_1436), .C2(n_1442), .Y(n_1434) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g793 ( .A(n_369), .Y(n_793) );
AND2x4_ASAP7_75t_L g401 ( .A(n_371), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g575 ( .A(n_371), .Y(n_575) );
BUFx2_ASAP7_75t_L g579 ( .A(n_371), .Y(n_579) );
AND2x4_ASAP7_75t_L g583 ( .A(n_371), .B(n_416), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_378), .B2(n_379), .Y(n_372) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g397 ( .A(n_375), .Y(n_397) );
BUFx3_ASAP7_75t_L g549 ( .A(n_375), .Y(n_549) );
BUFx3_ASAP7_75t_L g991 ( .A(n_375), .Y(n_991) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g587 ( .A(n_376), .Y(n_587) );
BUFx4f_ASAP7_75t_L g852 ( .A(n_376), .Y(n_852) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_379), .A2(n_396), .B1(n_1373), .B2(n_1374), .C(n_1375), .Y(n_1372) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx8_ASAP7_75t_L g552 ( .A(n_380), .Y(n_552) );
OR2x2_ASAP7_75t_L g591 ( .A(n_380), .B(n_579), .Y(n_591) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_385), .A2(n_854), .B1(n_1126), .B2(n_1136), .C(n_1149), .Y(n_1148) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g392 ( .A(n_387), .Y(n_392) );
INVx2_ASAP7_75t_L g555 ( .A(n_387), .Y(n_555) );
BUFx3_ASAP7_75t_L g562 ( .A(n_387), .Y(n_562) );
BUFx2_ASAP7_75t_L g750 ( .A(n_387), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_388), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_752) );
BUFx2_ASAP7_75t_L g930 ( .A(n_388), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_388), .A2(n_549), .B1(n_1123), .B2(n_1132), .Y(n_1145) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g434 ( .A(n_389), .B(n_429), .Y(n_434) );
INVx2_ASAP7_75t_SL g644 ( .A(n_389), .Y(n_644) );
OR2x2_ASAP7_75t_L g841 ( .A(n_389), .B(n_429), .Y(n_841) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_390), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_393), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x6_ASAP7_75t_L g418 ( .A(n_394), .B(n_419), .Y(n_418) );
INVx4_ASAP7_75t_L g558 ( .A(n_394), .Y(n_558) );
BUFx4f_ASAP7_75t_L g563 ( .A(n_394), .Y(n_563) );
BUFx4f_ASAP7_75t_L g982 ( .A(n_394), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_396), .A2(n_652), .B1(n_653), .B2(n_656), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_396), .A2(n_568), .B1(n_1009), .B2(n_1017), .C(n_1030), .Y(n_1029) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g762 ( .A(n_400), .Y(n_762) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_401), .B(n_403), .Y(n_400) );
AND2x4_ASAP7_75t_L g499 ( .A(n_401), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_401), .B(n_500), .Y(n_566) );
INVx4_ASAP7_75t_L g672 ( .A(n_401), .Y(n_672) );
INVx4_ASAP7_75t_L g1033 ( .A(n_401), .Y(n_1033) );
INVx1_ASAP7_75t_SL g1364 ( .A(n_401), .Y(n_1364) );
INVx1_ASAP7_75t_L g601 ( .A(n_402), .Y(n_601) );
AND2x4_ASAP7_75t_L g650 ( .A(n_402), .B(n_575), .Y(n_650) );
INVx1_ASAP7_75t_L g501 ( .A(n_403), .Y(n_501) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_403), .Y(n_633) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g1086 ( .A(n_407), .Y(n_1086) );
NAND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g419 ( .A(n_408), .Y(n_419) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_410), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g660 ( .A(n_410), .Y(n_660) );
AND2x6_ASAP7_75t_L g676 ( .A(n_410), .B(n_491), .Y(n_676) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g578 ( .A(n_413), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g659 ( .A(n_413), .Y(n_659) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_418), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g856 ( .A1(n_418), .A2(n_857), .B(n_863), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g1146 ( .A1(n_418), .A2(n_1147), .B(n_1148), .Y(n_1146) );
AOI332xp33_ASAP7_75t_L g487 ( .A1(n_421), .A2(n_488), .A3(n_493), .B1(n_495), .B2(n_497), .B3(n_499), .C1(n_502), .C2(n_506), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g764 ( .A1(n_421), .A2(n_427), .B1(n_433), .B2(n_765), .C1(n_766), .C2(n_767), .Y(n_764) );
AOI222xp33_ASAP7_75t_L g972 ( .A1(n_421), .A2(n_427), .B1(n_433), .B2(n_953), .C1(n_973), .C2(n_974), .Y(n_972) );
AOI322xp5_ASAP7_75t_L g1090 ( .A1(n_421), .A2(n_499), .A3(n_1091), .B1(n_1093), .B2(n_1096), .C1(n_1097), .C2(n_1098), .Y(n_1090) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g697 ( .A(n_423), .B(n_426), .Y(n_697) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g538 ( .A(n_424), .Y(n_538) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g483 ( .A1(n_427), .A2(n_484), .B(n_485), .Y(n_483) );
INVxp67_ASAP7_75t_L g840 ( .A(n_427), .Y(n_840) );
INVx1_ASAP7_75t_L g1083 ( .A(n_427), .Y(n_1083) );
AOI222xp33_ASAP7_75t_L g1431 ( .A1(n_427), .A2(n_1086), .B1(n_1088), .B2(n_1423), .C1(n_1432), .C2(n_1433), .Y(n_1431) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g505 ( .A(n_432), .Y(n_505) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_432), .Y(n_664) );
BUFx3_ASAP7_75t_L g862 ( .A(n_432), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_433), .A2(n_454), .B(n_480), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g1448 ( .A1(n_433), .A2(n_480), .B(n_1449), .Y(n_1448) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_437), .B(n_482), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g794 ( .A(n_437), .B(n_795), .Y(n_794) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_437), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_437), .B(n_976), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_437), .B(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1429 ( .A(n_437), .Y(n_1429) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g598 ( .A(n_440), .B(n_588), .Y(n_598) );
INVx2_ASAP7_75t_L g671 ( .A(n_440), .Y(n_671) );
BUFx3_ASAP7_75t_L g1043 ( .A(n_440), .Y(n_1043) );
XOR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_507), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_478), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_463), .B1(n_471), .B2(n_475), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_459), .B2(n_460), .C(n_461), .Y(n_456) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_457), .A2(n_518), .B1(n_519), .B2(n_522), .Y(n_517) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_457), .Y(n_919) );
OAI21xp33_ASAP7_75t_L g958 ( .A1(n_459), .A2(n_461), .B(n_959), .Y(n_958) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_461), .A2(n_542), .B1(n_751), .B2(n_755), .C(n_785), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_461), .A2(n_805), .B1(n_1067), .B2(n_1068), .C(n_1069), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1414 ( .A1(n_461), .A2(n_542), .B1(n_811), .B2(n_1415), .C(n_1416), .Y(n_1414) );
INVx3_ASAP7_75t_L g615 ( .A(n_462), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_463) );
BUFx4f_ASAP7_75t_SL g1133 ( .A(n_465), .Y(n_1133) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g927 ( .A(n_466), .Y(n_927) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g473 ( .A(n_467), .Y(n_473) );
BUFx4f_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
OR2x4_ASAP7_75t_L g624 ( .A(n_467), .B(n_608), .Y(n_624) );
BUFx3_ASAP7_75t_L g773 ( .A(n_467), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_469), .A2(n_747), .B1(n_761), .B2(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
INVx3_ASAP7_75t_L g921 ( .A(n_470), .Y(n_921) );
INVx1_ASAP7_75t_L g962 ( .A(n_470), .Y(n_962) );
INVx1_ASAP7_75t_L g918 ( .A(n_473), .Y(n_918) );
NAND4xp25_ASAP7_75t_SL g478 ( .A(n_479), .B(n_481), .C(n_483), .D(n_487), .Y(n_478) );
OR3x1_ASAP7_75t_L g977 ( .A(n_480), .B(n_978), .C(n_979), .Y(n_977) );
AND2x4_ASAP7_75t_L g685 ( .A(n_486), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_486), .Y(n_1088) );
BUFx3_ASAP7_75t_L g1092 ( .A(n_489), .Y(n_1092) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g498 ( .A(n_491), .Y(n_498) );
AND2x2_ASAP7_75t_L g573 ( .A(n_491), .B(n_574), .Y(n_573) );
BUFx3_ASAP7_75t_L g667 ( .A(n_491), .Y(n_667) );
BUFx3_ASAP7_75t_L g848 ( .A(n_491), .Y(n_848) );
INVx1_ASAP7_75t_L g1032 ( .A(n_491), .Y(n_1032) );
BUFx6f_ASAP7_75t_L g1100 ( .A(n_491), .Y(n_1100) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AOI211xp5_ASAP7_75t_L g845 ( .A1(n_499), .A2(n_846), .B(n_856), .C(n_865), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_499), .Y(n_1147) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g674 ( .A(n_504), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_505), .Y(n_675) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
XNOR2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_634), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_570), .C(n_603), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_544), .Y(n_513) );
OAI33xp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_517), .A3(n_523), .B1(n_529), .B2(n_534), .B3(n_539), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_L g915 ( .A(n_516), .Y(n_915) );
OAI22xp5_ASAP7_75t_SL g546 ( .A1(n_518), .A2(n_540), .B1(n_547), .B2(n_550), .Y(n_546) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_519), .A2(n_540), .B1(n_541), .B2(n_543), .Y(n_539) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_522), .A2(n_543), .B1(n_560), .B2(n_563), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_527), .B2(n_528), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_524), .A2(n_531), .B1(n_554), .B2(n_556), .Y(n_553) );
INVx1_ASAP7_75t_L g966 ( .A(n_525), .Y(n_966) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g607 ( .A(n_526), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g1063 ( .A(n_526), .Y(n_1063) );
BUFx6f_ASAP7_75t_L g1138 ( .A(n_526), .Y(n_1138) );
BUFx6f_ASAP7_75t_L g1387 ( .A(n_526), .Y(n_1387) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_527), .A2(n_533), .B1(n_547), .B2(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_532), .B2(n_533), .Y(n_529) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI33xp33_ASAP7_75t_L g713 ( .A1(n_535), .A2(n_714), .A3(n_716), .B1(n_719), .B2(n_723), .B3(n_725), .Y(n_713) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g925 ( .A(n_537), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_541), .A2(n_917), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI33xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .A3(n_553), .B1(n_559), .B2(n_564), .B3(n_567), .Y(n_544) );
OAI33xp33_ASAP7_75t_L g979 ( .A1(n_545), .A2(n_762), .A3(n_980), .B1(n_984), .B2(n_987), .B3(n_990), .Y(n_979) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g569 ( .A(n_551), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g1439 ( .A1(n_551), .A2(n_1421), .B1(n_1440), .B2(n_1441), .Y(n_1439) );
INVx4_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g655 ( .A(n_552), .Y(n_655) );
INVx2_ASAP7_75t_SL g745 ( .A(n_552), .Y(n_745) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_552), .Y(n_855) );
INVx1_ASAP7_75t_L g911 ( .A(n_552), .Y(n_911) );
INVx2_ASAP7_75t_L g986 ( .A(n_552), .Y(n_986) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g646 ( .A(n_555), .Y(n_646) );
BUFx2_ASAP7_75t_L g754 ( .A(n_555), .Y(n_754) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_557), .A2(n_747), .B1(n_748), .B2(n_751), .Y(n_746) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g859 ( .A(n_558), .Y(n_859) );
INVx1_ASAP7_75t_L g989 ( .A(n_558), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g857 ( .A1(n_560), .A2(n_858), .B1(n_859), .B2(n_860), .C(n_861), .Y(n_857) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI33xp33_ASAP7_75t_L g890 ( .A1(n_564), .A2(n_863), .A3(n_891), .B1(n_899), .B2(n_903), .B3(n_906), .Y(n_890) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_568), .A2(n_1011), .B1(n_1039), .B2(n_1041), .C(n_1042), .Y(n_1038) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI31xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_584), .A3(n_592), .B(n_599), .Y(n_570) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVxp67_ASAP7_75t_L g596 ( .A(n_575), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_580), .B2(n_581), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_577), .A2(n_613), .B1(n_617), .B2(n_620), .Y(n_612) );
BUFx3_ASAP7_75t_L g932 ( .A(n_578), .Y(n_932) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g935 ( .A(n_583), .Y(n_935) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g938 ( .A(n_586), .Y(n_938) );
OR2x6_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x6_ASAP7_75t_L g595 ( .A(n_587), .B(n_596), .Y(n_595) );
BUFx4f_ASAP7_75t_L g743 ( .A(n_587), .Y(n_743) );
INVxp67_ASAP7_75t_L g759 ( .A(n_587), .Y(n_759) );
INVx1_ASAP7_75t_L g896 ( .A(n_587), .Y(n_896) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx2_ASAP7_75t_L g940 ( .A(n_591), .Y(n_940) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_594), .B(n_1168), .Y(n_1167) );
AND2x4_ASAP7_75t_SL g1402 ( .A(n_594), .B(n_1403), .Y(n_1402) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx3_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
CKINVDCx16_ASAP7_75t_R g942 ( .A(n_598), .Y(n_942) );
OAI31xp33_ASAP7_75t_L g928 ( .A1(n_599), .A2(n_929), .A3(n_936), .B(n_941), .Y(n_928) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g1168 ( .A(n_601), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_601), .B(n_1160), .Y(n_1403) );
OAI31xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_609), .A3(n_621), .B(n_628), .Y(n_603) );
INVx2_ASAP7_75t_SL g876 ( .A(n_605), .Y(n_876) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g877 ( .A(n_607), .Y(n_877) );
CKINVDCx8_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx3_ASAP7_75t_L g882 ( .A(n_614), .Y(n_882) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x4_ASAP7_75t_L g618 ( .A(n_615), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_617), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g886 ( .A(n_624), .Y(n_886) );
BUFx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g888 ( .A(n_626), .Y(n_888) );
INVx1_ASAP7_75t_L g828 ( .A(n_627), .Y(n_828) );
BUFx3_ASAP7_75t_L g923 ( .A(n_627), .Y(n_923) );
BUFx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AND2x4_ASAP7_75t_L g872 ( .A(n_630), .B(n_632), .Y(n_872) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND3x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_693), .C(n_699), .Y(n_635) );
O2A1O1Ixp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_661), .B(n_683), .C(n_684), .Y(n_636) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g1028 ( .A(n_639), .Y(n_1028) );
INVx4_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_643), .A2(n_901), .B1(n_904), .B2(n_905), .Y(n_903) );
INVx5_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx3_ASAP7_75t_L g1044 ( .A(n_650), .Y(n_1044) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g1371 ( .A(n_658), .Y(n_1371) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_SL g1361 ( .A(n_663), .Y(n_1361) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_673), .B(n_676), .Y(n_665) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g847 ( .A(n_671), .Y(n_847) );
INVx1_ASAP7_75t_L g1034 ( .A(n_676), .Y(n_1034) );
AOI21xp5_ASAP7_75t_SL g1362 ( .A1(n_676), .A2(n_1363), .B(n_1365), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g1046 ( .A(n_678), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_678), .A2(n_1037), .B1(n_1367), .B2(n_1368), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_679), .A2(n_682), .B1(n_689), .B2(n_692), .Y(n_688) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_681), .Y(n_1037) );
A2O1A1Ixp33_ASAP7_75t_L g1055 ( .A1(n_683), .A2(n_1056), .B(n_1060), .C(n_1077), .Y(n_1055) );
INVx1_ASAP7_75t_L g691 ( .A(n_687), .Y(n_691) );
INVx1_ASAP7_75t_L g1022 ( .A(n_687), .Y(n_1022) );
AND2x4_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx2_ASAP7_75t_L g999 ( .A(n_692), .Y(n_999) );
INVx2_ASAP7_75t_L g1398 ( .A(n_692), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_698), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g1023 ( .A1(n_694), .A2(n_1024), .B(n_1025), .Y(n_1023) );
AOI21xp33_ASAP7_75t_SL g1379 ( .A1(n_694), .A2(n_1380), .B(n_1381), .Y(n_1379) );
INVx8_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g839 ( .A(n_697), .Y(n_839) );
AND4x1_ASAP7_75t_SL g699 ( .A(n_700), .B(n_708), .C(n_713), .D(n_728), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_704), .B2(n_705), .Y(n_700) );
AND2x4_ASAP7_75t_L g705 ( .A(n_703), .B(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g729 ( .A(n_703), .B(n_718), .Y(n_729) );
INVx1_ASAP7_75t_L g1003 ( .A(n_705), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_705), .A2(n_1002), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx5_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI33xp33_ASAP7_75t_L g1384 ( .A1(n_715), .A2(n_1385), .A3(n_1386), .B1(n_1389), .B2(n_1390), .B3(n_1392), .Y(n_1384) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx8_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g1117 ( .A1(n_726), .A2(n_1118), .B(n_1119), .C(n_1120), .Y(n_1117) );
INVx3_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx3_ASAP7_75t_L g1400 ( .A(n_729), .Y(n_1400) );
INVx1_ASAP7_75t_L g1158 ( .A(n_731), .Y(n_1158) );
XNOR2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_946), .Y(n_731) );
XOR2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_796), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
XNOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_770), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_764), .C(n_768), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_763), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_743), .A2(n_898), .B1(n_1069), .B2(n_1095), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_745), .A2(n_758), .B1(n_760), .B2(n_761), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_745), .A2(n_963), .B1(n_991), .B2(n_992), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_745), .A2(n_895), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
INVx4_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g901 ( .A(n_749), .Y(n_901) );
INVx2_ASAP7_75t_L g981 ( .A(n_749), .Y(n_981) );
INVx4_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_753), .A2(n_968), .B1(n_988), .B2(n_989), .Y(n_987) );
INVx4_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_778), .B(n_791), .C(n_794), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_773), .A2(n_961), .B1(n_962), .B2(n_963), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_774), .A2(n_897), .B1(n_905), .B2(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1110 ( .A(n_775), .Y(n_1110) );
BUFx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g823 ( .A(n_776), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .C(n_787), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI221xp5_ASAP7_75t_SL g1111 ( .A1(n_783), .A2(n_1112), .B1(n_1113), .B2(n_1115), .C(n_1116), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_785), .A2(n_902), .B1(n_912), .B2(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g970 ( .A(n_791), .Y(n_970) );
A2O1A1Ixp33_ASAP7_75t_L g1410 ( .A1(n_791), .A2(n_1411), .B(n_1422), .C(n_1426), .Y(n_1410) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_792), .A2(n_801), .B(n_835), .Y(n_800) );
INVx1_ASAP7_75t_L g1047 ( .A(n_792), .Y(n_1047) );
BUFx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g1141 ( .A(n_793), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_868), .B1(n_869), .B2(n_945), .Y(n_796) );
INVx1_ASAP7_75t_L g945 ( .A(n_797), .Y(n_945) );
BUFx2_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_866), .B(n_867), .Y(n_798) );
AND3x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_836), .C(n_845), .Y(n_799) );
AOI31xp33_ASAP7_75t_L g867 ( .A1(n_800), .A2(n_836), .A3(n_845), .B(n_866), .Y(n_867) );
NAND3xp33_ASAP7_75t_SL g801 ( .A(n_802), .B(n_818), .C(n_821), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_808), .B1(n_812), .B2(n_815), .Y(n_802) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_811), .A2(n_900), .B1(n_909), .B2(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g1016 ( .A(n_825), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_826), .A2(n_1132), .B1(n_1133), .B2(n_1134), .Y(n_1131) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_829) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_842), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B1(n_853), .B2(n_854), .Y(n_849) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_851), .Y(n_1040) );
INVx3_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_852), .Y(n_908) );
INVx4_ASAP7_75t_L g1441 ( .A(n_852), .Y(n_1441) );
INVx6_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx5_ASAP7_75t_L g898 ( .A(n_855), .Y(n_898) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g943 ( .A(n_870), .Y(n_943) );
OAI211xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_873), .B(n_889), .C(n_928), .Y(n_870) );
CKINVDCx14_ASAP7_75t_R g871 ( .A(n_872), .Y(n_871) );
NOR3xp33_ASAP7_75t_SL g873 ( .A(n_874), .B(n_878), .C(n_885), .Y(n_873) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_883), .A2(n_932), .B1(n_933), .B2(n_934), .Y(n_931) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_913), .Y(n_889) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_897), .B2(n_898), .Y(n_891) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_892), .A2(n_904), .B1(n_917), .B2(n_919), .Y(n_916) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_909), .B1(n_910), .B2(n_912), .Y(n_906) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
INVx3_ASAP7_75t_L g985 ( .A(n_908), .Y(n_985) );
BUFx3_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
OAI33xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_916), .A3(n_920), .B1(n_922), .B2(n_924), .B3(n_926), .Y(n_913) );
BUFx3_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_923), .A2(n_1006), .B1(n_1007), .B2(n_1009), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_923), .A2(n_1014), .B1(n_1015), .B2(n_1017), .C(n_1018), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_923), .A2(n_1123), .B1(n_1124), .B2(n_1126), .Y(n_1122) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_927), .B(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_948), .A2(n_1051), .B1(n_1052), .B2(n_1156), .Y(n_947) );
INVx1_ASAP7_75t_L g1156 ( .A(n_948), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_993), .B1(n_1049), .B2(n_1050), .Y(n_948) );
INVx2_ASAP7_75t_L g1049 ( .A(n_949), .Y(n_1049) );
AOI211x1_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_970), .B(n_971), .C(n_977), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_952), .B(n_956), .Y(n_951) );
NOR3xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_964), .C(n_965), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_959), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_961), .A2(n_969), .B1(n_985), .B2(n_986), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_986), .A2(n_991), .B1(n_1068), .B2(n_1103), .Y(n_1102) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
AND3x2_ASAP7_75t_L g995 ( .A(n_996), .B(n_1023), .C(n_1026), .Y(n_995) );
AOI211xp5_ASAP7_75t_SL g996 ( .A1(n_997), .A2(n_998), .B(n_1000), .C(n_1004), .Y(n_996) );
INVxp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVxp67_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
OAI31xp33_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1035), .A3(n_1045), .B(n_1047), .Y(n_1026) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1032), .Y(n_1376) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_1043), .Y(n_1101) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1043), .Y(n_1438) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1104), .B1(n_1105), .B2(n_1155), .Y(n_1052) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1053), .Y(n_1155) );
NOR2x1_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1079), .Y(n_1054) );
NOR3xp33_ASAP7_75t_SL g1060 ( .A(n_1061), .B(n_1070), .C(n_1071), .Y(n_1060) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_L g1388 ( .A(n_1067), .Y(n_1388) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1090), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1086), .B1(n_1087), .B2(n_1088), .Y(n_1084) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
NAND4xp75_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1142), .C(n_1151), .D(n_1152), .Y(n_1107) );
OAI21x1_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1121), .B(n_1140), .Y(n_1108) );
OAI21xp5_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1111), .B(n_1117), .Y(n_1109) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1114), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1127), .B1(n_1131), .B2(n_1135), .Y(n_1121) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
AOI211x1_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1144), .B(n_1146), .C(n_1150), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1166), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
NOR2xp33_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1164), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1162), .B(n_1165), .Y(n_1451) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1162), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
NOR2xp33_ASAP7_75t_L g1455 ( .A(n_1165), .B(n_1453), .Y(n_1455) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
OAI21xp33_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1175), .B(n_1355), .Y(n_1169) );
INVx4_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1235 ( .A(n_1172), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
AND2x6_ASAP7_75t_L g1183 ( .A(n_1173), .B(n_1184), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1187 ( .A(n_1173), .B(n_1188), .Y(n_1187) );
AND2x6_ASAP7_75t_L g1190 ( .A(n_1173), .B(n_1191), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1173), .B(n_1174), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1173), .B(n_1174), .Y(n_1225) );
OAI21xp5_ASAP7_75t_L g1452 ( .A1(n_1174), .A2(n_1453), .B(n_1454), .Y(n_1452) );
AOI221xp5_ASAP7_75t_SL g1175 ( .A1(n_1176), .A2(n_1236), .B1(n_1293), .B2(n_1295), .C(n_1322), .Y(n_1175) );
A2O1A1Ixp33_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1210), .B(n_1221), .C(n_1230), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1205), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1195), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1180), .B(n_1202), .Y(n_1247) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1180), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1180), .B(n_1317), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1192), .Y(n_1180) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1181), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1181), .B(n_1220), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1181), .B(n_1215), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1186), .Y(n_1181) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1183), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1185), .B(n_1189), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1192), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1192), .Y(n_1220) );
AND3x1_ASAP7_75t_L g1265 ( .A(n_1192), .B(n_1196), .C(n_1217), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1192), .B(n_1215), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1192), .B(n_1196), .Y(n_1274) );
OAI32xp33_ASAP7_75t_L g1351 ( .A1(n_1192), .A2(n_1266), .A3(n_1276), .B1(n_1352), .B2(n_1354), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1195), .B(n_1281), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1195), .B(n_1216), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1201), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1196), .B(n_1219), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1196), .B(n_1288), .Y(n_1334) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_1197), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1197), .B(n_1219), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1197), .B(n_1247), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1197), .B(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1197), .B(n_1281), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1243 ( .A(n_1201), .B(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1201), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1201), .B(n_1267), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1269 ( .A(n_1201), .B(n_1270), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1201), .B(n_1262), .Y(n_1321) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1202), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1202), .B(n_1207), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1202), .B(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1202), .B(n_1227), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1202), .B(n_1207), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1202), .B(n_1244), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1202), .B(n_1215), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1202), .B(n_1273), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1202), .B(n_1223), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1205), .Y(n_1238) );
A2O1A1Ixp33_ASAP7_75t_L g1241 ( .A1(n_1205), .A2(n_1242), .B(n_1243), .C(n_1245), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1205), .B(n_1256), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1205), .B(n_1339), .Y(n_1338) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1206), .B(n_1227), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1206), .B(n_1256), .Y(n_1329) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1207), .B(n_1227), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1207), .B(n_1263), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1207), .B(n_1227), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1212), .B1(n_1214), .B2(n_1218), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1212), .B(n_1240), .Y(n_1239) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1213), .B(n_1281), .Y(n_1288) );
O2A1O1Ixp33_ASAP7_75t_SL g1290 ( .A1(n_1213), .A2(n_1217), .B(n_1291), .C(n_1292), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1213), .B(n_1214), .Y(n_1324) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1214), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .Y(n_1214) );
AOI221xp5_ASAP7_75t_L g1248 ( .A1(n_1215), .A2(n_1249), .B1(n_1253), .B2(n_1255), .C(n_1258), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1215), .B(n_1217), .Y(n_1254) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1216), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1216), .B(n_1219), .Y(n_1298) );
OAI332xp33_ASAP7_75t_L g1258 ( .A1(n_1217), .A2(n_1223), .A3(n_1227), .B1(n_1259), .B2(n_1261), .B3(n_1262), .C1(n_1264), .C2(n_1266), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1217), .B(n_1220), .Y(n_1281) );
O2A1O1Ixp33_ASAP7_75t_L g1303 ( .A1(n_1218), .A2(n_1304), .B(n_1306), .C(n_1307), .Y(n_1303) );
AOI22xp5_ASAP7_75t_L g1296 ( .A1(n_1220), .A2(n_1297), .B1(n_1299), .B2(n_1301), .Y(n_1296) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1227), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1223), .B(n_1251), .Y(n_1250) );
CKINVDCx6p67_ASAP7_75t_R g1256 ( .A(n_1223), .Y(n_1256) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_1223), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1223), .B(n_1227), .Y(n_1309) );
OR2x6_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1226), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1224), .B(n_1226), .Y(n_1242) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1227), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1227), .B(n_1256), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1227), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1227), .B(n_1256), .Y(n_1335) );
AND2x4_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1229), .Y(n_1227) );
INVx2_ASAP7_75t_SL g1282 ( .A(n_1230), .Y(n_1282) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_1230), .Y(n_1294) );
OAI22xp5_ASAP7_75t_SL g1231 ( .A1(n_1232), .A2(n_1233), .B1(n_1234), .B2(n_1235), .Y(n_1231) );
NAND5xp2_ASAP7_75t_SL g1236 ( .A(n_1237), .B(n_1241), .C(n_1248), .D(n_1268), .E(n_1283), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1238), .B(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1240), .Y(n_1291) );
OAI211xp5_ASAP7_75t_SL g1295 ( .A1(n_1242), .A2(n_1296), .B(n_1303), .C(n_1312), .Y(n_1295) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1244), .Y(n_1354) );
OAI21xp5_ASAP7_75t_L g1336 ( .A1(n_1245), .A2(n_1261), .B(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1250), .B(n_1285), .Y(n_1348) );
CKINVDCx6p67_ASAP7_75t_R g1251 ( .A(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1252), .B(n_1260), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_1252), .A2(n_1269), .B1(n_1271), .B2(n_1273), .C(n_1275), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_1252), .A2(n_1313), .B1(n_1318), .B2(n_1321), .Y(n_1312) );
O2A1O1Ixp33_ASAP7_75t_L g1349 ( .A1(n_1252), .A2(n_1311), .B(n_1350), .C(n_1351), .Y(n_1349) );
A2O1A1Ixp33_ASAP7_75t_L g1332 ( .A1(n_1253), .A2(n_1260), .B(n_1333), .C(n_1335), .Y(n_1332) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_1255), .A2(n_1267), .B1(n_1324), .B2(n_1325), .C(n_1330), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1257), .Y(n_1255) );
NOR2xp33_ASAP7_75t_L g1271 ( .A(n_1256), .B(n_1272), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1256), .B(n_1279), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1256), .B(n_1262), .Y(n_1347) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1257), .Y(n_1279) );
AOI21xp33_ASAP7_75t_L g1330 ( .A1(n_1257), .A2(n_1308), .B(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1262), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1262), .B(n_1353), .Y(n_1352) );
A2O1A1Ixp33_ASAP7_75t_L g1307 ( .A1(n_1264), .A2(n_1308), .B(n_1309), .C(n_1310), .Y(n_1307) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1267), .Y(n_1277) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1272), .Y(n_1306) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
OAI211xp5_ASAP7_75t_SL g1275 ( .A1(n_1276), .A2(n_1277), .B(n_1278), .C(n_1282), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1280), .Y(n_1278) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1281), .Y(n_1341) );
O2A1O1Ixp33_ASAP7_75t_L g1283 ( .A1(n_1284), .A2(n_1287), .B(n_1289), .C(n_1290), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
NAND3xp33_ASAP7_75t_SL g1343 ( .A(n_1288), .B(n_1344), .C(n_1345), .Y(n_1343) );
NOR2xp33_ASAP7_75t_L g1318 ( .A(n_1292), .B(n_1319), .Y(n_1318) );
INVx3_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
AOI21xp33_ASAP7_75t_L g1325 ( .A1(n_1294), .A2(n_1326), .B(n_1328), .Y(n_1325) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVxp67_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVxp67_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
NOR2xp33_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1316), .Y(n_1314) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1317), .Y(n_1340) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
NAND5xp2_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1332), .C(n_1336), .D(n_1342), .E(n_1349), .Y(n_1322) );
INVx2_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1335), .Y(n_1344) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1339), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1341), .Y(n_1339) );
AOI21xp5_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1347), .B(n_1348), .Y(n_1342) );
INVxp67_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND3xp33_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1379), .C(n_1382), .Y(n_1358) );
OAI21xp33_ASAP7_75t_L g1359 ( .A1(n_1360), .A2(n_1369), .B(n_1377), .Y(n_1359) );
BUFx2_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
NOR3xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1397), .C(n_1399), .Y(n_1382) );
NAND2xp5_ASAP7_75t_SL g1383 ( .A(n_1384), .B(n_1394), .Y(n_1383) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx2_ASAP7_75t_SL g1399 ( .A(n_1400), .Y(n_1399) );
BUFx4f_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVxp67_ASAP7_75t_SL g1404 ( .A(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
HB1xp67_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1430), .Y(n_1409) );
NOR3xp33_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1413), .C(n_1417), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1428), .Y(n_1426) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NAND4xp25_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1434), .C(n_1446), .D(n_1448), .Y(n_1430) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
HB1xp67_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
endmodule