module fake_jpeg_1888_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_60),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_70),
.B1(n_49),
.B2(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_48),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_44),
.B1(n_45),
.B2(n_39),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_49),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_40),
.B1(n_44),
.B2(n_53),
.Y(n_77)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_72),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_41),
.C(n_43),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_80),
.A3(n_81),
.B1(n_74),
.B2(n_83),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_82),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_57),
.B1(n_54),
.B2(n_66),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_51),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_62),
.B1(n_57),
.B2(n_54),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_94),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_78),
.B(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_11),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_111),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_17),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_20),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_8),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_9),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_113),
.B(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_11),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_13),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_34),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_93),
.C(n_16),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_119),
.C(n_126),
.Y(n_137)
);

XOR2x2_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_93),
.B1(n_14),
.B2(n_19),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_102),
.B1(n_106),
.B2(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_127),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_21),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.C1(n_27),
.C2(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_125),
.B1(n_101),
.B2(n_122),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_119),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_126),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_141),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_137),
.B(n_131),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_143),
.C(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_139),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_146),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_35),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);


endmodule