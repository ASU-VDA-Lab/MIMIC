module fake_jpeg_2888_n_297 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_256;
wire n_151;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_32),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_60),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_39),
.B(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_54),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_74),
.B1(n_79),
.B2(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_90),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_54),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_53),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_26),
.B1(n_23),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_32),
.B1(n_14),
.B2(n_25),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_84),
.B1(n_88),
.B2(n_19),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_27),
.B1(n_19),
.B2(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_34),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_18),
.B1(n_15),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_27),
.B1(n_19),
.B2(n_16),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_15),
.B1(n_18),
.B2(n_34),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_53),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx10_ASAP7_75t_R g155 ( 
.A(n_96),
.Y(n_155)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_127),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_29),
.B1(n_57),
.B2(n_49),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_120),
.B1(n_125),
.B2(n_129),
.Y(n_148)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_40),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_118),
.Y(n_137)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_115),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_31),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_60),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_91),
.B(n_63),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_49),
.B1(n_48),
.B2(n_57),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_126),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_35),
.B(n_33),
.C(n_28),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_133),
.Y(n_140)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_28),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_131),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_67),
.B(n_53),
.Y(n_127)
);

CKINVDCx11_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_67),
.A2(n_83),
.B1(n_46),
.B2(n_16),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_59),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_41),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_103),
.B(n_116),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_43),
.B(n_65),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_160),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_65),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_127),
.C(n_119),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_10),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_9),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_92),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_98),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_182),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_179),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_122),
.B1(n_120),
.B2(n_132),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_170),
.B1(n_174),
.B2(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_127),
.C(n_130),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_177),
.C(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_112),
.B1(n_110),
.B2(n_117),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_104),
.B1(n_101),
.B2(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_190),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_106),
.C(n_95),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_126),
.B1(n_102),
.B2(n_133),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_114),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_185),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_87),
.B1(n_108),
.B2(n_114),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_149),
.B1(n_152),
.B2(n_156),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_114),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_96),
.C(n_123),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_139),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_87),
.B1(n_25),
.B2(n_16),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_141),
.B1(n_163),
.B2(n_135),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_63),
.C(n_16),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_149),
.C(n_152),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_201),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_136),
.B(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_206),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_162),
.B(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_194),
.B(n_189),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_207),
.C(n_208),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_209),
.B1(n_175),
.B2(n_172),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_134),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_165),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_158),
.B1(n_156),
.B2(n_154),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_178),
.B1(n_167),
.B2(n_169),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_158),
.A3(n_157),
.B1(n_145),
.B2(n_161),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_221),
.B1(n_223),
.B2(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_203),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_225),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_168),
.B1(n_183),
.B2(n_186),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_177),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_226),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_193),
.B(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_230),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_196),
.B(n_164),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_157),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_188),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_145),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_198),
.C(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_236),
.C(n_248),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_198),
.C(n_228),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_247),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_210),
.B1(n_233),
.B2(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_204),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_249),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_223),
.C(n_221),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_199),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_218),
.B(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_251),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_257),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_215),
.B1(n_209),
.B2(n_227),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_254),
.Y(n_268)
);

AO221x1_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_200),
.B1(n_230),
.B2(n_227),
.C(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_260),
.Y(n_271)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_214),
.B1(n_229),
.B2(n_197),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_262),
.B1(n_25),
.B2(n_16),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_159),
.A3(n_197),
.B1(n_151),
.B2(n_13),
.C1(n_8),
.C2(n_161),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_8),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NOR2x1p5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_159),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_236),
.Y(n_266)
);

OAI321xp33_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_246),
.A3(n_248),
.B1(n_244),
.B2(n_249),
.C(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_264),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_151),
.C(n_159),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_260),
.C(n_263),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_151),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_272),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_280),
.B(n_271),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_250),
.C(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_281),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_261),
.B(n_250),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_285),
.B(n_0),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_268),
.C(n_270),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_279),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_265),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_278),
.C(n_8),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_275),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_291),
.A3(n_0),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_4),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_0),
.C(n_2),
.Y(n_294)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_0),
.A3(n_3),
.B1(n_4),
.B2(n_293),
.C(n_291),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_296),
.Y(n_297)
);


endmodule