module real_jpeg_17982_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_0),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_0),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_1),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_1),
.B(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_2),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_2),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_2),
.B(n_144),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_2),
.B(n_41),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_2),
.B(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_5),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_5),
.B(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_5),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_5),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_5),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_5),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_6),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_6),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_6),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_7),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_11),
.B1(n_39),
.B2(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_8),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_8),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_8),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_8),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_8),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_8),
.B(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_9),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_9),
.B(n_105),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_9),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_9),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_9),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_62),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_10),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_10),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_10),
.B(n_33),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_10),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_11),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_11),
.B(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_11),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_11),
.B(n_395),
.Y(n_394)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_12),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_14),
.Y(n_191)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_14),
.Y(n_289)
);

NAND2x1_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_15),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_15),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_15),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_15),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_15),
.B(n_297),
.Y(n_296)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_368),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_208),
.B(n_367),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_173),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_20),
.B(n_173),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_100),
.Y(n_20)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_21),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.C(n_85),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_23),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.C(n_50),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_24),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_28),
.C(n_32),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_25),
.B(n_143),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_37),
.A2(n_38),
.B1(n_50),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_38),
.A2(n_226),
.B(n_229),
.Y(n_225)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_48),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_61),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_51),
.A2(n_52),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_52),
.B(n_108),
.C(n_153),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_54),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_56),
.B(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_61),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_66),
.A2(n_86),
.B1(n_87),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_66),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.C(n_80),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_67),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.C(n_75),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_68),
.A2(n_75),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_68),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_68),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_70),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_71),
.B(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_75),
.Y(n_224)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_76),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_204),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_80),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_83),
.Y(n_228)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_90),
.C(n_96),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_90),
.A2(n_91),
.B1(n_240),
.B2(n_241),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_91),
.B(n_235),
.C(n_240),
.Y(n_234)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_99),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_149),
.B1(n_171),
.B2(n_172),
.Y(n_100)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_138),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_102),
.B(n_139),
.C(n_140),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.C(n_125),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_103),
.B(n_115),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_108),
.C(n_111),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_108),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_108),
.A2(n_114),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_109),
.Y(n_291)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_109),
.Y(n_319)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_113),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_116),
.A2(n_122),
.B1(n_123),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_118),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_120),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_122),
.B(n_260),
.C(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_122),
.A2(n_123),
.B1(n_260),
.B2(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_SL g178 ( 
.A(n_125),
.B(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_131),
.C(n_135),
.Y(n_148)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_134),
.Y(n_392)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_136),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_142),
.B(n_147),
.C(n_148),
.Y(n_408)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_149),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_150),
.B(n_157),
.C(n_158),
.Y(n_409)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_153),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_153),
.A2(n_155),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_154),
.B(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_159),
.B(n_163),
.C(n_167),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_166),
.Y(n_278)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_171),
.B(n_372),
.C(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_180),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_202),
.C(n_205),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_193),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_187),
.B(n_193),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_192),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_191),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_194),
.A2(n_197),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_197),
.A2(n_257),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_197),
.B(n_321),
.C(n_325),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_198),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_199),
.B(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_267),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.C(n_247),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_213),
.B(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_243),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_244),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.C(n_234),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_225),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_223),
.B(n_276),
.C(n_279),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_235),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_SL g309 ( 
.A(n_236),
.B(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_236),
.A2(n_316),
.B1(n_317),
.B2(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.C(n_265),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_251),
.B(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_253),
.B(n_265),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.C(n_263),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_254),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_259),
.B(n_264),
.Y(n_358)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

XOR2x1_ASAP7_75t_L g303 ( 
.A(n_261),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.C(n_366),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_361),
.B(n_365),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_347),
.B(n_360),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_312),
.B(n_346),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_300),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_273),
.B(n_300),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.C(n_292),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_283),
.A2(n_284),
.B1(n_292),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_285),
.B(n_290),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

AO22x1_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_292)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_293),
.Y(n_298)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_302),
.B(n_303),
.C(n_306),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_340),
.B(n_345),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_328),
.B(n_339),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_320),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_335),
.B(n_338),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_333),
.Y(n_338)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_344),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_359),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_SL g360 ( 
.A(n_348),
.B(n_359),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_356),
.B2(n_357),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_355),
.C(n_356),
.Y(n_364)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_364),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_410),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

AND2x2_ASAP7_75t_SL g410 ( 
.A(n_371),
.B(n_374),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_401),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_387),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_397),
.Y(n_393)
);

INVx8_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_409),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_408),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_406),
.B2(n_407),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_405),
.Y(n_407)
);


endmodule