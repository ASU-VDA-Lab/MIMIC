module fake_jpeg_2341_n_546 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_546);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_133;
wire n_419;
wire n_132;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_47),
.Y(n_111)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_53),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_56),
.Y(n_158)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_67),
.B(n_73),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_30),
.A2(n_12),
.B(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_76),
.B(n_77),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_17),
.B(n_12),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_88),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_93),
.Y(n_115)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_35),
.B(n_12),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_35),
.B(n_44),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_97),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_44),
.B(n_11),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_32),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_105),
.B(n_126),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_46),
.B(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_108),
.B(n_161),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_33),
.B1(n_21),
.B2(n_23),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_33),
.B1(n_99),
.B2(n_92),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_79),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_81),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_123),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_29),
.B1(n_22),
.B2(n_32),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_142),
.A2(n_144),
.B1(n_149),
.B2(n_34),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_57),
.A2(n_29),
.B1(n_22),
.B2(n_32),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_62),
.A2(n_32),
.B1(n_39),
.B2(n_34),
.Y(n_149)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_53),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

BUFx16f_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

CKINVDCx6p67_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_53),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_32),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_74),
.B(n_42),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_49),
.Y(n_162)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_23),
.B1(n_33),
.B2(n_94),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_178),
.B1(n_189),
.B2(n_142),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_114),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_173),
.Y(n_212)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_188),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_73),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_190),
.Y(n_217)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_47),
.B1(n_61),
.B2(n_50),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_138),
.B1(n_143),
.B2(n_158),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_56),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_72),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_83),
.B1(n_87),
.B2(n_86),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_32),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_91),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_192),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_52),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_140),
.B(n_28),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_201),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_146),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_197),
.Y(n_237)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_113),
.B(n_96),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_235)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_199),
.Y(n_229)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_107),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_75),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_203),
.B(n_208),
.Y(n_240)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_100),
.B(n_75),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_127),
.B(n_78),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_143),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_214),
.A2(n_215),
.B1(n_234),
.B2(n_238),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_149),
.B1(n_152),
.B2(n_136),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_138),
.A3(n_102),
.B1(n_148),
.B2(n_137),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_196),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_172),
.B1(n_181),
.B2(n_131),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_187),
.B(n_109),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_175),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_148),
.C(n_103),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_211),
.C(n_179),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_178),
.A2(n_133),
.B1(n_147),
.B2(n_121),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_168),
.A2(n_129),
.B1(n_117),
.B2(n_118),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_SL g239 ( 
.A(n_194),
.B(n_104),
.C(n_28),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_195),
.B(n_133),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_175),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_198),
.A2(n_145),
.B1(n_141),
.B2(n_119),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_245),
.B1(n_199),
.B2(n_182),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_201),
.A2(n_68),
.B1(n_104),
.B2(n_131),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_274),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_251),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_227),
.B(n_217),
.C(n_171),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_270),
.B(n_248),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_253),
.A2(n_262),
.B1(n_270),
.B2(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_166),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_256),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_255),
.A2(n_260),
.B(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_217),
.Y(n_256)
);

OAI32xp33_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_166),
.A3(n_167),
.B1(n_206),
.B2(n_193),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_167),
.Y(n_261)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_216),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_215),
.A2(n_202),
.B1(n_200),
.B2(n_209),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_213),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_271),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_207),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_183),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_275),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_237),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_218),
.B(n_228),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_235),
.B1(n_238),
.B2(n_231),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_278),
.A2(n_292),
.B1(n_299),
.B2(n_275),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_231),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_288),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_286),
.A2(n_297),
.B(n_229),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_287),
.A2(n_286),
.B1(n_285),
.B2(n_277),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_232),
.C(n_222),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_290),
.B(n_259),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_233),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_271),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_255),
.B1(n_270),
.B2(n_249),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_239),
.B1(n_221),
.B2(n_220),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_261),
.B1(n_272),
.B2(n_254),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_253),
.A2(n_239),
.B(n_243),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_230),
.B1(n_186),
.B2(n_169),
.Y(n_299)
);

AO22x2_ASAP7_75t_L g303 ( 
.A1(n_252),
.A2(n_230),
.B1(n_236),
.B2(n_225),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_257),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_233),
.C(n_220),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_304),
.B(n_182),
.CI(n_176),
.CON(n_334),
.SN(n_334)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_247),
.C(n_263),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_307),
.A2(n_311),
.B1(n_312),
.B2(n_316),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_308),
.B(n_297),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_274),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_309),
.B(n_313),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_329),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_302),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_276),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_285),
.A2(n_266),
.B1(n_252),
.B2(n_260),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_314),
.A2(n_317),
.B1(n_337),
.B2(n_278),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_332),
.Y(n_339)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_262),
.B1(n_275),
.B2(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_319),
.Y(n_346)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_295),
.B(n_263),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_326),
.C(n_336),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_SL g322 ( 
.A(n_288),
.B(n_182),
.C(n_243),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_322),
.B(n_331),
.Y(n_355)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_258),
.Y(n_324)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_325),
.B(n_338),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_306),
.Y(n_327)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_333),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_284),
.B(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_228),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_291),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_279),
.B(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_267),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_352),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_342),
.A2(n_343),
.B1(n_356),
.B2(n_366),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_294),
.B1(n_290),
.B2(n_281),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_277),
.Y(n_347)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_309),
.B(n_300),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_350),
.B(n_358),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_336),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_281),
.B1(n_305),
.B2(n_304),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_338),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_303),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_335),
.B(n_296),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_361),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_280),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_287),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_303),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_321),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_365),
.B(n_370),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_311),
.A2(n_299),
.B1(n_298),
.B2(n_284),
.Y(n_366)
);

NOR3xp33_ASAP7_75t_SL g371 ( 
.A(n_368),
.B(n_334),
.C(n_322),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_228),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_385),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_372),
.B(n_400),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_316),
.C(n_330),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_386),
.C(n_388),
.Y(n_401)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_342),
.A2(n_307),
.B1(n_317),
.B2(n_328),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_377),
.A2(n_380),
.B1(n_363),
.B2(n_357),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_344),
.A2(n_333),
.B1(n_323),
.B2(n_320),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_348),
.Y(n_381)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_347),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_334),
.C(n_318),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_341),
.Y(n_387)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_297),
.C(n_319),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_392),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_344),
.A2(n_303),
.B(n_183),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_394),
.B(n_360),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_339),
.B(n_229),
.C(n_219),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_362),
.C(n_353),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_352),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_396),
.B(n_230),
.Y(n_429)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_399),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_339),
.B(n_229),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_360),
.Y(n_420)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_355),
.B(n_267),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_390),
.A2(n_391),
.B1(n_377),
.B2(n_393),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_408),
.B1(n_392),
.B2(n_384),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_410),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_340),
.B1(n_343),
.B2(n_367),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_407),
.B(n_415),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_351),
.B1(n_344),
.B2(n_363),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_364),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_369),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_418),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_413),
.A2(n_389),
.B1(n_394),
.B2(n_371),
.Y(n_437)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_376),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_414),
.B(n_225),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_369),
.C(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_422),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_346),
.C(n_219),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_421),
.B(n_425),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_393),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_219),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_225),
.C(n_236),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_398),
.C(n_375),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_182),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_204),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_28),
.C(n_40),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_432),
.A2(n_444),
.B1(n_446),
.B2(n_449),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_439),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_412),
.Y(n_436)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_453),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_SL g443 ( 
.A1(n_428),
.A2(n_38),
.B(n_42),
.C(n_40),
.Y(n_443)
);

OAI31xp33_ASAP7_75t_L g469 ( 
.A1(n_443),
.A2(n_36),
.A3(n_37),
.B(n_38),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_424),
.A2(n_210),
.B1(n_205),
.B2(n_177),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_401),
.B(n_118),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_448),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_417),
.A2(n_129),
.B1(n_117),
.B2(n_155),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_406),
.B(n_125),
.Y(n_447)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_416),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_48),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_450),
.A2(n_455),
.B(n_440),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_422),
.A2(n_124),
.B1(n_155),
.B2(n_125),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_451),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_409),
.B(n_8),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_419),
.A2(n_403),
.B1(n_427),
.B2(n_410),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_426),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_132),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_452),
.B(n_411),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_450),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_415),
.C(n_421),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_458),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_401),
.C(n_405),
.Y(n_458)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_460),
.A2(n_431),
.B1(n_441),
.B2(n_430),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_423),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_466),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_420),
.C(n_85),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_469),
.B(n_472),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_132),
.C(n_176),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_154),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_473),
.B(n_476),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_54),
.C(n_51),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_474),
.B(n_462),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_154),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_454),
.Y(n_477)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_477),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_430),
.C(n_431),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_479),
.B(n_481),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_441),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_447),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_482),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_453),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_483),
.A2(n_475),
.B(n_467),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_466),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_487),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_472),
.C(n_463),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_489),
.C(n_494),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_451),
.C(n_443),
.Y(n_489)
);

AOI221xp5_ASAP7_75t_L g492 ( 
.A1(n_465),
.A2(n_443),
.B1(n_37),
.B2(n_38),
.C(n_42),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_492),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_151),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_443),
.C(n_70),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_501),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_490),
.A2(n_55),
.B(n_45),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_498),
.A2(n_504),
.B(n_507),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_502),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_151),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_503),
.B(n_39),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_485),
.A2(n_69),
.B(n_58),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_36),
.B1(n_151),
.B2(n_68),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_505),
.A2(n_34),
.B1(n_39),
.B2(n_31),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_479),
.A2(n_78),
.B(n_8),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_31),
.C(n_39),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_0),
.Y(n_520)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_496),
.A2(n_484),
.A3(n_491),
.B1(n_478),
.B2(n_487),
.C1(n_494),
.C2(n_31),
.Y(n_512)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_512),
.A2(n_520),
.B(n_509),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_10),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_513),
.B(n_514),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_508),
.C(n_500),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_515),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_516),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_31),
.C(n_10),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_519),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_10),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_522),
.B(n_498),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_31),
.C(n_10),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_1),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_9),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_511),
.A2(n_507),
.B(n_505),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_524),
.A2(n_9),
.B(n_2),
.Y(n_536)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_527),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_531),
.C(n_510),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_519),
.C(n_517),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_514),
.A2(n_503),
.B(n_31),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_532),
.A2(n_535),
.B(n_5),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_SL g541 ( 
.A1(n_534),
.A2(n_6),
.B(n_7),
.C(n_533),
.Y(n_541)
);

A2O1A1O1Ixp25_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_9),
.B(n_2),
.C(n_3),
.D(n_5),
.Y(n_535)
);

AOI21xp33_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_525),
.B(n_530),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_523),
.A2(n_1),
.B(n_3),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_537),
.A2(n_5),
.B(n_6),
.Y(n_540)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_538),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_539),
.A2(n_540),
.B(n_541),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_6),
.B(n_7),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_542),
.C(n_6),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_6),
.B(n_7),
.Y(n_546)
);


endmodule