module real_jpeg_10631_n_1 (n_0, n_1);

input n_0;

output n_1;

wire n_2;

CKINVDCx20_ASAP7_75t_R g2 ( 
.A(n_0),
.Y(n_2)
);

CKINVDCx20_ASAP7_75t_R g1 ( 
.A(n_2),
.Y(n_1)
);


endmodule