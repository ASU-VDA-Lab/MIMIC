module fake_aes_9591_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_0), .B(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_16), .B(n_3), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_17), .B(n_15), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_13), .B1(n_11), .B2(n_5), .Y(n_22) );
AOI22x1_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_11), .B1(n_7), .B2(n_10), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
OA21x2_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_18), .B(n_11), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_24), .B(n_21), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_26), .Y(n_29) );
O2A1O1Ixp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_21), .B(n_26), .C(n_27), .Y(n_30) );
OAI211xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_23), .B(n_25), .C(n_21), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
INVxp33_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_30), .B(n_4), .Y(n_34) );
NOR2xp33_ASAP7_75t_L g35 ( .A(n_32), .B(n_4), .Y(n_35) );
BUFx3_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_33), .B(n_31), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_5), .B1(n_34), .B2(n_37), .Y(n_38) );
XNOR2xp5_ASAP7_75t_L g39 ( .A(n_38), .B(n_36), .Y(n_39) );
endmodule