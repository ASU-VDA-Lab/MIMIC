module fake_jpeg_2566_n_685 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_685);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_685;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_8),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_11),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_72),
.Y(n_171)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_74),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_76),
.Y(n_193)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_79),
.Y(n_222)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_85),
.Y(n_206)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_86),
.Y(n_197)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_89),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_91),
.Y(n_203)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_94),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_127),
.Y(n_136)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_99),
.Y(n_205)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_100),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_50),
.A2(n_31),
.B1(n_35),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_101),
.A2(n_47),
.B1(n_34),
.B2(n_32),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_105),
.Y(n_210)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_57),
.Y(n_114)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_116),
.Y(n_217)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_57),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_124),
.Y(n_226)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_38),
.Y(n_149)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_132),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_39),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_25),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_70),
.B(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_145),
.B(n_173),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_30),
.B1(n_21),
.B2(n_36),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_148),
.B(n_1),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_149),
.B(n_162),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_35),
.B1(n_21),
.B2(n_36),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_151),
.A2(n_160),
.B1(n_167),
.B2(n_172),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_21),
.B1(n_26),
.B2(n_36),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_158),
.A2(n_174),
.B1(n_202),
.B2(n_177),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_26),
.B1(n_41),
.B2(n_43),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_65),
.A2(n_43),
.B1(n_41),
.B2(n_26),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_91),
.A2(n_41),
.B1(n_43),
.B2(n_38),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_133),
.B(n_25),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_63),
.A2(n_93),
.B1(n_99),
.B2(n_62),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_75),
.A2(n_25),
.B1(n_45),
.B2(n_38),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_176),
.A2(n_208),
.B1(n_216),
.B2(n_220),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_58),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_177),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_75),
.B(n_110),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_180),
.B(n_183),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_110),
.B(n_23),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_73),
.B(n_23),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_192),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_86),
.B(n_23),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_122),
.B(n_29),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_195),
.B(n_198),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_67),
.B(n_29),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_123),
.B(n_45),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_199),
.B(n_209),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_71),
.A2(n_45),
.B1(n_29),
.B2(n_52),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_76),
.A2(n_115),
.B1(n_113),
.B2(n_107),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_79),
.B(n_52),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_102),
.B(n_52),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_24),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_81),
.A2(n_58),
.B1(n_56),
.B2(n_47),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_90),
.A2(n_58),
.B1(n_56),
.B2(n_47),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_142),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_227),
.B(n_233),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_136),
.A2(n_95),
.B1(n_34),
.B2(n_56),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_229),
.A2(n_214),
.B1(n_164),
.B2(n_169),
.Y(n_346)
);

BUFx16f_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx4_ASAP7_75t_SL g322 ( 
.A(n_230),
.Y(n_322)
);

AO21x2_ASAP7_75t_L g318 ( 
.A1(n_231),
.A2(n_246),
.B(n_262),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_177),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_235),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_24),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_236),
.B(n_257),
.Y(n_309)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_237),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_140),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_238),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_239),
.B(n_244),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_153),
.A2(n_28),
.B1(n_39),
.B2(n_97),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_240),
.A2(n_285),
.B1(n_287),
.B2(n_289),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_241),
.Y(n_345)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_143),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_134),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_243),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_146),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_245),
.A2(n_248),
.B1(n_252),
.B2(n_264),
.Y(n_330)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_137),
.A2(n_39),
.B1(n_10),
.B2(n_11),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_146),
.Y(n_249)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_176),
.A2(n_18),
.B(n_17),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_251),
.A2(n_217),
.B(n_159),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_252)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_254),
.Y(n_344)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_255),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_0),
.Y(n_257)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_259),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_168),
.B(n_0),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_147),
.Y(n_261)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_261),
.Y(n_317)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_263),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_157),
.A2(n_200),
.B1(n_188),
.B2(n_213),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_265),
.B(n_266),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_178),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_147),
.Y(n_269)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_270),
.Y(n_339)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_171),
.Y(n_271)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_272),
.B(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_150),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_278),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_182),
.B(n_141),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

BUFx6f_ASAP7_75t_SL g276 ( 
.A(n_194),
.Y(n_276)
);

INVx11_ASAP7_75t_L g368 ( 
.A(n_276),
.Y(n_368)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_170),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g280 ( 
.A(n_155),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_280),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_184),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_135),
.B(n_1),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_304),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_157),
.A2(n_188),
.B1(n_200),
.B2(n_205),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_292),
.B1(n_220),
.B2(n_167),
.Y(n_314)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_179),
.B(n_1),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_302),
.B(n_303),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_226),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_197),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_179),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_181),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_291),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_161),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_294),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_201),
.B(n_14),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_165),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_297),
.Y(n_356)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_296),
.Y(n_357)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_197),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_300),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_219),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_299),
.Y(n_360)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_139),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_159),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_151),
.B1(n_160),
.B2(n_172),
.Y(n_310)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_163),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_184),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_181),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_204),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_231),
.A2(n_161),
.B1(n_205),
.B2(n_225),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_308),
.A2(n_318),
.B1(n_338),
.B2(n_343),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_310),
.A2(n_277),
.B1(n_297),
.B2(n_288),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_314),
.A2(n_362),
.B1(n_286),
.B2(n_292),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_319),
.A2(n_254),
.B(n_296),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_219),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_348),
.C(n_367),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_234),
.A2(n_217),
.B(n_206),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_331),
.A2(n_334),
.B(n_281),
.Y(n_415)
);

O2A1O1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_155),
.B(n_184),
.C(n_187),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_279),
.A2(n_225),
.B1(n_222),
.B2(n_193),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_279),
.A2(n_222),
.B1(n_193),
.B2(n_207),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_253),
.B(n_164),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_207),
.B1(n_204),
.B2(n_196),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_353),
.A2(n_359),
.B1(n_284),
.B2(n_264),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_236),
.A2(n_196),
.B1(n_185),
.B2(n_13),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_245),
.A2(n_185),
.B1(n_3),
.B2(n_5),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_257),
.B(n_2),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_365),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_258),
.A2(n_2),
.A3(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_256),
.B(n_2),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_414),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_313),
.B(n_290),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_371),
.B(n_378),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_376),
.B1(n_383),
.B2(n_388),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_318),
.A2(n_274),
.B1(n_260),
.B2(n_283),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_375),
.A2(n_384),
.B1(n_390),
.B2(n_400),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_255),
.C(n_251),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_395),
.C(n_398),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_326),
.B(n_309),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_309),
.B(n_286),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_385),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_380),
.Y(n_427)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_318),
.A2(n_242),
.B1(n_247),
.B2(n_249),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_318),
.A2(n_293),
.B1(n_278),
.B2(n_263),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_312),
.B(n_298),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_316),
.B(n_235),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_389),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_387),
.A2(n_415),
.B1(n_349),
.B2(n_353),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_318),
.A2(n_305),
.B1(n_291),
.B2(n_275),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_312),
.B(n_268),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_276),
.B1(n_285),
.B2(n_241),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_393),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_367),
.B(n_270),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_394),
.B(n_408),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_332),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_271),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_402),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_272),
.C(n_259),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_308),
.A2(n_250),
.B1(n_299),
.B2(n_267),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_399),
.A2(n_404),
.B1(n_417),
.B2(n_362),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_314),
.A2(n_331),
.B1(n_330),
.B2(n_321),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_343),
.B(n_299),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_401),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_228),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_230),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_405),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_321),
.A2(n_304),
.B1(n_230),
.B2(n_280),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_6),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_340),
.Y(n_407)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_6),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_330),
.A2(n_280),
.B1(n_281),
.B2(n_8),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_410),
.A2(n_361),
.B1(n_360),
.B2(n_357),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_6),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_411),
.B(n_337),
.Y(n_451)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_339),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_413),
.A2(n_322),
.B1(n_360),
.B2(n_341),
.Y(n_442)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_311),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_358),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_359),
.A2(n_281),
.B1(n_8),
.B2(n_9),
.Y(n_417)
);

OAI211xp5_ASAP7_75t_L g418 ( 
.A1(n_319),
.A2(n_7),
.B(n_9),
.C(n_364),
.Y(n_418)
);

OAI31xp33_ASAP7_75t_L g434 ( 
.A1(n_418),
.A2(n_334),
.A3(n_355),
.B(n_356),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_422),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_315),
.C(n_364),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_449),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_426),
.A2(n_457),
.B1(n_383),
.B2(n_409),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_375),
.A2(n_338),
.B1(n_310),
.B2(n_347),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_439),
.B1(n_445),
.B2(n_455),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_432),
.B(n_451),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_434),
.A2(n_442),
.B1(n_454),
.B2(n_415),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_372),
.A2(n_341),
.B1(n_315),
.B2(n_357),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_342),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_323),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_446),
.C(n_452),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_355),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_377),
.C(n_379),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_361),
.B(n_337),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_450),
.A2(n_380),
.B(n_411),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_328),
.C(n_355),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_350),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_453),
.B(n_456),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_400),
.A2(n_307),
.B1(n_345),
.B2(n_329),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_384),
.A2(n_307),
.B1(n_345),
.B2(n_329),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_370),
.B(n_371),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_390),
.A2(n_307),
.B1(n_328),
.B2(n_350),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_373),
.A2(n_339),
.B1(n_352),
.B2(n_340),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_376),
.B1(n_401),
.B2(n_399),
.Y(n_489)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_462),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_374),
.Y(n_463)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_398),
.C(n_389),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_465),
.B(n_488),
.C(n_424),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_423),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_466),
.B(n_479),
.Y(n_529)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_467),
.A2(n_472),
.B(n_481),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_419),
.A2(n_373),
.B1(n_374),
.B2(n_408),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_468),
.A2(n_489),
.B1(n_494),
.B2(n_433),
.Y(n_505)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_469),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_470),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_471),
.B(n_473),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_431),
.B(n_378),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_474),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_385),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_475),
.B(n_484),
.Y(n_509)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_476),
.Y(n_511)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_477),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_478),
.A2(n_493),
.B1(n_447),
.B2(n_433),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_432),
.Y(n_479)
);

AO22x1_ASAP7_75t_L g480 ( 
.A1(n_439),
.A2(n_388),
.B1(n_409),
.B2(n_401),
.Y(n_480)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_480),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_427),
.A2(n_402),
.B(n_387),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_398),
.Y(n_482)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_431),
.B(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_483),
.B(n_492),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_394),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_429),
.B(n_405),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_486),
.Y(n_498)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_491),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_440),
.B(n_412),
.C(n_414),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_427),
.A2(n_404),
.B(n_410),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_490),
.A2(n_450),
.B(n_434),
.Y(n_526)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_419),
.A2(n_401),
.B1(n_381),
.B2(n_393),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_428),
.A2(n_382),
.B1(n_413),
.B2(n_397),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_456),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_495),
.B(n_435),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_497),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_500),
.B(n_502),
.Y(n_536)
);

XOR2x2_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_484),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_501),
.B(n_512),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_497),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_505),
.A2(n_507),
.B1(n_518),
.B2(n_520),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_464),
.B(n_449),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_506),
.B(n_333),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_461),
.B(n_446),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_485),
.A2(n_472),
.B1(n_460),
.B2(n_489),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_513),
.A2(n_528),
.B1(n_531),
.B2(n_480),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_461),
.B(n_452),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_517),
.B(n_521),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_485),
.A2(n_430),
.B1(n_458),
.B2(n_454),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_420),
.B1(n_428),
.B2(n_447),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_465),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_524),
.C(n_532),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_424),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g545 ( 
.A(n_525),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_526),
.A2(n_496),
.B(n_413),
.Y(n_554)
);

OAI22x1_ASAP7_75t_SL g528 ( 
.A1(n_460),
.A2(n_422),
.B1(n_435),
.B2(n_445),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_495),
.A2(n_420),
.B1(n_451),
.B2(n_444),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_444),
.C(n_448),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_466),
.A2(n_455),
.B1(n_436),
.B2(n_425),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_533),
.A2(n_474),
.B1(n_425),
.B2(n_413),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_463),
.B(n_333),
.C(n_436),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_492),
.C(n_491),
.Y(n_546)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_499),
.Y(n_537)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_537),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_529),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_540),
.B(n_536),
.Y(n_571)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_529),
.Y(n_541)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_541),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_542),
.A2(n_544),
.B1(n_551),
.B2(n_564),
.Y(n_591)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_510),
.Y(n_543)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_543),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_513),
.A2(n_480),
.B1(n_468),
.B2(n_469),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_546),
.B(n_557),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_514),
.B(n_479),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_547),
.B(n_532),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_494),
.C(n_486),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_548),
.B(n_549),
.C(n_550),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_512),
.B(n_467),
.C(n_481),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_517),
.B(n_487),
.C(n_477),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_528),
.A2(n_490),
.B1(n_496),
.B2(n_476),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_498),
.B(n_462),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_552),
.B(n_558),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_553),
.A2(n_519),
.B1(n_511),
.B2(n_508),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_554),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_524),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_527),
.A2(n_366),
.B(n_351),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_556),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_522),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_391),
.Y(n_558)
);

INVx3_ASAP7_75t_SL g559 ( 
.A(n_504),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_560),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_503),
.B(n_392),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_509),
.B(n_407),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_562),
.B(n_369),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_506),
.B(n_351),
.C(n_366),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_563),
.B(n_501),
.C(n_534),
.Y(n_581)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_515),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_508),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_566),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_527),
.A2(n_470),
.B(n_417),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_470),
.B1(n_438),
.B2(n_396),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_567),
.A2(n_516),
.B1(n_533),
.B2(n_518),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_569),
.A2(n_578),
.B1(n_583),
.B2(n_584),
.Y(n_600)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_542),
.A2(n_507),
.B1(n_523),
.B2(n_505),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_572),
.A2(n_573),
.B1(n_566),
.B2(n_556),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_SL g606 ( 
.A(n_575),
.B(n_539),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_539),
.B(n_530),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_579),
.B(n_589),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_538),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_530),
.C(n_520),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_586),
.C(n_565),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_535),
.A2(n_526),
.B1(n_531),
.B2(n_519),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_541),
.A2(n_511),
.B1(n_516),
.B2(n_504),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_561),
.B(n_369),
.C(n_352),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_552),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_590),
.B(n_592),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_545),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_550),
.B(n_344),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_594),
.B(n_586),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_SL g625 ( 
.A(n_595),
.B(n_612),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_596),
.A2(n_607),
.B1(n_574),
.B2(n_578),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_548),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_597),
.B(n_602),
.Y(n_621)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_577),
.Y(n_599)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_599),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_537),
.Y(n_601)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_601),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_580),
.B(n_562),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_546),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_605),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_593),
.A2(n_551),
.B(n_554),
.Y(n_604)
);

MAJx2_ASAP7_75t_L g628 ( 
.A(n_604),
.B(n_617),
.C(n_570),
.Y(n_628)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_568),
.Y(n_605)
);

XNOR2x1_ASAP7_75t_L g631 ( 
.A(n_606),
.B(n_555),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_591),
.A2(n_553),
.B1(n_549),
.B2(n_544),
.Y(n_607)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_588),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_609),
.B(n_610),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_576),
.B(n_543),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_611),
.B(n_614),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_576),
.B(n_538),
.Y(n_612)
);

OAI21x1_ASAP7_75t_SL g614 ( 
.A1(n_583),
.A2(n_587),
.B(n_585),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_560),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_616),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_593),
.A2(n_567),
.B(n_558),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_600),
.A2(n_587),
.B1(n_573),
.B2(n_585),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_628),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_612),
.B(n_557),
.C(n_579),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_620),
.B(n_627),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_610),
.B(n_581),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_622),
.B(n_631),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_SL g649 ( 
.A1(n_626),
.A2(n_438),
.B1(n_396),
.B2(n_322),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_595),
.B(n_589),
.C(n_572),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_604),
.A2(n_568),
.B(n_584),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_629),
.A2(n_617),
.B(n_615),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_563),
.C(n_575),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_630),
.B(n_344),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_613),
.B(n_606),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_633),
.B(n_634),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_613),
.B(n_588),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_623),
.B(n_598),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_637),
.B(n_647),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_635),
.B(n_601),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_641),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_609),
.Y(n_641)
);

AO21x1_ASAP7_75t_L g654 ( 
.A1(n_642),
.A2(n_643),
.B(n_645),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_629),
.A2(n_607),
.B(n_596),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_624),
.A2(n_608),
.B(n_602),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_621),
.B(n_559),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_648),
.B(n_650),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_649),
.B(n_626),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_621),
.B(n_322),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_618),
.B(n_7),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_651),
.B(n_652),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_9),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_641),
.B(n_619),
.Y(n_656)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_656),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_657),
.B(n_658),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_L g658 ( 
.A(n_646),
.B(n_638),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_639),
.B(n_645),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_660),
.B(n_661),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_642),
.B(n_628),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_644),
.B(n_625),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_663),
.B(n_620),
.Y(n_670)
);

NOR2x1_ASAP7_75t_L g664 ( 
.A(n_643),
.B(n_634),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_664),
.A2(n_627),
.B(n_646),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_654),
.A2(n_644),
.B(n_622),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_668),
.A2(n_669),
.B1(n_670),
.B2(n_662),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_654),
.A2(n_640),
.B(n_633),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_671),
.A2(n_672),
.B(n_658),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_630),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_673),
.A2(n_675),
.B(n_676),
.Y(n_679)
);

AO21x1_ASAP7_75t_L g680 ( 
.A1(n_674),
.A2(n_677),
.B(n_655),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_672),
.B(n_664),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_665),
.B(n_662),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_667),
.A2(n_666),
.B(n_656),
.Y(n_677)
);

NOR2x1_ASAP7_75t_L g678 ( 
.A(n_676),
.B(n_640),
.Y(n_678)
);

AO21x1_ASAP7_75t_L g682 ( 
.A1(n_678),
.A2(n_659),
.B(n_368),
.Y(n_682)
);

MAJx2_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_657),
.C(n_631),
.Y(n_681)
);

BUFx24_ASAP7_75t_SL g683 ( 
.A(n_681),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_683),
.B(n_682),
.Y(n_684)
);

XOR2xp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_679),
.Y(n_685)
);


endmodule