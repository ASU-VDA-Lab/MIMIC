module fake_jpeg_23551_n_172 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_22),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_1),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_22),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_23),
.B1(n_31),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_53),
.B1(n_15),
.B2(n_3),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_23),
.B1(n_35),
.B2(n_30),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_27),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_25),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_28),
.B(n_15),
.C(n_25),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_57),
.B(n_40),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_29),
.C(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_36),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_81),
.C(n_44),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_63),
.B1(n_50),
.B2(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_42),
.B1(n_24),
.B2(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_11),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_74),
.B(n_81),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_36),
.B(n_37),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_82),
.B(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_74),
.Y(n_87)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_50),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_2),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_86),
.B(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_59),
.C(n_50),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_72),
.C(n_78),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_81),
.B(n_65),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_100),
.Y(n_106)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_104),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_65),
.B1(n_72),
.B2(n_76),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_3),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_98),
.B1(n_121),
.B2(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_68),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_109),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_89),
.C(n_100),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_60),
.B1(n_71),
.B2(n_75),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_102),
.B1(n_95),
.B2(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_85),
.C(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_75),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_104),
.B1(n_95),
.B2(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_135),
.C(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_90),
.B(n_86),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_135),
.C(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_119),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_146),
.B1(n_126),
.B2(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_120),
.Y(n_145)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_117),
.A3(n_75),
.B1(n_133),
.B2(n_123),
.C(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_114),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_128),
.A3(n_117),
.B1(n_123),
.B2(n_110),
.C1(n_132),
.C2(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_152),
.B(n_141),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_127),
.B1(n_125),
.B2(n_88),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_88),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_113),
.C(n_134),
.Y(n_153)
);

NOR2xp67_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_117),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_155),
.A2(n_160),
.B(n_101),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_7),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_8),
.B1(n_11),
.B2(n_5),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_143),
.B(n_99),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_153),
.B1(n_143),
.B2(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_164),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_4),
.B(n_5),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_164),
.CI(n_163),
.CON(n_169),
.SN(n_169)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_170),
.B1(n_6),
.B2(n_167),
.C(n_159),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_6),
.B1(n_166),
.B2(n_137),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_170),
.Y(n_172)
);


endmodule