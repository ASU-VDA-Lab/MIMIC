module fake_netlist_1_6411_n_1907 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_407, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_431, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_448, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_383, n_6, n_400, n_296, n_157, n_79, n_202, n_386, n_432, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_389, n_436, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_387, n_163, n_434, n_105, n_227, n_384, n_231, n_298, n_411, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_401, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_443, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_392, n_39, n_279, n_303, n_437, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_447, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_426, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_417, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_393, n_24, n_247, n_381, n_304, n_399, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_402, n_32, n_413, n_391, n_427, n_235, n_243, n_415, n_394, n_442, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_404, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_412, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_430, n_88, n_33, n_107, n_403, n_254, n_262, n_10, n_239, n_439, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_420, n_423, n_342, n_446, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_388, n_193, n_273, n_390, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_416, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_409, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_428, n_75, n_376, n_344, n_136, n_283, n_76, n_435, n_216, n_147, n_148, n_212, n_92, n_11, n_419, n_396, n_168, n_398, n_445, n_438, n_134, n_429, n_233, n_82, n_106, n_440, n_173, n_422, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_449, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_441, n_104, n_74, n_335, n_272, n_146, n_397, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_424, n_156, n_124, n_297, n_128, n_129, n_410, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_418, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_444, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_425, n_332, n_414, n_350, n_433, n_164, n_421, n_175, n_145, n_408, n_290, n_405, n_280, n_21, n_99, n_109, n_132, n_395, n_406, n_151, n_385, n_257, n_269, n_1907, n_1903);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_407;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_431;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_448;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_383;
input n_6;
input n_400;
input n_296;
input n_157;
input n_79;
input n_202;
input n_386;
input n_432;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_389;
input n_436;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_387;
input n_163;
input n_434;
input n_105;
input n_227;
input n_384;
input n_231;
input n_298;
input n_411;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_401;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_443;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_392;
input n_39;
input n_279;
input n_303;
input n_437;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_447;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_426;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_417;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_393;
input n_24;
input n_247;
input n_381;
input n_304;
input n_399;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_402;
input n_32;
input n_413;
input n_391;
input n_427;
input n_235;
input n_243;
input n_415;
input n_394;
input n_442;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_404;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_412;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_430;
input n_88;
input n_33;
input n_107;
input n_403;
input n_254;
input n_262;
input n_10;
input n_239;
input n_439;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_420;
input n_423;
input n_342;
input n_446;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_388;
input n_193;
input n_273;
input n_390;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_416;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_409;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_428;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_435;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_419;
input n_396;
input n_168;
input n_398;
input n_445;
input n_438;
input n_134;
input n_429;
input n_233;
input n_82;
input n_106;
input n_440;
input n_173;
input n_422;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_449;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_441;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_397;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_424;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_410;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_418;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_444;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_425;
input n_332;
input n_414;
input n_350;
input n_433;
input n_164;
input n_421;
input n_175;
input n_145;
input n_408;
input n_290;
input n_405;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_395;
input n_406;
input n_151;
input n_385;
input n_257;
input n_269;
output n_1907;
output n_1903;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_1671;
wire n_646;
wire n_1334;
wire n_1698;
wire n_1627;
wire n_1858;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_1812;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_1785;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_1667;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_1782;
wire n_877;
wire n_1445;
wire n_1663;
wire n_545;
wire n_896;
wire n_588;
wire n_1743;
wire n_1019;
wire n_1714;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_452;
wire n_518;
wire n_1336;
wire n_1341;
wire n_1381;
wire n_1760;
wire n_1884;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1672;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1840;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1906;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_1874;
wire n_979;
wire n_499;
wire n_1683;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_1895;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_950;
wire n_676;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_1744;
wire n_501;
wire n_1898;
wire n_699;
wire n_1654;
wire n_551;
wire n_1061;
wire n_509;
wire n_849;
wire n_1732;
wire n_864;
wire n_1772;
wire n_961;
wire n_1525;
wire n_1718;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1882;
wire n_1500;
wire n_1209;
wire n_1739;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1775;
wire n_1620;
wire n_537;
wire n_1764;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1758;
wire n_1406;
wire n_1789;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_1831;
wire n_556;
wire n_1891;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_1900;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_1707;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_1731;
wire n_1871;
wire n_1902;
wire n_514;
wire n_1693;
wire n_1690;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1877;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1790;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1703;
wire n_1377;
wire n_1079;
wire n_1582;
wire n_1321;
wire n_1801;
wire n_1890;
wire n_1838;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1728;
wire n_1385;
wire n_1711;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1716;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_1193;
wire n_1119;
wire n_825;
wire n_815;
wire n_477;
wire n_1695;
wire n_908;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_1819;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1788;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1682;
wire n_1740;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1826;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_1730;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_1768;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1802;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1694;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_1792;
wire n_753;
wire n_1753;
wire n_658;
wire n_691;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_1893;
wire n_1542;
wire n_1892;
wire n_1311;
wire n_1558;
wire n_483;
wire n_992;
wire n_1748;
wire n_1754;
wire n_1077;
wire n_838;
wire n_705;
wire n_1741;
wire n_964;
wire n_590;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1681;
wire n_1289;
wire n_957;
wire n_808;
wire n_484;
wire n_862;
wire n_852;
wire n_1602;
wire n_1769;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1868;
wire n_1886;
wire n_1202;
wire n_1897;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_1733;
wire n_911;
wire n_980;
wire n_1847;
wire n_1675;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1709;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1852;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_1825;
wire n_973;
wire n_587;
wire n_1818;
wire n_1468;
wire n_476;
wire n_1725;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_1787;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_1829;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1834;
wire n_1670;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_1515;
wire n_897;
wire n_1810;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1807;
wire n_1791;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1861;
wire n_1643;
wire n_1687;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_1854;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_1811;
wire n_767;
wire n_550;
wire n_826;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_478;
wire n_482;
wire n_485;
wire n_1248;
wire n_1828;
wire n_519;
wire n_1465;
wire n_1777;
wire n_1851;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1778;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_1710;
wire n_1781;
wire n_842;
wire n_1269;
wire n_614;
wire n_1346;
wire n_1107;
wire n_799;
wire n_1427;
wire n_1765;
wire n_1050;
wire n_1593;
wire n_1763;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_1844;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1668;
wire n_1692;
wire n_1845;
wire n_1153;
wire n_1797;
wire n_1657;
wire n_1655;
wire n_1771;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_1875;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_1762;
wire n_942;
wire n_1862;
wire n_1029;
wire n_1665;
wire n_508;
wire n_721;
wire n_1060;
wire n_640;
wire n_1766;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_1817;
wire n_811;
wire n_1849;
wire n_530;
wire n_737;
wire n_1696;
wire n_1832;
wire n_1266;
wire n_795;
wire n_1232;
wire n_1796;
wire n_734;
wire n_919;
wire n_763;
wire n_1724;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1752;
wire n_1645;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_1633;
wire n_1784;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1837;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_1894;
wire n_688;
wire n_1800;
wire n_515;
wire n_1577;
wire n_1719;
wire n_1290;
wire n_1813;
wire n_1888;
wire n_1234;
wire n_592;
wire n_1878;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1798;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_1705;
wire n_457;
wire n_1799;
wire n_1757;
wire n_736;
wire n_1495;
wire n_1822;
wire n_1583;
wire n_606;
wire n_1729;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_1697;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_1720;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1679;
wire n_1881;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_1688;
wire n_1767;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1904;
wire n_1554;
wire n_1455;
wire n_659;
wire n_1329;
wire n_1750;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_1896;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1830;
wire n_1101;
wire n_1857;
wire n_1072;
wire n_1761;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_1508;
wire n_1375;
wire n_969;
wire n_1835;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1795;
wire n_1659;
wire n_1816;
wire n_1901;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1734;
wire n_1701;
wire n_1332;
wire n_1480;
wire n_703;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1704;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1870;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_1823;
wire n_546;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1759;
wire n_1774;
wire n_1846;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_516;
wire n_1864;
wire n_1873;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_1794;
wire n_1684;
wire n_1089;
wire n_1717;
wire n_1434;
wire n_1058;
wire n_1396;
wire n_1400;
wire n_1842;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_1706;
wire n_1473;
wire n_1678;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1674;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1755;
wire n_1804;
wire n_1773;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1712;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1779;
wire n_1170;
wire n_1887;
wire n_1523;
wire n_1700;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_1550;
wire n_1827;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1722;
wire n_1872;
wire n_1288;
wire n_1340;
wire n_1903;
wire n_1042;
wire n_1130;
wire n_584;
wire n_1325;
wire n_912;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_1726;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1735;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1689;
wire n_1756;
wire n_1805;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1824;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_1850;
wire n_473;
wire n_1699;
wire n_991;
wire n_1865;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_1713;
wire n_1905;
wire n_913;
wire n_845;
wire n_1776;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_1780;
wire n_934;
wire n_1737;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1749;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_1786;
wire n_757;
wire n_1568;
wire n_750;
wire n_1855;
wire n_645;
wire n_1022;
wire n_1880;
wire n_1856;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_1806;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_1821;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1833;
wire n_1379;
wire n_1003;
wire n_1676;
wire n_678;
wire n_1200;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_1708;
wire n_481;
wire n_694;
wire n_1601;
wire n_1863;
wire n_1262;
wire n_1479;
wire n_1885;
wire n_1486;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_1666;
wire n_1169;
wire n_975;
wire n_1721;
wire n_1081;
wire n_1680;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_1669;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_1815;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1859;
wire n_1673;
wire n_1180;
wire n_647;
wire n_1839;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1742;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1736;
wire n_1245;
wire n_1195;
wire n_1866;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_1876;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1843;
wire n_1076;
wire n_1808;
wire n_1879;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1793;
wire n_1041;
wire n_1745;
wire n_1080;
wire n_1727;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1738;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1809;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_881;
wire n_653;
wire n_1820;
wire n_1853;
wire n_1867;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1814;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_1883;
wire n_861;
wire n_654;
wire n_1221;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_1702;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1685;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_1836;
wire n_1848;
wire n_1285;
wire n_1860;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1677;
wire n_1296;
wire n_1751;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1723;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1783;
wire n_1390;
wire n_1691;
wire n_1715;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1889;
wire n_1487;
wire n_1747;
wire n_1686;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_1770;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_1137;
wire n_1841;
wire n_1869;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_1803;
wire n_1398;
wire n_491;
wire n_1746;
wire n_1291;
INVx1_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_18), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_407), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_292), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_130), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_176), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_373), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_190), .B(n_252), .Y(n_457) );
INVxp33_ASAP7_75t_SL g458 ( .A(n_151), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_83), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_285), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_411), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_440), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_259), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_439), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_87), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_6), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_140), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_15), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_102), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_135), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_116), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_291), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_243), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_189), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_438), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_155), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_207), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_427), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_421), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_372), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_376), .Y(n_481) );
BUFx10_ASAP7_75t_L g482 ( .A(n_77), .Y(n_482) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_130), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_80), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_335), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_310), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_272), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_206), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_131), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_265), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_166), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_64), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_173), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_155), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_33), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_168), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_184), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_225), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_221), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_176), .Y(n_502) );
INVxp33_ASAP7_75t_L g503 ( .A(n_15), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_305), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_63), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_21), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_420), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_288), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_9), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_77), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_172), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_235), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_230), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_331), .Y(n_514) );
INVxp33_ASAP7_75t_L g515 ( .A(n_127), .Y(n_515) );
INVx4_ASAP7_75t_R g516 ( .A(n_446), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_46), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_136), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_201), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_98), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_281), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_181), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_7), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_328), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_114), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_177), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_101), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_256), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_428), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_415), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_14), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_410), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_85), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_21), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_390), .Y(n_535) );
BUFx5_ASAP7_75t_L g536 ( .A(n_356), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_177), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_46), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_398), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_49), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_119), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_228), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_436), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_279), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_419), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_120), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_278), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_208), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_360), .Y(n_549) );
BUFx8_ASAP7_75t_SL g550 ( .A(n_432), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_296), .Y(n_551) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_245), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_445), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_139), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_4), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_391), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_113), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_72), .B(n_11), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_0), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_142), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_129), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_416), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_113), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_413), .Y(n_564) );
CKINVDCx16_ASAP7_75t_R g565 ( .A(n_132), .Y(n_565) );
BUFx3_ASAP7_75t_L g566 ( .A(n_257), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_290), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_39), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_324), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_326), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_267), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_388), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_332), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_111), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_271), .Y(n_575) );
CKINVDCx16_ASAP7_75t_R g576 ( .A(n_145), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_301), .B(n_338), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_270), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_85), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_131), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_94), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_167), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_3), .B(n_375), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_196), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_91), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_280), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_183), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_304), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_128), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_409), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_105), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_447), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_261), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_192), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_95), .Y(n_595) );
BUFx3_ASAP7_75t_L g596 ( .A(n_18), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_402), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_175), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_358), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_263), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_395), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_67), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_57), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_444), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_61), .Y(n_605) );
CKINVDCx16_ASAP7_75t_R g606 ( .A(n_325), .Y(n_606) );
INVxp33_ASAP7_75t_L g607 ( .A(n_64), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_277), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_442), .Y(n_609) );
BUFx3_ASAP7_75t_L g610 ( .A(n_318), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_406), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_369), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_308), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_96), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_340), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_125), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_217), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_254), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_62), .Y(n_619) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_28), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_128), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_4), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_63), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_306), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_70), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_381), .Y(n_626) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_365), .Y(n_627) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_260), .Y(n_628) );
BUFx8_ASAP7_75t_SL g629 ( .A(n_30), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_127), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_213), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_249), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_80), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_101), .Y(n_634) );
INVxp33_ASAP7_75t_L g635 ( .A(n_187), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_392), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_333), .Y(n_637) );
BUFx3_ASAP7_75t_L g638 ( .A(n_53), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_354), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_210), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_12), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_345), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_339), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_156), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_48), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_94), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_307), .Y(n_647) );
INVxp67_ASAP7_75t_SL g648 ( .A(n_366), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_139), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_72), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_274), .Y(n_651) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_23), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_370), .Y(n_653) );
CKINVDCx16_ASAP7_75t_R g654 ( .A(n_321), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_173), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_144), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_6), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_317), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_137), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_312), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_404), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_224), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_170), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_319), .Y(n_664) );
CKINVDCx16_ASAP7_75t_R g665 ( .A(n_253), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_242), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_289), .Y(n_667) );
INVxp33_ASAP7_75t_L g668 ( .A(n_241), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_33), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_313), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_146), .B(n_342), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g672 ( .A(n_329), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_384), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_133), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_377), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_268), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_297), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_505), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_536), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_458), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_458), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_470), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_465), .B(n_5), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_536), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_503), .B(n_5), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_536), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_455), .B(n_7), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_503), .B(n_8), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_515), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_515), .B(n_8), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_607), .B(n_9), .Y(n_691) );
CKINVDCx8_ASAP7_75t_R g692 ( .A(n_552), .Y(n_692) );
INVx6_ASAP7_75t_L g693 ( .A(n_536), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_465), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_607), .B(n_10), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_536), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_502), .B(n_10), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_505), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_536), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_534), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_550), .Y(n_701) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_632), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_534), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_536), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_559), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_502), .B(n_11), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_472), .B(n_12), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_471), .Y(n_708) );
AND2x4_ASAP7_75t_L g709 ( .A(n_596), .B(n_13), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_635), .B(n_13), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_596), .B(n_14), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_635), .B(n_16), .Y(n_712) );
BUFx2_ASAP7_75t_L g713 ( .A(n_669), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_565), .B(n_16), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_638), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_638), .B(n_17), .Y(n_716) );
INVx3_ASAP7_75t_L g717 ( .A(n_645), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_550), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_601), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_689), .B(n_576), .Y(n_720) );
BUFx3_ASAP7_75t_L g721 ( .A(n_694), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_715), .B(n_530), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_715), .B(n_645), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_689), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_708), .B(n_468), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_708), .B(n_668), .Y(n_726) );
AND2x6_ASAP7_75t_L g727 ( .A(n_683), .B(n_479), .Y(n_727) );
INVx2_ASAP7_75t_SL g728 ( .A(n_693), .Y(n_728) );
INVx4_ASAP7_75t_SL g729 ( .A(n_693), .Y(n_729) );
CKINVDCx11_ASAP7_75t_R g730 ( .A(n_682), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_694), .B(n_631), .Y(n_731) );
AO22x2_ASAP7_75t_L g732 ( .A1(n_683), .A2(n_583), .B1(n_483), .B2(n_554), .Y(n_732) );
INVx3_ASAP7_75t_L g733 ( .A(n_683), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_679), .Y(n_734) );
NOR2x1p5_ASAP7_75t_L g735 ( .A(n_701), .B(n_468), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_679), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_694), .B(n_668), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_719), .B(n_613), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_702), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_694), .B(n_453), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_702), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_702), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_679), .Y(n_743) );
INVx1_ASAP7_75t_SL g744 ( .A(n_718), .Y(n_744) );
NOR2xp33_ASAP7_75t_SL g745 ( .A(n_692), .B(n_606), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_713), .B(n_627), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_702), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_684), .Y(n_748) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_687), .A2(n_455), .B1(n_531), .B2(n_495), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_702), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_719), .B(n_654), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_684), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_717), .B(n_453), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_717), .B(n_569), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_719), .B(n_665), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_684), .Y(n_756) );
BUFx4f_ASAP7_75t_L g757 ( .A(n_683), .Y(n_757) );
INVx2_ASAP7_75t_SL g758 ( .A(n_693), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_686), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_721), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_757), .A2(n_706), .B(n_709), .C(n_697), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_737), .B(n_712), .Y(n_762) );
NAND3xp33_ASAP7_75t_SL g763 ( .A(n_744), .B(n_718), .C(n_692), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_721), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_737), .B(n_712), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_723), .B(n_690), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_723), .B(n_690), .Y(n_767) );
NOR2x2_ASAP7_75t_L g768 ( .A(n_730), .B(n_687), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_723), .B(n_713), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_723), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_757), .B(n_692), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_721), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_734), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_757), .A2(n_697), .B1(n_709), .B2(n_706), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_738), .B(n_722), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_734), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_726), .B(n_685), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_732), .A2(n_706), .B1(n_709), .B2(n_697), .Y(n_778) );
BUFx3_ASAP7_75t_L g779 ( .A(n_727), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_732), .A2(n_706), .B1(n_709), .B2(n_697), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_757), .A2(n_716), .B(n_711), .C(n_696), .Y(n_781) );
NAND2x1_ASAP7_75t_L g782 ( .A(n_727), .B(n_693), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_L g783 ( .A1(n_724), .A2(n_688), .B(n_691), .C(n_685), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_731), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_726), .B(n_688), .Y(n_785) );
INVx4_ASAP7_75t_L g786 ( .A(n_727), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_722), .B(n_707), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_725), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_732), .A2(n_716), .B1(n_711), .B2(n_695), .Y(n_789) );
INVx8_ASAP7_75t_L g790 ( .A(n_727), .Y(n_790) );
INVx8_ASAP7_75t_L g791 ( .A(n_727), .Y(n_791) );
INVx2_ASAP7_75t_SL g792 ( .A(n_725), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_727), .A2(n_711), .B1(n_716), .B2(n_693), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_751), .B(n_691), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_731), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_736), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_720), .A2(n_714), .B1(n_681), .B2(n_680), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g798 ( .A(n_733), .B(n_711), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_746), .B(n_714), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g800 ( .A(n_733), .B(n_716), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_736), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_727), .B(n_695), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_727), .B(n_710), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_733), .Y(n_804) );
NOR2x1p5_ASAP7_75t_L g805 ( .A(n_720), .B(n_710), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_746), .B(n_717), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g807 ( .A(n_733), .B(n_686), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_740), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_743), .B(n_686), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_755), .B(n_678), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_732), .A2(n_553), .B1(n_570), .B2(n_512), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_732), .A2(n_696), .B1(n_704), .B2(n_699), .Y(n_812) );
AND2x4_ASAP7_75t_SL g813 ( .A(n_745), .B(n_512), .Y(n_813) );
AND2x2_ASAP7_75t_SL g814 ( .A(n_745), .B(n_672), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_740), .Y(n_815) );
NAND2x1p5_ASAP7_75t_L g816 ( .A(n_744), .B(n_680), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_729), .B(n_473), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_743), .B(n_717), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_753), .B(n_678), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_735), .B(n_482), .Y(n_820) );
AND2x6_ASAP7_75t_SL g821 ( .A(n_749), .B(n_451), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_749), .B(n_520), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_748), .B(n_473), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_748), .B(n_681), .C(n_603), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_752), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_752), .B(n_475), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_756), .B(n_475), .Y(n_827) );
INVx4_ASAP7_75t_L g828 ( .A(n_729), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_756), .B(n_481), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_735), .A2(n_553), .B1(n_593), .B2(n_570), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_759), .B(n_481), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_753), .B(n_698), .Y(n_832) );
NAND2xp5_ASAP7_75t_SL g833 ( .A(n_729), .B(n_487), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_759), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_754), .B(n_482), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_754), .B(n_698), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_728), .B(n_758), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_728), .A2(n_696), .B1(n_704), .B2(n_699), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_729), .Y(n_839) );
INVx4_ASAP7_75t_L g840 ( .A(n_729), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_758), .B(n_487), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g842 ( .A(n_739), .B(n_699), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g843 ( .A(n_750), .B(n_521), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_739), .B(n_561), .C(n_541), .Y(n_844) );
NOR2x1_ASAP7_75t_L g845 ( .A(n_763), .B(n_593), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_770), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_808), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_799), .B(n_495), .Y(n_848) );
NOR3xp33_ASAP7_75t_SL g849 ( .A(n_797), .B(n_603), .C(n_520), .Y(n_849) );
AND2x4_ASAP7_75t_L g850 ( .A(n_835), .B(n_784), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_813), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_792), .B(n_629), .Y(n_852) );
O2A1O1Ixp33_ASAP7_75t_L g853 ( .A1(n_761), .A2(n_703), .B(n_705), .C(n_700), .Y(n_853) );
NAND2xp5_ASAP7_75t_SL g854 ( .A(n_786), .B(n_521), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_778), .A2(n_662), .B1(n_600), .B2(n_555), .Y(n_855) );
BUFx12f_ASAP7_75t_L g856 ( .A(n_821), .Y(n_856) );
OR2x6_ASAP7_75t_SL g857 ( .A(n_822), .B(n_619), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_762), .B(n_619), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_815), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_765), .B(n_630), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_834), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_807), .A2(n_704), .B(n_671), .Y(n_862) );
AO32x1_ASAP7_75t_L g863 ( .A1(n_773), .A2(n_456), .A3(n_461), .B1(n_460), .B2(n_450), .Y(n_863) );
OAI21xp33_ASAP7_75t_L g864 ( .A1(n_775), .A2(n_630), .B(n_496), .Y(n_864) );
NOR2xp33_ASAP7_75t_SL g865 ( .A(n_786), .B(n_600), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_807), .A2(n_508), .B(n_452), .Y(n_866) );
CKINVDCx16_ASAP7_75t_R g867 ( .A(n_788), .Y(n_867) );
INVxp67_ASAP7_75t_L g868 ( .A(n_777), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g869 ( .A(n_779), .B(n_535), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_775), .A2(n_459), .B(n_467), .C(n_466), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_834), .Y(n_871) );
O2A1O1Ixp33_ASAP7_75t_L g872 ( .A1(n_781), .A2(n_703), .B(n_705), .C(n_700), .Y(n_872) );
O2A1O1Ixp33_ASAP7_75t_L g873 ( .A1(n_783), .A2(n_469), .B(n_484), .C(n_476), .Y(n_873) );
O2A1O1Ixp5_ASAP7_75t_L g874 ( .A1(n_787), .A2(n_628), .B(n_648), .C(n_519), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_804), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_804), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_795), .Y(n_877) );
OR2x6_ASAP7_75t_SL g878 ( .A(n_768), .B(n_535), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_773), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_780), .A2(n_662), .B1(n_555), .B2(n_574), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_776), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_776), .Y(n_882) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_812), .B(n_499), .C(n_493), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_794), .B(n_580), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_813), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_785), .B(n_649), .Y(n_886) );
A2O1A1Ixp33_ASAP7_75t_L g887 ( .A1(n_789), .A2(n_494), .B(n_498), .C(n_497), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_812), .A2(n_558), .B1(n_574), .B2(n_531), .Y(n_888) );
OAI22x1_ASAP7_75t_L g889 ( .A1(n_811), .A2(n_587), .B1(n_629), .B2(n_568), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_830), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_796), .Y(n_891) );
NOR2xp67_ASAP7_75t_SL g892 ( .A(n_779), .B(n_543), .Y(n_892) );
BUFx6f_ASAP7_75t_L g893 ( .A(n_790), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_766), .B(n_581), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_796), .Y(n_895) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_824), .B(n_620), .C(n_454), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_767), .B(n_633), .Y(n_897) );
NAND2xp5_ASAP7_75t_SL g898 ( .A(n_793), .B(n_543), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_774), .A2(n_587), .B1(n_578), .B2(n_564), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_769), .B(n_656), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_787), .B(n_652), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_801), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_805), .B(n_564), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_819), .B(n_578), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_801), .Y(n_905) );
INVx3_ASAP7_75t_L g906 ( .A(n_790), .Y(n_906) );
O2A1O1Ixp33_ASAP7_75t_L g907 ( .A1(n_806), .A2(n_509), .B(n_510), .C(n_506), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_819), .B(n_594), .Y(n_908) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_798), .A2(n_464), .B(n_462), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_816), .B(n_579), .Y(n_910) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_832), .Y(n_911) );
INVx3_ASAP7_75t_L g912 ( .A(n_790), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_832), .B(n_594), .Y(n_913) );
BUFx3_ASAP7_75t_L g914 ( .A(n_825), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_836), .B(n_597), .Y(n_915) );
NAND2xp5_ASAP7_75t_SL g916 ( .A(n_793), .B(n_597), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g917 ( .A1(n_774), .A2(n_517), .B(n_518), .C(n_511), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_836), .B(n_599), .Y(n_918) );
NAND3xp33_ASAP7_75t_SL g919 ( .A(n_816), .B(n_585), .C(n_599), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_825), .Y(n_920) );
NOR3xp33_ASAP7_75t_SL g921 ( .A(n_810), .B(n_612), .C(n_604), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_820), .B(n_522), .Y(n_922) );
OAI21xp33_ASAP7_75t_SL g923 ( .A1(n_814), .A2(n_525), .B(n_523), .Y(n_923) );
BUFx2_ASAP7_75t_L g924 ( .A(n_814), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_771), .B(n_482), .Y(n_925) );
OAI22x1_ASAP7_75t_L g926 ( .A1(n_810), .A2(n_612), .B1(n_615), .B2(n_604), .Y(n_926) );
OAI21xp33_ASAP7_75t_L g927 ( .A1(n_802), .A2(n_527), .B(n_526), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_844), .A2(n_533), .B1(n_538), .B2(n_537), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_803), .B(n_540), .Y(n_929) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_782), .Y(n_930) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_823), .Y(n_931) );
OAI21xp33_ASAP7_75t_L g932 ( .A1(n_826), .A2(n_557), .B(n_546), .Y(n_932) );
NOR3xp33_ASAP7_75t_SL g933 ( .A(n_841), .B(n_618), .C(n_615), .Y(n_933) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_827), .Y(n_934) );
BUFx2_ASAP7_75t_L g935 ( .A(n_791), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_798), .A2(n_477), .B(n_474), .Y(n_936) );
NAND2xp5_ASAP7_75t_SL g937 ( .A(n_791), .B(n_618), .Y(n_937) );
OAI22xp5_ASAP7_75t_SL g938 ( .A1(n_829), .A2(n_626), .B1(n_560), .B2(n_582), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_831), .B(n_800), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_800), .B(n_563), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_818), .Y(n_941) );
NAND2xp33_ASAP7_75t_SL g942 ( .A(n_791), .B(n_626), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_760), .Y(n_943) );
NOR2xp33_ASAP7_75t_R g944 ( .A(n_837), .B(n_463), .Y(n_944) );
AOI21xp5_ASAP7_75t_L g945 ( .A1(n_809), .A2(n_480), .B(n_478), .Y(n_945) );
BUFx2_ASAP7_75t_SL g946 ( .A(n_828), .Y(n_946) );
INVx1_ASAP7_75t_SL g947 ( .A(n_843), .Y(n_947) );
OAI21x1_ASAP7_75t_L g948 ( .A1(n_842), .A2(n_457), .B(n_739), .Y(n_948) );
INVxp67_ASAP7_75t_SL g949 ( .A(n_760), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_764), .B(n_589), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_764), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_772), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_772), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_838), .B(n_591), .Y(n_954) );
O2A1O1Ixp33_ASAP7_75t_L g955 ( .A1(n_809), .A2(n_602), .B(n_605), .C(n_598), .Y(n_955) );
BUFx2_ASAP7_75t_L g956 ( .A(n_828), .Y(n_956) );
NOR2xp33_ASAP7_75t_R g957 ( .A(n_839), .B(n_507), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_838), .Y(n_958) );
NAND3xp33_ASAP7_75t_SL g959 ( .A(n_817), .B(n_514), .C(n_513), .Y(n_959) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_833), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_842), .A2(n_486), .B(n_485), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g962 ( .A(n_840), .B(n_616), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_840), .Y(n_963) );
NAND2xp5_ASAP7_75t_SL g964 ( .A(n_786), .B(n_528), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_788), .B(n_621), .Y(n_965) );
AOI21xp5_ASAP7_75t_L g966 ( .A1(n_807), .A2(n_489), .B(n_488), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_807), .A2(n_492), .B(n_490), .Y(n_967) );
NOR2xp33_ASAP7_75t_R g968 ( .A(n_763), .B(n_549), .Y(n_968) );
NAND2x2_ASAP7_75t_L g969 ( .A(n_805), .B(n_479), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_799), .B(n_622), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_762), .B(n_623), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_805), .A2(n_641), .B1(n_644), .B2(n_625), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_762), .B(n_650), .Y(n_973) );
A2O1A1Ixp33_ASAP7_75t_L g974 ( .A1(n_775), .A2(n_663), .B(n_674), .C(n_657), .Y(n_974) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_813), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g976 ( .A(n_786), .B(n_551), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_778), .A2(n_559), .B1(n_634), .B2(n_595), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_770), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_807), .A2(n_501), .B(n_500), .Y(n_979) );
INVxp67_ASAP7_75t_L g980 ( .A(n_788), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g981 ( .A1(n_807), .A2(n_524), .B(n_504), .Y(n_981) );
BUFx6f_ASAP7_75t_L g982 ( .A(n_790), .Y(n_982) );
NAND2xp5_ASAP7_75t_SL g983 ( .A(n_786), .B(n_556), .Y(n_983) );
AOI21xp5_ASAP7_75t_L g984 ( .A1(n_807), .A2(n_532), .B(n_529), .Y(n_984) );
O2A1O1Ixp33_ASAP7_75t_L g985 ( .A1(n_761), .A2(n_634), .B(n_646), .C(n_595), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_770), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_770), .Y(n_987) );
BUFx3_ASAP7_75t_L g988 ( .A(n_851), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_877), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_939), .A2(n_542), .B(n_539), .Y(n_990) );
NOR4xp25_ASAP7_75t_L g991 ( .A(n_923), .B(n_659), .C(n_646), .D(n_545), .Y(n_991) );
OR2x6_ASAP7_75t_L g992 ( .A(n_855), .B(n_659), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_865), .A2(n_677), .B1(n_544), .B2(n_548), .Y(n_993) );
BUFx12f_ASAP7_75t_L g994 ( .A(n_885), .Y(n_994) );
AND2x4_ASAP7_75t_L g995 ( .A(n_850), .B(n_547), .Y(n_995) );
AO31x2_ASAP7_75t_L g996 ( .A1(n_977), .A2(n_590), .A3(n_647), .B(n_569), .Y(n_996) );
A2O1A1Ixp33_ASAP7_75t_L g997 ( .A1(n_985), .A2(n_572), .B(n_575), .C(n_567), .Y(n_997) );
AOI21xp5_ASAP7_75t_L g998 ( .A1(n_862), .A2(n_586), .B(n_584), .Y(n_998) );
INVx6_ASAP7_75t_L g999 ( .A(n_969), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_847), .Y(n_1000) );
BUFx6f_ASAP7_75t_L g1001 ( .A(n_893), .Y(n_1001) );
O2A1O1Ixp33_ASAP7_75t_L g1002 ( .A1(n_870), .A2(n_588), .B(n_608), .C(n_592), .Y(n_1002) );
NAND3xp33_ASAP7_75t_L g1003 ( .A(n_849), .B(n_614), .C(n_491), .Y(n_1003) );
AOI21xp5_ASAP7_75t_L g1004 ( .A1(n_862), .A2(n_611), .B(n_609), .Y(n_1004) );
INVxp67_ASAP7_75t_SL g1005 ( .A(n_914), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_911), .B(n_491), .Y(n_1006) );
OAI211xp5_ASAP7_75t_L g1007 ( .A1(n_873), .A2(n_624), .B(n_636), .C(n_617), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g1008 ( .A(n_893), .Y(n_1008) );
BUFx6f_ASAP7_75t_L g1009 ( .A(n_893), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_881), .A2(n_639), .B(n_637), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_867), .B(n_17), .Y(n_1011) );
A2O1A1Ixp33_ASAP7_75t_L g1012 ( .A1(n_985), .A2(n_640), .B(n_651), .C(n_642), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_868), .B(n_491), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_859), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_850), .A2(n_614), .B1(n_655), .B2(n_491), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_980), .B(n_614), .Y(n_1016) );
OAI21x1_ASAP7_75t_L g1017 ( .A1(n_948), .A2(n_647), .B(n_590), .Y(n_1017) );
AO31x2_ASAP7_75t_L g1018 ( .A1(n_887), .A2(n_653), .A3(n_660), .B(n_658), .Y(n_1018) );
OAI22x1_ASAP7_75t_L g1019 ( .A1(n_924), .A2(n_667), .B1(n_670), .B2(n_666), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_879), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_950), .Y(n_1021) );
AO32x2_ASAP7_75t_L g1022 ( .A1(n_938), .A2(n_702), .A3(n_655), .B1(n_614), .B2(n_516), .Y(n_1022) );
AOI221x1_ASAP7_75t_L g1023 ( .A1(n_919), .A2(n_676), .B1(n_673), .B2(n_632), .C(n_655), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_880), .B(n_19), .Y(n_1024) );
AO21x2_ASAP7_75t_L g1025 ( .A1(n_961), .A2(n_577), .B(n_741), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g1026 ( .A1(n_882), .A2(n_750), .B(n_742), .Y(n_1026) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_891), .A2(n_750), .B(n_742), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_848), .A2(n_571), .B1(n_573), .B2(n_562), .Y(n_1028) );
O2A1O1Ixp33_ASAP7_75t_L g1029 ( .A1(n_974), .A2(n_610), .B(n_566), .C(n_741), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_846), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_975), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g1032 ( .A1(n_873), .A2(n_655), .B(n_610), .C(n_566), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_888), .A2(n_643), .B1(n_664), .B2(n_661), .Y(n_1033) );
AOI21xp5_ASAP7_75t_L g1034 ( .A1(n_895), .A2(n_747), .B(n_742), .Y(n_1034) );
OA21x2_ASAP7_75t_L g1035 ( .A1(n_961), .A2(n_747), .B(n_741), .Y(n_1035) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_878), .Y(n_1036) );
INVx3_ASAP7_75t_L g1037 ( .A(n_922), .Y(n_1037) );
A2O1A1Ixp33_ASAP7_75t_L g1038 ( .A1(n_853), .A2(n_632), .B(n_675), .C(n_747), .Y(n_1038) );
O2A1O1Ixp33_ASAP7_75t_SL g1039 ( .A1(n_853), .A2(n_191), .B(n_193), .C(n_188), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_902), .Y(n_1040) );
AND2x4_ASAP7_75t_L g1041 ( .A(n_931), .B(n_19), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_917), .B(n_20), .Y(n_1042) );
OAI21xp5_ASAP7_75t_L g1043 ( .A1(n_874), .A2(n_195), .B(n_194), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_909), .A2(n_198), .B(n_197), .Y(n_1044) );
AO31x2_ASAP7_75t_L g1045 ( .A1(n_958), .A2(n_23), .A3(n_20), .B(n_22), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_978), .Y(n_1046) );
AOI21xp5_ASAP7_75t_L g1047 ( .A1(n_905), .A2(n_200), .B(n_199), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_899), .Y(n_1048) );
OA21x2_ASAP7_75t_L g1049 ( .A1(n_945), .A2(n_203), .B(n_202), .Y(n_1049) );
INVx3_ASAP7_75t_L g1050 ( .A(n_922), .Y(n_1050) );
BUFx8_ASAP7_75t_SL g1051 ( .A(n_856), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g1052 ( .A(n_982), .Y(n_1052) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_852), .B(n_890), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_889), .A2(n_25), .B1(n_22), .B2(n_24), .Y(n_1054) );
INVx1_ASAP7_75t_SL g1055 ( .A(n_910), .Y(n_1055) );
A2O1A1Ixp33_ASAP7_75t_L g1056 ( .A1(n_872), .A2(n_26), .B(n_24), .C(n_25), .Y(n_1056) );
AO31x2_ASAP7_75t_L g1057 ( .A1(n_929), .A2(n_28), .A3(n_26), .B(n_27), .Y(n_1057) );
OAI21xp5_ASAP7_75t_L g1058 ( .A1(n_909), .A2(n_205), .B(n_204), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_857), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_903), .B(n_27), .Y(n_1060) );
AOI21xp5_ASAP7_75t_L g1061 ( .A1(n_920), .A2(n_211), .B(n_209), .Y(n_1061) );
O2A1O1Ixp33_ASAP7_75t_L g1062 ( .A1(n_907), .A2(n_901), .B(n_955), .C(n_896), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_934), .B(n_29), .Y(n_1063) );
A2O1A1Ixp33_ASAP7_75t_L g1064 ( .A1(n_955), .A2(n_31), .B(n_29), .C(n_30), .Y(n_1064) );
NAND2x1_ASAP7_75t_L g1065 ( .A(n_861), .B(n_212), .Y(n_1065) );
INVx1_ASAP7_75t_SL g1066 ( .A(n_965), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_858), .B(n_31), .Y(n_1067) );
O2A1O1Ixp33_ASAP7_75t_SL g1068 ( .A1(n_964), .A2(n_215), .B(n_216), .C(n_214), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_860), .B(n_32), .Y(n_1069) );
O2A1O1Ixp33_ASAP7_75t_L g1070 ( .A1(n_907), .A2(n_35), .B(n_32), .C(n_34), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_900), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_1071) );
BUFx10_ASAP7_75t_L g1072 ( .A(n_940), .Y(n_1072) );
AO31x2_ASAP7_75t_L g1073 ( .A1(n_936), .A2(n_38), .A3(n_36), .B(n_37), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_864), .A2(n_39), .B1(n_37), .B2(n_38), .Y(n_1074) );
AO32x2_ASAP7_75t_L g1075 ( .A1(n_863), .A2(n_40), .A3(n_41), .B1(n_42), .B2(n_43), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_970), .B(n_40), .Y(n_1076) );
AO31x2_ASAP7_75t_L g1077 ( .A1(n_936), .A2(n_43), .A3(n_41), .B(n_42), .Y(n_1077) );
BUFx10_ASAP7_75t_L g1078 ( .A(n_962), .Y(n_1078) );
AND2x4_ASAP7_75t_L g1079 ( .A(n_935), .B(n_44), .Y(n_1079) );
AO32x2_ASAP7_75t_L g1080 ( .A1(n_863), .A2(n_44), .A3(n_45), .B1(n_47), .B2(n_48), .Y(n_1080) );
AO31x2_ASAP7_75t_L g1081 ( .A1(n_945), .A2(n_49), .A3(n_45), .B(n_47), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_898), .A2(n_52), .B1(n_50), .B2(n_51), .Y(n_1082) );
AO32x2_ASAP7_75t_L g1083 ( .A1(n_863), .A2(n_50), .A3(n_51), .B1(n_52), .B2(n_53), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_906), .B(n_54), .Y(n_1084) );
AO21x1_ASAP7_75t_L g1085 ( .A1(n_966), .A2(n_219), .B(n_218), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_916), .A2(n_56), .B1(n_54), .B2(n_55), .Y(n_1086) );
AOI21xp5_ASAP7_75t_L g1087 ( .A1(n_871), .A2(n_222), .B(n_220), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_884), .B(n_55), .Y(n_1088) );
A2O1A1Ixp33_ASAP7_75t_L g1089 ( .A1(n_932), .A2(n_58), .B(n_56), .C(n_57), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_944), .Y(n_1090) );
NOR2xp33_ASAP7_75t_L g1091 ( .A(n_886), .B(n_58), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_951), .Y(n_1092) );
AOI21xp5_ASAP7_75t_L g1093 ( .A1(n_949), .A2(n_226), .B(n_223), .Y(n_1093) );
A2O1A1Ixp33_ASAP7_75t_L g1094 ( .A1(n_966), .A2(n_61), .B(n_59), .C(n_60), .Y(n_1094) );
AOI21xp5_ASAP7_75t_L g1095 ( .A1(n_854), .A2(n_229), .B(n_227), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_986), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_845), .A2(n_62), .B1(n_59), .B2(n_60), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_941), .A2(n_67), .B1(n_65), .B2(n_66), .Y(n_1098) );
INVx1_ASAP7_75t_SL g1099 ( .A(n_926), .Y(n_1099) );
INVx3_ASAP7_75t_L g1100 ( .A(n_982), .Y(n_1100) );
O2A1O1Ixp33_ASAP7_75t_L g1101 ( .A1(n_971), .A2(n_68), .B(n_65), .C(n_66), .Y(n_1101) );
INVxp67_ASAP7_75t_L g1102 ( .A(n_904), .Y(n_1102) );
INVx2_ASAP7_75t_L g1103 ( .A(n_953), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_943), .Y(n_1104) );
INVx3_ASAP7_75t_L g1105 ( .A(n_982), .Y(n_1105) );
BUFx10_ASAP7_75t_L g1106 ( .A(n_925), .Y(n_1106) );
O2A1O1Ixp33_ASAP7_75t_L g1107 ( .A1(n_973), .A2(n_70), .B(n_68), .C(n_69), .Y(n_1107) );
A2O1A1Ixp33_ASAP7_75t_L g1108 ( .A1(n_967), .A2(n_73), .B(n_69), .C(n_71), .Y(n_1108) );
INVx1_ASAP7_75t_SL g1109 ( .A(n_947), .Y(n_1109) );
O2A1O1Ixp33_ASAP7_75t_L g1110 ( .A1(n_894), .A2(n_74), .B(n_71), .C(n_73), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_957), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_972), .B(n_74), .Y(n_1112) );
AOI21xp5_ASAP7_75t_L g1113 ( .A1(n_908), .A2(n_232), .B(n_231), .Y(n_1113) );
INVx3_ASAP7_75t_L g1114 ( .A(n_875), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_987), .Y(n_1115) );
OAI21x1_ASAP7_75t_L g1116 ( .A1(n_967), .A2(n_234), .B(n_233), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_913), .A2(n_918), .B(n_915), .Y(n_1117) );
AOI221xp5_ASAP7_75t_L g1118 ( .A1(n_928), .A2(n_897), .B1(n_954), .B2(n_927), .C(n_921), .Y(n_1118) );
NOR2xp67_ASAP7_75t_SL g1119 ( .A(n_946), .B(n_75), .Y(n_1119) );
OAI22x1_ASAP7_75t_L g1120 ( .A1(n_883), .A2(n_78), .B1(n_75), .B2(n_76), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_976), .A2(n_237), .B(n_236), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_952), .A2(n_79), .B1(n_76), .B2(n_78), .Y(n_1122) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_983), .A2(n_239), .B(n_238), .Y(n_1123) );
O2A1O1Ixp33_ASAP7_75t_SL g1124 ( .A1(n_960), .A2(n_244), .B(n_246), .C(n_240), .Y(n_1124) );
AOI21xp5_ASAP7_75t_L g1125 ( .A1(n_979), .A2(n_248), .B(n_247), .Y(n_1125) );
NOR2xp33_ASAP7_75t_L g1126 ( .A(n_876), .B(n_79), .Y(n_1126) );
OAI21x1_ASAP7_75t_L g1127 ( .A1(n_979), .A2(n_251), .B(n_250), .Y(n_1127) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_981), .A2(n_258), .B(n_255), .Y(n_1128) );
AO31x2_ASAP7_75t_L g1129 ( .A1(n_984), .A2(n_83), .A3(n_81), .B(n_82), .Y(n_1129) );
AO32x2_ASAP7_75t_L g1130 ( .A1(n_984), .A2(n_933), .A3(n_866), .B1(n_968), .B2(n_942), .Y(n_1130) );
AOI21xp5_ASAP7_75t_L g1131 ( .A1(n_869), .A2(n_264), .B(n_262), .Y(n_1131) );
CKINVDCx8_ASAP7_75t_R g1132 ( .A(n_956), .Y(n_1132) );
AO31x2_ASAP7_75t_L g1133 ( .A1(n_866), .A2(n_81), .A3(n_82), .B(n_84), .Y(n_1133) );
A2O1A1Ixp33_ASAP7_75t_L g1134 ( .A1(n_930), .A2(n_84), .B(n_86), .C(n_87), .Y(n_1134) );
A2O1A1Ixp33_ASAP7_75t_L g1135 ( .A1(n_906), .A2(n_86), .B(n_88), .C(n_89), .Y(n_1135) );
INVx2_ASAP7_75t_L g1136 ( .A(n_963), .Y(n_1136) );
NAND2x1p5_ASAP7_75t_L g1137 ( .A(n_912), .B(n_88), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_912), .B(n_89), .Y(n_1138) );
O2A1O1Ixp33_ASAP7_75t_L g1139 ( .A1(n_937), .A2(n_90), .B(n_91), .C(n_92), .Y(n_1139) );
OAI22x1_ASAP7_75t_L g1140 ( .A1(n_892), .A2(n_90), .B1(n_92), .B2(n_93), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_959), .Y(n_1141) );
INVx2_ASAP7_75t_L g1142 ( .A(n_847), .Y(n_1142) );
A2O1A1Ixp33_ASAP7_75t_L g1143 ( .A1(n_939), .A2(n_93), .B(n_95), .C(n_96), .Y(n_1143) );
BUFx6f_ASAP7_75t_L g1144 ( .A(n_893), .Y(n_1144) );
OAI21xp5_ASAP7_75t_L g1145 ( .A1(n_939), .A2(n_269), .B(n_266), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_867), .B(n_97), .Y(n_1146) );
A2O1A1Ixp33_ASAP7_75t_L g1147 ( .A1(n_939), .A2(n_97), .B(n_98), .C(n_99), .Y(n_1147) );
AOI21xp33_ASAP7_75t_L g1148 ( .A1(n_852), .A2(n_99), .B(n_100), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_867), .B(n_100), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1150 ( .A(n_867), .B(n_102), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g1151 ( .A(n_865), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_911), .B(n_103), .Y(n_1152) );
INVx3_ASAP7_75t_L g1153 ( .A(n_850), .Y(n_1153) );
A2O1A1Ixp33_ASAP7_75t_L g1154 ( .A1(n_939), .A2(n_103), .B(n_104), .C(n_105), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_877), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_877), .Y(n_1156) );
OR2x6_ASAP7_75t_L g1157 ( .A(n_855), .B(n_104), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_877), .Y(n_1158) );
OAI21xp5_ASAP7_75t_L g1159 ( .A1(n_939), .A2(n_275), .B(n_273), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_877), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_877), .Y(n_1161) );
O2A1O1Ixp33_ASAP7_75t_SL g1162 ( .A1(n_881), .A2(n_295), .B(n_448), .C(n_443), .Y(n_1162) );
A2O1A1Ixp33_ASAP7_75t_L g1163 ( .A1(n_939), .A2(n_106), .B(n_107), .C(n_108), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_867), .B(n_106), .Y(n_1164) );
AOI21xp5_ASAP7_75t_L g1165 ( .A1(n_939), .A2(n_282), .B(n_276), .Y(n_1165) );
AOI21xp5_ASAP7_75t_L g1166 ( .A1(n_1117), .A2(n_284), .B(n_283), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1066), .B(n_107), .Y(n_1167) );
AO21x2_ASAP7_75t_L g1168 ( .A1(n_1043), .A2(n_287), .B(n_286), .Y(n_1168) );
AOI21x1_ASAP7_75t_L g1169 ( .A1(n_1017), .A2(n_294), .B(n_293), .Y(n_1169) );
AOI21xp5_ASAP7_75t_L g1170 ( .A1(n_1039), .A2(n_299), .B(n_298), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_1157), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_1171) );
AOI21xp5_ASAP7_75t_L g1172 ( .A1(n_998), .A2(n_302), .B(n_300), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_989), .Y(n_1173) );
OAI21xp33_ASAP7_75t_L g1174 ( .A1(n_991), .A2(n_109), .B(n_110), .Y(n_1174) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_1051), .Y(n_1175) );
INVxp67_ASAP7_75t_L g1176 ( .A(n_1041), .Y(n_1176) );
AO31x2_ASAP7_75t_L g1177 ( .A1(n_1085), .A2(n_111), .A3(n_112), .B(n_114), .Y(n_1177) );
AOI22xp33_ASAP7_75t_SL g1178 ( .A1(n_1157), .A2(n_112), .B1(n_115), .B2(n_116), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1000), .B(n_115), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1155), .B(n_117), .Y(n_1180) );
AOI21xp5_ASAP7_75t_L g1181 ( .A1(n_1004), .A2(n_309), .B(n_303), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_1014), .B(n_117), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_988), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_992), .A2(n_118), .B1(n_119), .B2(n_120), .Y(n_1184) );
AOI21xp33_ASAP7_75t_SL g1185 ( .A1(n_1036), .A2(n_118), .B(n_121), .Y(n_1185) );
INVx2_ASAP7_75t_SL g1186 ( .A(n_999), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1156), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1158), .Y(n_1188) );
INVx3_ASAP7_75t_L g1189 ( .A(n_1008), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1160), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1055), .B(n_121), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1161), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1142), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1102), .B(n_122), .Y(n_1194) );
BUFx3_ASAP7_75t_L g1195 ( .A(n_994), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_1153), .B(n_1115), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1048), .B(n_122), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_992), .B(n_123), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1030), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1046), .Y(n_1200) );
OAI21xp5_ASAP7_75t_L g1201 ( .A1(n_997), .A2(n_123), .B(n_124), .Y(n_1201) );
OR2x6_ASAP7_75t_L g1202 ( .A(n_1079), .B(n_124), .Y(n_1202) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_999), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g1204 ( .A1(n_1035), .A2(n_330), .B(n_441), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1041), .B(n_125), .Y(n_1205) );
A2O1A1Ixp33_ASAP7_75t_L g1206 ( .A1(n_1062), .A2(n_126), .B(n_129), .C(n_132), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1096), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1076), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_993), .A2(n_126), .B1(n_133), .B2(n_134), .Y(n_1209) );
OAI21x1_ASAP7_75t_L g1210 ( .A1(n_1035), .A2(n_336), .B(n_437), .Y(n_1210) );
BUFx2_ASAP7_75t_L g1211 ( .A(n_1031), .Y(n_1211) );
AOI21xp5_ASAP7_75t_L g1212 ( .A1(n_1118), .A2(n_334), .B(n_435), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1006), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1091), .B(n_134), .Y(n_1214) );
AOI21xp5_ASAP7_75t_L g1215 ( .A1(n_1038), .A2(n_337), .B(n_434), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_1151), .A2(n_135), .B1(n_136), .B2(n_137), .Y(n_1216) );
AOI21xp5_ASAP7_75t_L g1217 ( .A1(n_990), .A2(n_341), .B(n_433), .Y(n_1217) );
AOI221xp5_ASAP7_75t_L g1218 ( .A1(n_1002), .A2(n_138), .B1(n_140), .B2(n_141), .C(n_142), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1021), .B(n_138), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1024), .B(n_141), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_1079), .Y(n_1221) );
OA21x2_ASAP7_75t_L g1222 ( .A1(n_1023), .A2(n_344), .B(n_431), .Y(n_1222) );
AO21x2_ASAP7_75t_L g1223 ( .A1(n_1145), .A2(n_343), .B(n_429), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1037), .B(n_143), .Y(n_1224) );
AOI21x1_ASAP7_75t_L g1225 ( .A1(n_1049), .A2(n_327), .B(n_426), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1013), .Y(n_1226) );
A2O1A1Ixp33_ASAP7_75t_L g1227 ( .A1(n_1060), .A2(n_143), .B(n_144), .C(n_145), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1152), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1104), .Y(n_1229) );
INVx6_ASAP7_75t_L g1230 ( .A(n_1106), .Y(n_1230) );
INVxp67_ASAP7_75t_SL g1231 ( .A(n_1005), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1232 ( .A(n_1050), .Y(n_1232) );
BUFx6f_ASAP7_75t_L g1233 ( .A(n_1001), .Y(n_1233) );
OA21x2_ASAP7_75t_L g1234 ( .A1(n_1159), .A2(n_347), .B(n_424), .Y(n_1234) );
AOI21xp5_ASAP7_75t_L g1235 ( .A1(n_1067), .A2(n_346), .B(n_423), .Y(n_1235) );
AOI21xp5_ASAP7_75t_L g1236 ( .A1(n_1069), .A2(n_323), .B(n_422), .Y(n_1236) );
AOI21xp33_ASAP7_75t_L g1237 ( .A1(n_1029), .A2(n_146), .B(n_147), .Y(n_1237) );
HB1xp67_ASAP7_75t_L g1238 ( .A(n_1132), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1088), .B(n_147), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1084), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1084), .B(n_148), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1020), .Y(n_1242) );
OAI221xp5_ASAP7_75t_L g1243 ( .A1(n_1053), .A2(n_148), .B1(n_149), .B2(n_150), .C(n_151), .Y(n_1243) );
AOI21x1_ASAP7_75t_L g1244 ( .A1(n_1049), .A2(n_349), .B(n_418), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_995), .B(n_149), .Y(n_1245) );
A2O1A1Ixp33_ASAP7_75t_L g1246 ( .A1(n_1070), .A2(n_150), .B(n_152), .C(n_153), .Y(n_1246) );
BUFx6f_ASAP7_75t_L g1247 ( .A(n_1001), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1138), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1109), .B(n_152), .Y(n_1249) );
A2O1A1Ixp33_ASAP7_75t_L g1250 ( .A1(n_1003), .A2(n_153), .B(n_154), .C(n_156), .Y(n_1250) );
OAI21xp33_ASAP7_75t_SL g1251 ( .A1(n_1044), .A2(n_154), .B(n_157), .Y(n_1251) );
A2O1A1Ixp33_ASAP7_75t_L g1252 ( .A1(n_1110), .A2(n_157), .B(n_158), .C(n_159), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1138), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1040), .Y(n_1254) );
OAI221xp5_ASAP7_75t_L g1255 ( .A1(n_1059), .A2(n_158), .B1(n_159), .B2(n_160), .C(n_161), .Y(n_1255) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1092), .Y(n_1256) );
NOR4xp25_ASAP7_75t_L g1257 ( .A(n_1007), .B(n_160), .C(n_161), .D(n_162), .Y(n_1257) );
BUFx10_ASAP7_75t_L g1258 ( .A(n_1090), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1137), .Y(n_1259) );
AOI21xp5_ASAP7_75t_L g1260 ( .A1(n_1025), .A2(n_355), .B(n_417), .Y(n_1260) );
AOI222xp33_ASAP7_75t_L g1261 ( .A1(n_1164), .A2(n_162), .B1(n_163), .B2(n_164), .C1(n_165), .C2(n_166), .Y(n_1261) );
OA21x2_ASAP7_75t_L g1262 ( .A1(n_1058), .A2(n_357), .B(n_414), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1133), .Y(n_1263) );
AOI21xp5_ASAP7_75t_L g1264 ( .A1(n_1026), .A2(n_353), .B(n_412), .Y(n_1264) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_1027), .A2(n_352), .B(n_408), .Y(n_1265) );
AOI21xp5_ASAP7_75t_L g1266 ( .A1(n_1034), .A2(n_351), .B(n_405), .Y(n_1266) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1103), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1072), .B(n_163), .Y(n_1268) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1073), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1133), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1078), .Y(n_1271) );
AOI21xp5_ASAP7_75t_L g1272 ( .A1(n_1113), .A2(n_359), .B(n_403), .Y(n_1272) );
NOR3xp33_ASAP7_75t_L g1273 ( .A(n_1148), .B(n_164), .C(n_165), .Y(n_1273) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_1111), .Y(n_1274) );
OAI21x1_ASAP7_75t_L g1275 ( .A1(n_1116), .A2(n_361), .B(n_401), .Y(n_1275) );
HB1xp67_ASAP7_75t_L g1276 ( .A(n_1136), .Y(n_1276) );
AND2x4_ASAP7_75t_SL g1277 ( .A(n_1008), .B(n_167), .Y(n_1277) );
A2O1A1Ixp33_ASAP7_75t_L g1278 ( .A1(n_1139), .A2(n_168), .B(n_169), .C(n_170), .Y(n_1278) );
AOI21xp5_ASAP7_75t_L g1279 ( .A1(n_1124), .A2(n_362), .B(n_400), .Y(n_1279) );
AND2x4_ASAP7_75t_L g1280 ( .A(n_1001), .B(n_169), .Y(n_1280) );
NAND2x1_ASAP7_75t_L g1281 ( .A(n_1052), .B(n_363), .Y(n_1281) );
AOI21xp5_ASAP7_75t_L g1282 ( .A1(n_1162), .A2(n_350), .B(n_399), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_995), .B(n_171), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1112), .B(n_171), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1033), .B(n_172), .Y(n_1285) );
AOI21xp5_ASAP7_75t_L g1286 ( .A1(n_1165), .A2(n_364), .B(n_397), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1073), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_1052), .B(n_174), .Y(n_1288) );
AO31x2_ASAP7_75t_L g1289 ( .A1(n_1012), .A2(n_1120), .A3(n_1056), .B(n_1089), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_1063), .A2(n_174), .B1(n_175), .B2(n_178), .Y(n_1290) );
A2O1A1Ixp33_ASAP7_75t_L g1291 ( .A1(n_1101), .A2(n_178), .B(n_179), .C(n_180), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1122), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1099), .B(n_179), .Y(n_1293) );
AND2x4_ASAP7_75t_L g1294 ( .A(n_1052), .B(n_180), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1011), .B(n_181), .Y(n_1295) );
OR2x4_ASAP7_75t_L g1296 ( .A(n_1146), .B(n_182), .Y(n_1296) );
OR2x6_ASAP7_75t_L g1297 ( .A(n_1149), .B(n_182), .Y(n_1297) );
OA21x2_ASAP7_75t_L g1298 ( .A1(n_1128), .A2(n_371), .B(n_394), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1119), .Y(n_1299) );
OAI21x1_ASAP7_75t_L g1300 ( .A1(n_1127), .A2(n_368), .B(n_393), .Y(n_1300) );
AO21x2_ASAP7_75t_L g1301 ( .A1(n_1032), .A2(n_367), .B(n_389), .Y(n_1301) );
OAI21xp5_ASAP7_75t_L g1302 ( .A1(n_1042), .A2(n_183), .B(n_184), .Y(n_1302) );
AOI21xp5_ASAP7_75t_L g1303 ( .A1(n_1068), .A2(n_374), .B(n_387), .Y(n_1303) );
INVx2_ASAP7_75t_L g1304 ( .A(n_1077), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1077), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1019), .B(n_185), .Y(n_1306) );
AOI21xp33_ASAP7_75t_L g1307 ( .A1(n_1141), .A2(n_185), .B(n_186), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1077), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1016), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_1126), .A2(n_186), .B1(n_187), .B2(n_311), .Y(n_1310) );
AO31x2_ASAP7_75t_L g1311 ( .A1(n_1064), .A2(n_314), .A3(n_315), .B(n_316), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1028), .B(n_320), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1010), .B(n_322), .Y(n_1313) );
OA21x2_ASAP7_75t_L g1314 ( .A1(n_1093), .A2(n_348), .B(n_378), .Y(n_1314) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1150), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1018), .B(n_449), .Y(n_1316) );
A2O1A1Ixp33_ASAP7_75t_L g1317 ( .A1(n_1107), .A2(n_379), .B(n_380), .C(n_382), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1081), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_1054), .A2(n_383), .B1(n_385), .B2(n_386), .Y(n_1319) );
AO31x2_ASAP7_75t_L g1320 ( .A1(n_1143), .A2(n_1163), .A3(n_1154), .B(n_1147), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1081), .Y(n_1321) );
A2O1A1Ixp33_ASAP7_75t_L g1322 ( .A1(n_1094), .A2(n_1108), .B(n_1135), .C(n_1134), .Y(n_1322) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1129), .Y(n_1323) );
OAI21x1_ASAP7_75t_L g1324 ( .A1(n_1065), .A2(n_1047), .B(n_1061), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1018), .B(n_1114), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1081), .Y(n_1326) );
BUFx6f_ASAP7_75t_L g1327 ( .A(n_1144), .Y(n_1327) );
BUFx3_ASAP7_75t_L g1328 ( .A(n_1009), .Y(n_1328) );
AOI22xp33_ASAP7_75t_SL g1329 ( .A1(n_1144), .A2(n_1009), .B1(n_1105), .B2(n_1100), .Y(n_1329) );
AOI21x1_ASAP7_75t_L g1330 ( .A1(n_1121), .A2(n_1123), .B(n_1095), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1018), .B(n_1071), .Y(n_1331) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_1144), .A2(n_1140), .B1(n_1130), .B2(n_1125), .Y(n_1332) );
OAI21xp5_ASAP7_75t_L g1333 ( .A1(n_1131), .A2(n_1087), .B(n_1082), .Y(n_1333) );
AND2x6_ASAP7_75t_L g1334 ( .A(n_1130), .B(n_1022), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1129), .Y(n_1335) );
AOI21xp5_ASAP7_75t_L g1336 ( .A1(n_1015), .A2(n_1086), .B(n_1074), .Y(n_1336) );
A2O1A1Ixp33_ASAP7_75t_L g1337 ( .A1(n_1097), .A2(n_1098), .B(n_1130), .C(n_1022), .Y(n_1337) );
AOI21xp5_ASAP7_75t_L g1338 ( .A1(n_996), .A2(n_1022), .B(n_1075), .Y(n_1338) );
BUFx12f_ASAP7_75t_L g1339 ( .A(n_1057), .Y(n_1339) );
OAI21x1_ASAP7_75t_L g1340 ( .A1(n_996), .A2(n_1045), .B(n_1129), .Y(n_1340) );
OAI21x1_ASAP7_75t_L g1341 ( .A1(n_996), .A2(n_1045), .B(n_1075), .Y(n_1341) );
INVxp67_ASAP7_75t_L g1342 ( .A(n_1057), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1057), .Y(n_1343) );
OAI21x1_ASAP7_75t_L g1344 ( .A1(n_1045), .A2(n_1083), .B(n_1075), .Y(n_1344) );
AOI21xp5_ASAP7_75t_L g1345 ( .A1(n_1080), .A2(n_1117), .B(n_1017), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1080), .Y(n_1346) );
OAI221xp5_ASAP7_75t_L g1347 ( .A1(n_1080), .A2(n_849), .B1(n_816), .B2(n_1102), .C(n_923), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1173), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1202), .B(n_1083), .Y(n_1349) );
NAND3xp33_ASAP7_75t_L g1350 ( .A(n_1273), .B(n_1178), .C(n_1343), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1202), .B(n_1276), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1187), .Y(n_1352) );
BUFx3_ASAP7_75t_L g1353 ( .A(n_1328), .Y(n_1353) );
INVx1_ASAP7_75t_SL g1354 ( .A(n_1230), .Y(n_1354) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1287), .Y(n_1355) );
AO21x2_ASAP7_75t_L g1356 ( .A1(n_1345), .A2(n_1338), .B(n_1340), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1325), .Y(n_1357) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1304), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1188), .Y(n_1359) );
INVx3_ASAP7_75t_L g1360 ( .A(n_1233), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1190), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1362 ( .A(n_1233), .B(n_1247), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1192), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1199), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1200), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1202), .B(n_1229), .Y(n_1366) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1323), .Y(n_1367) );
INVx3_ASAP7_75t_L g1368 ( .A(n_1233), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1242), .B(n_1254), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1207), .B(n_1220), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1193), .B(n_1167), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1182), .Y(n_1372) );
INVx3_ASAP7_75t_L g1373 ( .A(n_1247), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1182), .Y(n_1374) );
OAI22xp33_ASAP7_75t_L g1375 ( .A1(n_1171), .A2(n_1221), .B1(n_1297), .B2(n_1347), .Y(n_1375) );
OR2x6_ASAP7_75t_L g1376 ( .A(n_1241), .B(n_1297), .Y(n_1376) );
OA21x2_ASAP7_75t_L g1377 ( .A1(n_1341), .A2(n_1344), .B(n_1308), .Y(n_1377) );
OR2x6_ASAP7_75t_L g1378 ( .A(n_1241), .B(n_1297), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1208), .B(n_1292), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1179), .Y(n_1380) );
OAI21xp5_ASAP7_75t_L g1381 ( .A1(n_1336), .A2(n_1322), .B(n_1251), .Y(n_1381) );
INVx2_ASAP7_75t_SL g1382 ( .A(n_1230), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1228), .B(n_1315), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1205), .B(n_1261), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1176), .B(n_1196), .Y(n_1385) );
INVx1_ASAP7_75t_SL g1386 ( .A(n_1271), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1180), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1256), .Y(n_1388) );
AO31x2_ASAP7_75t_L g1389 ( .A1(n_1305), .A2(n_1335), .A3(n_1318), .B(n_1326), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1261), .B(n_1295), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1267), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1219), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1196), .B(n_1240), .Y(n_1393) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_1247), .Y(n_1394) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1191), .B(n_1198), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1302), .B(n_1231), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1224), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_1171), .A2(n_1243), .B1(n_1174), .B2(n_1201), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1248), .B(n_1253), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1306), .Y(n_1400) );
OR2x6_ASAP7_75t_L g1401 ( .A(n_1259), .B(n_1280), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1194), .Y(n_1402) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1210), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1299), .Y(n_1404) );
AOI22xp33_ASAP7_75t_SL g1405 ( .A1(n_1251), .A2(n_1201), .B1(n_1277), .B2(n_1339), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1245), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1283), .Y(n_1407) );
HB1xp67_ASAP7_75t_L g1408 ( .A(n_1327), .Y(n_1408) );
AND2x4_ASAP7_75t_SL g1409 ( .A(n_1258), .B(n_1238), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1280), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1411 ( .A(n_1211), .B(n_1232), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1302), .B(n_1321), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1263), .B(n_1270), .Y(n_1413) );
HB1xp67_ASAP7_75t_L g1414 ( .A(n_1327), .Y(n_1414) );
INVx2_ASAP7_75t_L g1415 ( .A(n_1346), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1288), .Y(n_1416) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1169), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1288), .Y(n_1418) );
INVx2_ASAP7_75t_SL g1419 ( .A(n_1327), .Y(n_1419) );
OR2x6_ASAP7_75t_L g1420 ( .A(n_1294), .B(n_1274), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1249), .B(n_1183), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1294), .Y(n_1422) );
OA21x2_ASAP7_75t_L g1423 ( .A1(n_1342), .A2(n_1337), .B(n_1331), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1257), .B(n_1177), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1197), .Y(n_1425) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1225), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1268), .B(n_1184), .Y(n_1427) );
OR2x6_ASAP7_75t_L g1428 ( .A(n_1195), .B(n_1189), .Y(n_1428) );
BUFx3_ASAP7_75t_L g1429 ( .A(n_1189), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1293), .Y(n_1430) );
AND2x4_ASAP7_75t_L g1431 ( .A(n_1213), .B(n_1309), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1257), .B(n_1177), .Y(n_1432) );
HB1xp67_ASAP7_75t_L g1433 ( .A(n_1334), .Y(n_1433) );
OA21x2_ASAP7_75t_L g1434 ( .A1(n_1174), .A2(n_1316), .B(n_1170), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1290), .Y(n_1435) );
AOI22xp5_ASAP7_75t_L g1436 ( .A1(n_1209), .A2(n_1214), .B1(n_1285), .B2(n_1312), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1216), .Y(n_1437) );
AO21x2_ASAP7_75t_L g1438 ( .A1(n_1244), .A2(n_1279), .B(n_1237), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1177), .B(n_1320), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1320), .B(n_1289), .Y(n_1440) );
AOI21xp33_ASAP7_75t_L g1441 ( .A1(n_1239), .A2(n_1284), .B(n_1226), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1296), .Y(n_1442) );
AO21x2_ASAP7_75t_L g1443 ( .A1(n_1168), .A2(n_1282), .B(n_1260), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1227), .B(n_1255), .Y(n_1444) );
BUFx6f_ASAP7_75t_L g1445 ( .A(n_1281), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1320), .B(n_1289), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1185), .B(n_1307), .Y(n_1447) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1206), .Y(n_1448) );
BUFx3_ASAP7_75t_L g1449 ( .A(n_1186), .Y(n_1449) );
HB1xp67_ASAP7_75t_L g1450 ( .A(n_1334), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1185), .Y(n_1451) );
NOR2xp33_ASAP7_75t_L g1452 ( .A(n_1246), .B(n_1203), .Y(n_1452) );
BUFx2_ASAP7_75t_L g1453 ( .A(n_1334), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1289), .B(n_1332), .Y(n_1454) );
INVx3_ASAP7_75t_L g1455 ( .A(n_1275), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1311), .B(n_1291), .Y(n_1456) );
OR2x6_ASAP7_75t_L g1457 ( .A(n_1212), .B(n_1166), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1218), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1252), .Y(n_1459) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1310), .B(n_1278), .Y(n_1460) );
AND2x4_ASAP7_75t_L g1461 ( .A(n_1311), .B(n_1300), .Y(n_1461) );
BUFx3_ASAP7_75t_L g1462 ( .A(n_1258), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1329), .B(n_1175), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1250), .Y(n_1464) );
AOI21xp5_ASAP7_75t_SL g1465 ( .A1(n_1234), .A2(n_1262), .B(n_1298), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1313), .B(n_1311), .Y(n_1466) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1222), .Y(n_1467) );
OR2x6_ASAP7_75t_L g1468 ( .A(n_1286), .B(n_1217), .Y(n_1468) );
INVx2_ASAP7_75t_SL g1469 ( .A(n_1223), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1334), .B(n_1333), .Y(n_1470) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1262), .Y(n_1471) );
OA21x2_ASAP7_75t_L g1472 ( .A1(n_1204), .A2(n_1324), .B(n_1333), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1172), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1181), .Y(n_1474) );
HB1xp67_ASAP7_75t_L g1475 ( .A(n_1223), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1235), .Y(n_1476) );
INVx2_ASAP7_75t_L g1477 ( .A(n_1298), .Y(n_1477) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1317), .B(n_1319), .Y(n_1478) );
OAI22xp5_ASAP7_75t_L g1479 ( .A1(n_1215), .A2(n_1236), .B1(n_1272), .B2(n_1314), .Y(n_1479) );
OAI31xp33_ASAP7_75t_L g1480 ( .A1(n_1264), .A2(n_1265), .A3(n_1266), .B(n_1303), .Y(n_1480) );
AO21x2_ASAP7_75t_L g1481 ( .A1(n_1168), .A2(n_1301), .B(n_1330), .Y(n_1481) );
INVx2_ASAP7_75t_L g1482 ( .A(n_1269), .Y(n_1482) );
BUFx2_ASAP7_75t_L g1483 ( .A(n_1231), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1202), .B(n_1066), .Y(n_1484) );
OA21x2_ASAP7_75t_L g1485 ( .A1(n_1340), .A2(n_1341), .B(n_1344), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1202), .B(n_1066), .Y(n_1486) );
OR2x6_ASAP7_75t_L g1487 ( .A(n_1202), .B(n_1241), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1202), .B(n_1055), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1173), .Y(n_1489) );
HB1xp67_ASAP7_75t_L g1490 ( .A(n_1325), .Y(n_1490) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1173), .Y(n_1491) );
BUFx3_ASAP7_75t_L g1492 ( .A(n_1328), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1173), .Y(n_1493) );
HB1xp67_ASAP7_75t_L g1494 ( .A(n_1325), .Y(n_1494) );
INVx5_ASAP7_75t_SL g1495 ( .A(n_1202), .Y(n_1495) );
HB1xp67_ASAP7_75t_L g1496 ( .A(n_1325), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1202), .B(n_1055), .Y(n_1497) );
HB1xp67_ASAP7_75t_L g1498 ( .A(n_1325), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1202), .B(n_1066), .Y(n_1499) );
NOR2xp33_ASAP7_75t_L g1500 ( .A(n_1176), .B(n_867), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1242), .B(n_1254), .Y(n_1501) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1269), .Y(n_1502) );
OR2x2_ASAP7_75t_L g1503 ( .A(n_1483), .B(n_1357), .Y(n_1503) );
OR2x6_ASAP7_75t_L g1504 ( .A(n_1487), .B(n_1376), .Y(n_1504) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1348), .Y(n_1505) );
BUFx3_ASAP7_75t_L g1506 ( .A(n_1353), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1357), .B(n_1490), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1440), .B(n_1446), .Y(n_1508) );
HB1xp67_ASAP7_75t_L g1509 ( .A(n_1431), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1352), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1359), .Y(n_1511) );
HB1xp67_ASAP7_75t_L g1512 ( .A(n_1431), .Y(n_1512) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1413), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1440), .B(n_1446), .Y(n_1514) );
HB1xp67_ASAP7_75t_L g1515 ( .A(n_1431), .Y(n_1515) );
INVx2_ASAP7_75t_SL g1516 ( .A(n_1362), .Y(n_1516) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1413), .Y(n_1517) );
AND2x4_ASAP7_75t_L g1518 ( .A(n_1470), .B(n_1433), .Y(n_1518) );
OR2x2_ASAP7_75t_L g1519 ( .A(n_1490), .B(n_1494), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1470), .B(n_1439), .Y(n_1520) );
OR2x2_ASAP7_75t_L g1521 ( .A(n_1494), .B(n_1496), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1415), .Y(n_1522) );
INVxp67_ASAP7_75t_L g1523 ( .A(n_1500), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1439), .B(n_1412), .Y(n_1524) );
INVx3_ASAP7_75t_L g1525 ( .A(n_1362), .Y(n_1525) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1361), .Y(n_1526) );
AND2x4_ASAP7_75t_L g1527 ( .A(n_1433), .B(n_1450), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1363), .B(n_1364), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1412), .B(n_1454), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1454), .B(n_1369), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1369), .B(n_1501), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1365), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1501), .B(n_1496), .Y(n_1533) );
INVx1_ASAP7_75t_SL g1534 ( .A(n_1354), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1498), .B(n_1423), .Y(n_1535) );
INVx2_ASAP7_75t_SL g1536 ( .A(n_1362), .Y(n_1536) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1489), .Y(n_1537) );
HB1xp67_ASAP7_75t_L g1538 ( .A(n_1487), .Y(n_1538) );
BUFx2_ASAP7_75t_L g1539 ( .A(n_1498), .Y(n_1539) );
HB1xp67_ASAP7_75t_L g1540 ( .A(n_1487), .Y(n_1540) );
INVxp67_ASAP7_75t_SL g1541 ( .A(n_1394), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1423), .B(n_1424), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1423), .B(n_1424), .Y(n_1543) );
AOI221x1_ASAP7_75t_L g1544 ( .A1(n_1451), .A2(n_1350), .B1(n_1441), .B2(n_1432), .C(n_1465), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1432), .B(n_1450), .Y(n_1545) );
INVxp67_ASAP7_75t_L g1546 ( .A(n_1500), .Y(n_1546) );
AND2x4_ASAP7_75t_L g1547 ( .A(n_1453), .B(n_1415), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1381), .B(n_1491), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1493), .B(n_1389), .Y(n_1549) );
NOR2xp33_ASAP7_75t_L g1550 ( .A(n_1386), .B(n_1376), .Y(n_1550) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1388), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1389), .B(n_1396), .Y(n_1552) );
AOI21xp33_ASAP7_75t_SL g1553 ( .A1(n_1376), .A2(n_1378), .B(n_1375), .Y(n_1553) );
OAI221xp5_ASAP7_75t_L g1554 ( .A1(n_1400), .A2(n_1452), .B1(n_1436), .B2(n_1442), .C(n_1378), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1391), .Y(n_1555) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1355), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1389), .B(n_1396), .Y(n_1557) );
AOI33xp33_ASAP7_75t_L g1558 ( .A1(n_1430), .A2(n_1390), .A3(n_1425), .B1(n_1384), .B2(n_1402), .B3(n_1404), .Y(n_1558) );
AOI22xp5_ASAP7_75t_L g1559 ( .A1(n_1427), .A2(n_1452), .B1(n_1375), .B2(n_1378), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1389), .B(n_1349), .Y(n_1560) );
BUFx6f_ASAP7_75t_L g1561 ( .A(n_1445), .Y(n_1561) );
INVx2_ASAP7_75t_L g1562 ( .A(n_1358), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1358), .B(n_1367), .Y(n_1563) );
NAND2xp5_ASAP7_75t_L g1564 ( .A(n_1379), .B(n_1370), .Y(n_1564) );
AOI22xp5_ASAP7_75t_L g1565 ( .A1(n_1458), .A2(n_1447), .B1(n_1435), .B2(n_1495), .Y(n_1565) );
NAND2xp5_ASAP7_75t_SL g1566 ( .A(n_1495), .B(n_1405), .Y(n_1566) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1383), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1482), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1406), .B(n_1407), .Y(n_1569) );
NOR2xp67_ASAP7_75t_L g1570 ( .A(n_1382), .B(n_1462), .Y(n_1570) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1502), .Y(n_1571) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_1437), .A2(n_1444), .B1(n_1495), .B2(n_1398), .Y(n_1572) );
HB1xp67_ASAP7_75t_L g1573 ( .A(n_1411), .Y(n_1573) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1377), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1371), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1377), .B(n_1456), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1377), .B(n_1456), .Y(n_1577) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1366), .Y(n_1578) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1395), .B(n_1397), .Y(n_1579) );
INVx2_ASAP7_75t_SL g1580 ( .A(n_1394), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_1380), .B(n_1387), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1420), .B(n_1372), .Y(n_1582) );
NOR2xp67_ASAP7_75t_L g1583 ( .A(n_1382), .B(n_1462), .Y(n_1583) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1399), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1485), .B(n_1356), .Y(n_1585) );
INVx2_ASAP7_75t_L g1586 ( .A(n_1356), .Y(n_1586) );
NAND2x1_ASAP7_75t_L g1587 ( .A(n_1465), .B(n_1455), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1374), .B(n_1408), .Y(n_1588) );
INVx1_ASAP7_75t_SL g1589 ( .A(n_1409), .Y(n_1589) );
NAND4xp25_ASAP7_75t_L g1590 ( .A(n_1398), .B(n_1497), .C(n_1488), .D(n_1499), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1408), .B(n_1414), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1414), .B(n_1392), .Y(n_1592) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1420), .B(n_1401), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1410), .B(n_1422), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1420), .B(n_1401), .Y(n_1595) );
HB1xp67_ASAP7_75t_L g1596 ( .A(n_1351), .Y(n_1596) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_1460), .A2(n_1448), .B1(n_1459), .B2(n_1486), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1416), .B(n_1418), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1461), .B(n_1466), .Y(n_1599) );
OR2x6_ASAP7_75t_L g1600 ( .A(n_1401), .B(n_1461), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1601 ( .A(n_1484), .B(n_1393), .Y(n_1601) );
BUFx2_ASAP7_75t_SL g1602 ( .A(n_1353), .Y(n_1602) );
INVxp67_ASAP7_75t_SL g1603 ( .A(n_1360), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1421), .B(n_1385), .Y(n_1604) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1429), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1360), .B(n_1368), .Y(n_1606) );
INVxp67_ASAP7_75t_L g1607 ( .A(n_1492), .Y(n_1607) );
BUFx2_ASAP7_75t_L g1608 ( .A(n_1368), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1368), .B(n_1373), .Y(n_1609) );
AND4x1_ASAP7_75t_L g1610 ( .A(n_1463), .B(n_1409), .C(n_1478), .D(n_1480), .Y(n_1610) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1429), .Y(n_1611) );
AND2x4_ASAP7_75t_L g1612 ( .A(n_1373), .B(n_1419), .Y(n_1612) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1522), .Y(n_1613) );
NAND2x1p5_ASAP7_75t_L g1614 ( .A(n_1570), .B(n_1373), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1529), .B(n_1475), .Y(n_1615) );
INVx3_ASAP7_75t_L g1616 ( .A(n_1561), .Y(n_1616) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1522), .Y(n_1617) );
HB1xp67_ASAP7_75t_L g1618 ( .A(n_1503), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1529), .B(n_1508), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1503), .B(n_1475), .Y(n_1620) );
HB1xp67_ASAP7_75t_L g1621 ( .A(n_1539), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1508), .B(n_1469), .Y(n_1622) );
INVx2_ASAP7_75t_L g1623 ( .A(n_1574), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1514), .B(n_1469), .Y(n_1624) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1568), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1626 ( .A(n_1531), .B(n_1492), .Y(n_1626) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1568), .Y(n_1627) );
BUFx3_ASAP7_75t_L g1628 ( .A(n_1506), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1524), .B(n_1477), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1524), .B(n_1471), .Y(n_1630) );
OR2x6_ASAP7_75t_L g1631 ( .A(n_1600), .B(n_1471), .Y(n_1631) );
OR2x2_ASAP7_75t_L g1632 ( .A(n_1507), .B(n_1519), .Y(n_1632) );
INVx3_ASAP7_75t_L g1633 ( .A(n_1561), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1520), .B(n_1472), .Y(n_1634) );
NOR3xp33_ASAP7_75t_L g1635 ( .A(n_1554), .B(n_1449), .C(n_1478), .Y(n_1635) );
HB1xp67_ASAP7_75t_L g1636 ( .A(n_1539), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1520), .B(n_1472), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1530), .B(n_1472), .Y(n_1638) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1571), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1531), .B(n_1449), .Y(n_1640) );
OR2x6_ASAP7_75t_L g1641 ( .A(n_1600), .B(n_1467), .Y(n_1641) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1519), .B(n_1419), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1571), .Y(n_1643) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1549), .Y(n_1644) );
AND2x4_ASAP7_75t_L g1645 ( .A(n_1599), .B(n_1455), .Y(n_1645) );
AND2x4_ASAP7_75t_L g1646 ( .A(n_1599), .B(n_1455), .Y(n_1646) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1542), .B(n_1481), .Y(n_1647) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1549), .Y(n_1648) );
HB1xp67_ASAP7_75t_L g1649 ( .A(n_1521), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1543), .B(n_1464), .Y(n_1650) );
OR2x2_ASAP7_75t_L g1651 ( .A(n_1521), .B(n_1428), .Y(n_1651) );
OR2x2_ASAP7_75t_L g1652 ( .A(n_1513), .B(n_1428), .Y(n_1652) );
AND2x4_ASAP7_75t_SL g1653 ( .A(n_1504), .B(n_1428), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1552), .B(n_1474), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1655 ( .A(n_1567), .B(n_1473), .Y(n_1655) );
OR2x2_ASAP7_75t_L g1656 ( .A(n_1513), .B(n_1476), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1657 ( .A(n_1552), .B(n_1434), .Y(n_1657) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1517), .Y(n_1658) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1517), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1557), .B(n_1434), .Y(n_1660) );
OR2x2_ASAP7_75t_L g1661 ( .A(n_1557), .B(n_1426), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1560), .B(n_1434), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1560), .B(n_1403), .Y(n_1663) );
NOR2xp33_ASAP7_75t_L g1664 ( .A(n_1534), .B(n_1468), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1576), .B(n_1417), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1666 ( .A(n_1575), .B(n_1468), .Y(n_1666) );
INVx2_ASAP7_75t_SL g1667 ( .A(n_1580), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1576), .B(n_1468), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1533), .B(n_1438), .Y(n_1669) );
AND2x4_ASAP7_75t_L g1670 ( .A(n_1577), .B(n_1445), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1577), .B(n_1443), .Y(n_1671) );
OR2x2_ASAP7_75t_L g1672 ( .A(n_1533), .B(n_1457), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1545), .B(n_1443), .Y(n_1673) );
OR2x2_ASAP7_75t_L g1674 ( .A(n_1545), .B(n_1518), .Y(n_1674) );
OAI22xp5_ASAP7_75t_L g1675 ( .A1(n_1559), .A2(n_1457), .B1(n_1445), .B2(n_1479), .Y(n_1675) );
NAND2x1_ASAP7_75t_L g1676 ( .A(n_1600), .B(n_1445), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1518), .B(n_1438), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1579), .B(n_1457), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1518), .B(n_1548), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1548), .B(n_1563), .Y(n_1680) );
AOI211xp5_ASAP7_75t_L g1681 ( .A1(n_1553), .A2(n_1566), .B(n_1583), .C(n_1590), .Y(n_1681) );
CKINVDCx5p33_ASAP7_75t_R g1682 ( .A(n_1602), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1563), .B(n_1547), .Y(n_1683) );
BUFx2_ASAP7_75t_L g1684 ( .A(n_1600), .Y(n_1684) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1579), .B(n_1564), .Y(n_1685) );
NAND3xp33_ASAP7_75t_L g1686 ( .A(n_1544), .B(n_1610), .C(n_1572), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1687 ( .A(n_1619), .B(n_1632), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1619), .B(n_1535), .Y(n_1688) );
AND2x4_ASAP7_75t_L g1689 ( .A(n_1684), .B(n_1527), .Y(n_1689) );
OR2x2_ASAP7_75t_L g1690 ( .A(n_1632), .B(n_1573), .Y(n_1690) );
OR2x6_ASAP7_75t_L g1691 ( .A(n_1631), .B(n_1504), .Y(n_1691) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1649), .Y(n_1692) );
NAND2xp5_ASAP7_75t_L g1693 ( .A(n_1618), .B(n_1558), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1683), .B(n_1596), .Y(n_1694) );
NOR2x1_ASAP7_75t_SL g1695 ( .A(n_1628), .B(n_1504), .Y(n_1695) );
OR2x2_ASAP7_75t_L g1696 ( .A(n_1674), .B(n_1601), .Y(n_1696) );
INVx2_ASAP7_75t_L g1697 ( .A(n_1623), .Y(n_1697) );
AND2x4_ASAP7_75t_L g1698 ( .A(n_1684), .B(n_1527), .Y(n_1698) );
NAND2xp5_ASAP7_75t_L g1699 ( .A(n_1650), .B(n_1592), .Y(n_1699) );
AOI22xp33_ASAP7_75t_SL g1700 ( .A1(n_1653), .A2(n_1504), .B1(n_1538), .B2(n_1540), .Y(n_1700) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1658), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1650), .B(n_1680), .Y(n_1702) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1658), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1704 ( .A(n_1680), .B(n_1592), .Y(n_1704) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1659), .Y(n_1705) );
NOR2xp33_ASAP7_75t_L g1706 ( .A(n_1626), .B(n_1565), .Y(n_1706) );
NAND2xp5_ASAP7_75t_L g1707 ( .A(n_1659), .B(n_1505), .Y(n_1707) );
INVxp67_ASAP7_75t_L g1708 ( .A(n_1621), .Y(n_1708) );
NOR2x1p5_ASAP7_75t_L g1709 ( .A(n_1682), .B(n_1506), .Y(n_1709) );
OR2x2_ASAP7_75t_L g1710 ( .A(n_1674), .B(n_1601), .Y(n_1710) );
INVx2_ASAP7_75t_SL g1711 ( .A(n_1628), .Y(n_1711) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1613), .Y(n_1712) );
OR2x2_ASAP7_75t_L g1713 ( .A(n_1685), .B(n_1604), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1683), .B(n_1527), .Y(n_1714) );
O2A1O1Ixp33_ASAP7_75t_L g1715 ( .A1(n_1635), .A2(n_1581), .B(n_1523), .C(n_1546), .Y(n_1715) );
OAI22xp5_ASAP7_75t_L g1716 ( .A1(n_1681), .A2(n_1597), .B1(n_1595), .B2(n_1593), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_1644), .B(n_1537), .Y(n_1717) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1613), .Y(n_1718) );
OR2x2_ASAP7_75t_L g1719 ( .A(n_1640), .B(n_1509), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1679), .B(n_1591), .Y(n_1720) );
NOR2xp33_ASAP7_75t_SL g1721 ( .A(n_1682), .B(n_1589), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1679), .B(n_1591), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1668), .B(n_1615), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1634), .B(n_1535), .Y(n_1724) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1644), .B(n_1512), .Y(n_1725) );
NAND2x1_ASAP7_75t_L g1726 ( .A(n_1631), .B(n_1547), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1668), .B(n_1515), .Y(n_1727) );
AND2x4_ASAP7_75t_L g1728 ( .A(n_1645), .B(n_1547), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1634), .B(n_1585), .Y(n_1729) );
AND2x4_ASAP7_75t_L g1730 ( .A(n_1645), .B(n_1544), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1648), .B(n_1532), .Y(n_1731) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1617), .Y(n_1732) );
INVx3_ASAP7_75t_L g1733 ( .A(n_1676), .Y(n_1733) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1617), .Y(n_1734) );
OR2x2_ASAP7_75t_L g1735 ( .A(n_1648), .B(n_1636), .Y(n_1735) );
INVxp67_ASAP7_75t_L g1736 ( .A(n_1667), .Y(n_1736) );
NOR2xp33_ASAP7_75t_L g1737 ( .A(n_1651), .B(n_1607), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1738 ( .A(n_1654), .B(n_1526), .Y(n_1738) );
OR2x2_ASAP7_75t_L g1739 ( .A(n_1620), .B(n_1578), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1615), .B(n_1580), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1637), .B(n_1585), .Y(n_1741) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1625), .Y(n_1742) );
AND2x4_ASAP7_75t_L g1743 ( .A(n_1645), .B(n_1586), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1637), .B(n_1586), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1638), .B(n_1562), .Y(n_1745) );
AND2x4_ASAP7_75t_L g1746 ( .A(n_1645), .B(n_1525), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1638), .B(n_1562), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1622), .B(n_1556), .Y(n_1748) );
INVx2_ASAP7_75t_SL g1749 ( .A(n_1667), .Y(n_1749) );
OR2x2_ASAP7_75t_L g1750 ( .A(n_1687), .B(n_1669), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1690), .B(n_1661), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1752 ( .A(n_1693), .B(n_1654), .Y(n_1752) );
AND2x2_ASAP7_75t_SL g1753 ( .A(n_1728), .B(n_1653), .Y(n_1753) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1701), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_1729), .B(n_1647), .Y(n_1755) );
NAND2xp5_ASAP7_75t_L g1756 ( .A(n_1692), .B(n_1647), .Y(n_1756) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1703), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1702), .B(n_1671), .Y(n_1758) );
HB1xp67_ASAP7_75t_L g1759 ( .A(n_1708), .Y(n_1759) );
INVxp67_ASAP7_75t_SL g1760 ( .A(n_1736), .Y(n_1760) );
INVx1_ASAP7_75t_SL g1761 ( .A(n_1711), .Y(n_1761) );
NAND2xp5_ASAP7_75t_L g1762 ( .A(n_1688), .B(n_1671), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1729), .B(n_1673), .Y(n_1763) );
INVxp67_ASAP7_75t_SL g1764 ( .A(n_1736), .Y(n_1764) );
INVxp67_ASAP7_75t_L g1765 ( .A(n_1749), .Y(n_1765) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1688), .B(n_1663), .Y(n_1766) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1705), .Y(n_1767) );
NOR2xp33_ASAP7_75t_SL g1768 ( .A(n_1721), .B(n_1686), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1738), .B(n_1663), .Y(n_1769) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1724), .B(n_1661), .Y(n_1770) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_1724), .B(n_1665), .Y(n_1771) );
NAND2xp5_ASAP7_75t_L g1772 ( .A(n_1741), .B(n_1665), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1773 ( .A(n_1741), .B(n_1629), .Y(n_1773) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1699), .B(n_1629), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1744), .B(n_1673), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1744), .B(n_1657), .Y(n_1776) );
INVx1_ASAP7_75t_SL g1777 ( .A(n_1711), .Y(n_1777) );
INVx1_ASAP7_75t_SL g1778 ( .A(n_1696), .Y(n_1778) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1712), .Y(n_1779) );
INVx1_ASAP7_75t_SL g1780 ( .A(n_1710), .Y(n_1780) );
OR2x2_ASAP7_75t_L g1781 ( .A(n_1704), .B(n_1620), .Y(n_1781) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1718), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1745), .B(n_1657), .Y(n_1783) );
INVx2_ASAP7_75t_L g1784 ( .A(n_1697), .Y(n_1784) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1732), .Y(n_1785) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1734), .Y(n_1786) );
NAND2xp5_ASAP7_75t_L g1787 ( .A(n_1708), .B(n_1630), .Y(n_1787) );
OAI22xp33_ASAP7_75t_L g1788 ( .A1(n_1691), .A2(n_1595), .B1(n_1593), .B2(n_1651), .Y(n_1788) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1742), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1790 ( .A(n_1735), .B(n_1630), .Y(n_1790) );
INVx2_ASAP7_75t_L g1791 ( .A(n_1697), .Y(n_1791) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1745), .B(n_1660), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1747), .B(n_1660), .Y(n_1793) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1754), .B(n_1747), .Y(n_1794) );
OR2x2_ASAP7_75t_L g1795 ( .A(n_1770), .B(n_1739), .Y(n_1795) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1759), .Y(n_1796) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1750), .Y(n_1797) );
OAI22xp5_ASAP7_75t_L g1798 ( .A1(n_1753), .A2(n_1700), .B1(n_1709), .B2(n_1691), .Y(n_1798) );
AOI22xp33_ASAP7_75t_SL g1799 ( .A1(n_1753), .A2(n_1695), .B1(n_1730), .B2(n_1716), .Y(n_1799) );
NAND2xp5_ASAP7_75t_L g1800 ( .A(n_1754), .B(n_1717), .Y(n_1800) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1750), .Y(n_1801) );
AOI221xp5_ASAP7_75t_L g1802 ( .A1(n_1752), .A2(n_1715), .B1(n_1706), .B2(n_1737), .C(n_1731), .Y(n_1802) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1751), .Y(n_1803) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1757), .B(n_1707), .Y(n_1804) );
OAI21xp33_ASAP7_75t_L g1805 ( .A1(n_1768), .A2(n_1730), .B(n_1706), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1763), .B(n_1723), .Y(n_1806) );
INVx2_ASAP7_75t_SL g1807 ( .A(n_1761), .Y(n_1807) );
NAND2x1_ASAP7_75t_L g1808 ( .A(n_1770), .B(n_1733), .Y(n_1808) );
INVx1_ASAP7_75t_SL g1809 ( .A(n_1777), .Y(n_1809) );
NAND2xp5_ASAP7_75t_L g1810 ( .A(n_1757), .B(n_1662), .Y(n_1810) );
AOI21xp5_ASAP7_75t_L g1811 ( .A1(n_1753), .A2(n_1726), .B(n_1691), .Y(n_1811) );
AND2x2_ASAP7_75t_L g1812 ( .A(n_1763), .B(n_1714), .Y(n_1812) );
AOI21xp5_ASAP7_75t_L g1813 ( .A1(n_1768), .A2(n_1700), .B(n_1749), .Y(n_1813) );
AOI22xp5_ASAP7_75t_L g1814 ( .A1(n_1788), .A2(n_1737), .B1(n_1664), .B2(n_1727), .Y(n_1814) );
INVx2_ASAP7_75t_SL g1815 ( .A(n_1751), .Y(n_1815) );
AOI22xp33_ASAP7_75t_L g1816 ( .A1(n_1778), .A2(n_1730), .B1(n_1646), .B2(n_1678), .Y(n_1816) );
AOI21xp33_ASAP7_75t_SL g1817 ( .A1(n_1765), .A2(n_1614), .B(n_1733), .Y(n_1817) );
AOI22xp5_ASAP7_75t_L g1818 ( .A1(n_1780), .A2(n_1675), .B1(n_1689), .B2(n_1698), .Y(n_1818) );
INVx2_ASAP7_75t_L g1819 ( .A(n_1784), .Y(n_1819) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1767), .Y(n_1820) );
AOI22xp5_ASAP7_75t_L g1821 ( .A1(n_1760), .A2(n_1698), .B1(n_1689), .B2(n_1740), .Y(n_1821) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1767), .Y(n_1822) );
INVx3_ASAP7_75t_L g1823 ( .A(n_1784), .Y(n_1823) );
AOI21xp33_ASAP7_75t_L g1824 ( .A1(n_1798), .A2(n_1550), .B(n_1666), .Y(n_1824) );
INVxp67_ASAP7_75t_L g1825 ( .A(n_1807), .Y(n_1825) );
NAND2xp5_ASAP7_75t_L g1826 ( .A(n_1797), .B(n_1755), .Y(n_1826) );
AOI222xp33_ASAP7_75t_L g1827 ( .A1(n_1798), .A2(n_1764), .B1(n_1756), .B2(n_1787), .C1(n_1755), .C2(n_1775), .Y(n_1827) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1794), .Y(n_1828) );
OAI22xp5_ASAP7_75t_L g1829 ( .A1(n_1799), .A2(n_1773), .B1(n_1781), .B2(n_1771), .Y(n_1829) );
AOI322xp5_ASAP7_75t_L g1830 ( .A1(n_1802), .A2(n_1762), .A3(n_1775), .B1(n_1776), .B2(n_1758), .C1(n_1793), .C2(n_1783), .Y(n_1830) );
OAI222xp33_ASAP7_75t_L g1831 ( .A1(n_1813), .A2(n_1713), .B1(n_1781), .B2(n_1772), .C1(n_1652), .C2(n_1719), .Y(n_1831) );
AOI211xp5_ASAP7_75t_L g1832 ( .A1(n_1805), .A2(n_1677), .B(n_1733), .C(n_1672), .Y(n_1832) );
OAI21xp5_ASAP7_75t_L g1833 ( .A1(n_1809), .A2(n_1614), .B(n_1792), .Y(n_1833) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1794), .Y(n_1834) );
AOI21xp5_ASAP7_75t_L g1835 ( .A1(n_1811), .A2(n_1676), .B(n_1790), .Y(n_1835) );
OAI22xp33_ASAP7_75t_L g1836 ( .A1(n_1808), .A2(n_1766), .B1(n_1774), .B2(n_1769), .Y(n_1836) );
AOI22xp5_ASAP7_75t_L g1837 ( .A1(n_1818), .A2(n_1694), .B1(n_1689), .B2(n_1698), .Y(n_1837) );
OAI322xp33_ASAP7_75t_SL g1838 ( .A1(n_1803), .A2(n_1569), .A3(n_1528), .B1(n_1510), .B2(n_1511), .C1(n_1789), .C2(n_1782), .Y(n_1838) );
AOI22xp33_ASAP7_75t_L g1839 ( .A1(n_1801), .A2(n_1646), .B1(n_1746), .B2(n_1672), .Y(n_1839) );
AOI221xp5_ASAP7_75t_L g1840 ( .A1(n_1796), .A2(n_1779), .B1(n_1782), .B2(n_1789), .C(n_1786), .Y(n_1840) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1804), .Y(n_1841) );
A2O1A1Ixp33_ASAP7_75t_L g1842 ( .A1(n_1817), .A2(n_1602), .B(n_1776), .C(n_1792), .Y(n_1842) );
AOI21xp33_ASAP7_75t_SL g1843 ( .A1(n_1815), .A2(n_1614), .B(n_1652), .Y(n_1843) );
AOI22xp33_ASAP7_75t_SL g1844 ( .A1(n_1823), .A2(n_1728), .B1(n_1746), .B2(n_1793), .Y(n_1844) );
NOR2xp33_ASAP7_75t_R g1845 ( .A(n_1825), .B(n_1795), .Y(n_1845) );
AOI221xp5_ASAP7_75t_L g1846 ( .A1(n_1838), .A2(n_1800), .B1(n_1804), .B2(n_1816), .C(n_1810), .Y(n_1846) );
NAND3xp33_ASAP7_75t_L g1847 ( .A(n_1827), .B(n_1814), .C(n_1821), .Y(n_1847) );
NAND3xp33_ASAP7_75t_L g1848 ( .A(n_1829), .B(n_1822), .C(n_1820), .Y(n_1848) );
OR2x2_ASAP7_75t_L g1849 ( .A(n_1828), .B(n_1810), .Y(n_1849) );
AOI21xp5_ASAP7_75t_L g1850 ( .A1(n_1831), .A2(n_1800), .B(n_1823), .Y(n_1850) );
AOI31xp33_ASAP7_75t_L g1851 ( .A1(n_1832), .A2(n_1582), .A3(n_1806), .B(n_1812), .Y(n_1851) );
AOI322xp5_ASAP7_75t_L g1852 ( .A1(n_1836), .A2(n_1783), .A3(n_1720), .B1(n_1722), .B2(n_1748), .C1(n_1662), .C2(n_1819), .Y(n_1852) );
NAND2xp5_ASAP7_75t_L g1853 ( .A(n_1830), .B(n_1779), .Y(n_1853) );
OAI211xp5_ASAP7_75t_SL g1854 ( .A1(n_1837), .A2(n_1582), .B(n_1655), .C(n_1642), .Y(n_1854) );
O2A1O1Ixp33_ASAP7_75t_L g1855 ( .A1(n_1831), .A2(n_1551), .B(n_1555), .C(n_1611), .Y(n_1855) );
OAI221xp5_ASAP7_75t_L g1856 ( .A1(n_1844), .A2(n_1785), .B1(n_1786), .B2(n_1725), .C(n_1631), .Y(n_1856) );
AOI221xp5_ASAP7_75t_L g1857 ( .A1(n_1841), .A2(n_1785), .B1(n_1677), .B2(n_1791), .C(n_1584), .Y(n_1857) );
NOR4xp75_ASAP7_75t_L g1858 ( .A(n_1833), .B(n_1587), .C(n_1516), .D(n_1536), .Y(n_1858) );
AOI21xp5_ASAP7_75t_L g1859 ( .A1(n_1842), .A2(n_1791), .B(n_1541), .Y(n_1859) );
AOI221xp5_ASAP7_75t_L g1860 ( .A1(n_1824), .A2(n_1748), .B1(n_1746), .B2(n_1622), .C(n_1624), .Y(n_1860) );
NAND2xp5_ASAP7_75t_L g1861 ( .A(n_1846), .B(n_1834), .Y(n_1861) );
OAI211xp5_ASAP7_75t_L g1862 ( .A1(n_1845), .A2(n_1847), .B(n_1853), .C(n_1852), .Y(n_1862) );
A2O1A1Ixp33_ASAP7_75t_L g1863 ( .A1(n_1855), .A2(n_1835), .B(n_1843), .C(n_1840), .Y(n_1863) );
NAND2xp5_ASAP7_75t_L g1864 ( .A(n_1860), .B(n_1826), .Y(n_1864) );
NAND3xp33_ASAP7_75t_L g1865 ( .A(n_1848), .B(n_1839), .C(n_1605), .Y(n_1865) );
NOR3xp33_ASAP7_75t_L g1866 ( .A(n_1856), .B(n_1525), .C(n_1616), .Y(n_1866) );
NAND2xp5_ASAP7_75t_SL g1867 ( .A(n_1851), .B(n_1728), .Y(n_1867) );
AOI21xp5_ASAP7_75t_L g1868 ( .A1(n_1850), .A2(n_1642), .B(n_1587), .Y(n_1868) );
NOR2xp33_ASAP7_75t_L g1869 ( .A(n_1849), .B(n_1743), .Y(n_1869) );
NAND4xp25_ASAP7_75t_L g1870 ( .A(n_1854), .B(n_1598), .C(n_1594), .D(n_1588), .Y(n_1870) );
NAND2xp5_ASAP7_75t_SL g1871 ( .A(n_1857), .B(n_1743), .Y(n_1871) );
OR2x2_ASAP7_75t_L g1872 ( .A(n_1861), .B(n_1859), .Y(n_1872) );
NAND4xp25_ASAP7_75t_L g1873 ( .A(n_1862), .B(n_1858), .C(n_1594), .D(n_1598), .Y(n_1873) );
NAND3xp33_ASAP7_75t_L g1874 ( .A(n_1863), .B(n_1868), .C(n_1866), .Y(n_1874) );
NAND2xp5_ASAP7_75t_L g1875 ( .A(n_1864), .B(n_1624), .Y(n_1875) );
NAND4xp75_ASAP7_75t_L g1876 ( .A(n_1867), .B(n_1588), .C(n_1606), .D(n_1609), .Y(n_1876) );
OAI211xp5_ASAP7_75t_SL g1877 ( .A1(n_1871), .A2(n_1525), .B(n_1656), .C(n_1516), .Y(n_1877) );
NAND3xp33_ASAP7_75t_SL g1878 ( .A(n_1865), .B(n_1656), .C(n_1608), .Y(n_1878) );
HB1xp67_ASAP7_75t_L g1879 ( .A(n_1869), .Y(n_1879) );
AND3x1_ASAP7_75t_L g1880 ( .A(n_1879), .B(n_1870), .C(n_1606), .Y(n_1880) );
NOR4xp25_ASAP7_75t_L g1881 ( .A(n_1874), .B(n_1609), .C(n_1625), .D(n_1627), .Y(n_1881) );
NOR2xp67_ASAP7_75t_L g1882 ( .A(n_1873), .B(n_1616), .Y(n_1882) );
AND2x4_ASAP7_75t_L g1883 ( .A(n_1875), .B(n_1743), .Y(n_1883) );
NOR3xp33_ASAP7_75t_L g1884 ( .A(n_1872), .B(n_1633), .C(n_1616), .Y(n_1884) );
INVx3_ASAP7_75t_SL g1885 ( .A(n_1877), .Y(n_1885) );
AND2x4_ASAP7_75t_L g1886 ( .A(n_1884), .B(n_1876), .Y(n_1886) );
INVx2_ASAP7_75t_L g1887 ( .A(n_1883), .Y(n_1887) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1882), .Y(n_1888) );
XNOR2xp5_ASAP7_75t_L g1889 ( .A(n_1880), .B(n_1878), .Y(n_1889) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1885), .Y(n_1890) );
NOR3xp33_ASAP7_75t_L g1891 ( .A(n_1890), .B(n_1881), .C(n_1603), .Y(n_1891) );
BUFx2_ASAP7_75t_L g1892 ( .A(n_1887), .Y(n_1892) );
BUFx2_ASAP7_75t_L g1893 ( .A(n_1887), .Y(n_1893) );
INVx1_ASAP7_75t_SL g1894 ( .A(n_1888), .Y(n_1894) );
AOI222xp33_ASAP7_75t_L g1895 ( .A1(n_1892), .A2(n_1889), .B1(n_1886), .B2(n_1612), .C1(n_1608), .C2(n_1670), .Y(n_1895) );
OAI21xp33_ASAP7_75t_L g1896 ( .A1(n_1894), .A2(n_1886), .B(n_1612), .Y(n_1896) );
XNOR2xp5_ASAP7_75t_L g1897 ( .A(n_1893), .B(n_1886), .Y(n_1897) );
AOI21xp5_ASAP7_75t_L g1898 ( .A1(n_1891), .A2(n_1612), .B(n_1631), .Y(n_1898) );
AOI21xp5_ASAP7_75t_L g1899 ( .A1(n_1897), .A2(n_1631), .B(n_1536), .Y(n_1899) );
OAI21xp5_ASAP7_75t_L g1900 ( .A1(n_1896), .A2(n_1670), .B(n_1646), .Y(n_1900) );
OAI21xp5_ASAP7_75t_L g1901 ( .A1(n_1895), .A2(n_1670), .B(n_1646), .Y(n_1901) );
OAI22xp33_ASAP7_75t_L g1902 ( .A1(n_1898), .A2(n_1641), .B1(n_1561), .B2(n_1633), .Y(n_1902) );
UNKNOWN g1903 ( );
OR2x6_ASAP7_75t_L g1904 ( .A(n_1900), .B(n_1561), .Y(n_1904) );
NAND2xp5_ASAP7_75t_L g1905 ( .A(n_1902), .B(n_1633), .Y(n_1905) );
AOI221x1_ASAP7_75t_L g1906 ( .A1(n_1901), .A2(n_1561), .B1(n_1670), .B2(n_1643), .C(n_1639), .Y(n_1906) );
AOI22xp5_ASAP7_75t_L g1907 ( .A1(n_1903), .A2(n_1904), .B1(n_1905), .B2(n_1906), .Y(n_1907) );
endmodule