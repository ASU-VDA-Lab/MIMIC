module fake_netlist_6_389_n_1662 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1662);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1662;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_10),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_13),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_57),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_21),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_104),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_14),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_16),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_26),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_35),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_56),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_24),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_76),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_30),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_113),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_86),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_75),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_7),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_54),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_48),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

INVxp67_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_66),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_42),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_77),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_85),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_25),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_44),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_38),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_51),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_28),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_44),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_41),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_14),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_55),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_20),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_95),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_81),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_67),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_19),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_62),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_90),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_23),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_52),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_49),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_3),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_72),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_12),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_120),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_98),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_80),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_12),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_43),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_25),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_84),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_137),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_39),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_105),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_88),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_112),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_59),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_15),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_60),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_36),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_26),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_31),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_15),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_111),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_106),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_89),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_16),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_110),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_129),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_33),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_107),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_31),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_74),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_79),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_143),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_46),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_101),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_41),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_40),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_133),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_38),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_149),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_42),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_3),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_97),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_40),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_123),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_39),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_94),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_32),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_18),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_11),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_48),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_0),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_162),
.B(n_1),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_151),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_168),
.B(n_1),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_214),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_168),
.B(n_2),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_151),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_150),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_234),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_186),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_154),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_150),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_172),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_186),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_152),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_172),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_155),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_153),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_160),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_4),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_161),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_188),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_188),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_157),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_193),
.B(n_4),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_194),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_158),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_164),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_171),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_191),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_203),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_206),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_196),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_207),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_196),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_R g337 ( 
.A(n_266),
.B(n_5),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_209),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_270),
.B(n_5),
.Y(n_339)
);

BUFx6f_ASAP7_75t_SL g340 ( 
.A(n_167),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_198),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_159),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_218),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_270),
.B(n_6),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_163),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_166),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_169),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_279),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_201),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_170),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_198),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_173),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_174),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_175),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_202),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_176),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_255),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_177),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_223),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_227),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_202),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_204),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_204),
.B(n_212),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_165),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_192),
.B(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_212),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_231),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_213),
.B(n_9),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_255),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_213),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_242),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_245),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_165),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_267),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_302),
.A2(n_256),
.B1(n_238),
.B2(n_295),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_267),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_365),
.A2(n_304),
.B(n_300),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_321),
.B(n_285),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_165),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_305),
.B(n_285),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_298),
.B(n_167),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_268),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_268),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_192),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_268),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_268),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_336),
.B(n_268),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_309),
.B(n_310),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_341),
.A2(n_208),
.B(n_199),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_178),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_199),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_309),
.B(n_215),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_362),
.B(n_208),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_366),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_310),
.B(n_335),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_299),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_299),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_301),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_193),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_303),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_325),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_314),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_314),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_317),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_318),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_318),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_320),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_320),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_328),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_329),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_306),
.A2(n_179),
.B1(n_228),
.B2(n_197),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_329),
.B(n_287),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_307),
.B(n_287),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_330),
.B(n_184),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_438),
.B(n_348),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_438),
.B(n_330),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_438),
.B(n_331),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_417),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_215),
.Y(n_453)
);

INVx4_ASAP7_75t_SL g454 ( 
.A(n_399),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_372),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_378),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_308),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_316),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_438),
.B(n_331),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_438),
.B(n_332),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_324),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_374),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_438),
.B(n_332),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_201),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_398),
.B(n_334),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_376),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_376),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_423),
.B(n_334),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_399),
.B(n_338),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_376),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_392),
.B(n_426),
.Y(n_489)
);

CKINVDCx11_ASAP7_75t_R g490 ( 
.A(n_390),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_408),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_380),
.B(n_327),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_379),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_421),
.A2(n_337),
.B1(n_399),
.B2(n_394),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_429),
.B(n_156),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_390),
.B(n_338),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_438),
.B(n_343),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_400),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_342),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_405),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_398),
.B(n_388),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_417),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_377),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_377),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_398),
.B(n_343),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_438),
.B(n_359),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_423),
.B(n_359),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_426),
.B(n_428),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_382),
.B(n_217),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_377),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_398),
.B(n_360),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_417),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_403),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_404),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_377),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_411),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_379),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_393),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_383),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_428),
.B(n_360),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_383),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_398),
.B(n_367),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_382),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_398),
.B(n_388),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_394),
.B(n_226),
.C(n_217),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_390),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_428),
.B(n_345),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_382),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_393),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_428),
.B(n_346),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_415),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_423),
.A2(n_356),
.B1(n_350),
.B2(n_352),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_423),
.B(n_367),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_382),
.B(n_371),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_383),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_382),
.B(n_371),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_383),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_386),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_393),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_404),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_421),
.A2(n_437),
.B1(n_436),
.B2(n_432),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_441),
.B(n_181),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_416),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_419),
.B(n_225),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_386),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_393),
.Y(n_564)
);

BUFx6f_ASAP7_75t_SL g565 ( 
.A(n_429),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_386),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_431),
.B(n_347),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_399),
.A2(n_182),
.B1(n_225),
.B2(n_205),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_381),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_377),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_386),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_389),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_381),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_431),
.B(n_353),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_379),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_389),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_381),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_431),
.B(n_358),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_381),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_379),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_431),
.B(n_180),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_432),
.A2(n_219),
.B1(n_279),
.B2(n_253),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_429),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_441),
.B(n_254),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_399),
.A2(n_292),
.B1(n_296),
.B2(n_297),
.Y(n_585)
);

INVxp33_ASAP7_75t_SL g586 ( 
.A(n_401),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_441),
.A2(n_183),
.B1(n_290),
.B2(n_248),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_389),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_434),
.B(n_435),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_381),
.Y(n_590)
);

BUFx5_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_489),
.B(n_494),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_508),
.B(n_432),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_562),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_559),
.B(n_434),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_519),
.B(n_434),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_550),
.B(n_434),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_581),
.B(n_432),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_521),
.A2(n_404),
.B(n_405),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_569),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_554),
.B(n_435),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_476),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_452),
.B(n_432),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_494),
.B(n_435),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_522),
.B(n_435),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_560),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_468),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_452),
.B(n_432),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_532),
.B(n_483),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_499),
.B(n_429),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_499),
.B(n_429),
.Y(n_614)
);

AND2x6_ASAP7_75t_SL g615 ( 
.A(n_466),
.B(n_162),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_497),
.A2(n_437),
.B1(n_436),
.B2(n_419),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_497),
.A2(n_419),
.B1(n_418),
.B2(n_183),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_573),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_562),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_472),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_511),
.B(n_436),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_541),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_526),
.B(n_436),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_526),
.B(n_436),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_522),
.A2(n_539),
.B(n_510),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_522),
.B(n_437),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_449),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_472),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_579),
.Y(n_631)
);

BUFx6f_ASAP7_75t_SL g632 ( 
.A(n_476),
.Y(n_632)
);

INVxp33_ASAP7_75t_L g633 ( 
.A(n_560),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_585),
.A2(n_419),
.B1(n_418),
.B2(n_420),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_532),
.B(n_437),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_483),
.B(n_429),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_579),
.Y(n_637)
);

BUFx5_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_575),
.B(n_382),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_457),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_518),
.B(n_549),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_590),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_474),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_484),
.B(n_583),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_583),
.B(n_399),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_484),
.B(n_404),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_589),
.A2(n_406),
.B(n_397),
.C(n_440),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_575),
.B(n_382),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_549),
.B(n_404),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_538),
.B(n_404),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_580),
.B(n_399),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_541),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_457),
.B(n_441),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_474),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_506),
.B(n_425),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_580),
.B(n_399),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_491),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_538),
.B(n_404),
.Y(n_659)
);

NOR2x1p5_ASAP7_75t_L g660 ( 
.A(n_584),
.B(n_427),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_469),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_455),
.A2(n_399),
.B1(n_440),
.B2(n_425),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_477),
.B(n_399),
.Y(n_663)
);

INVx8_ASAP7_75t_L g664 ( 
.A(n_453),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_516),
.B(n_410),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_475),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_584),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_542),
.B(n_420),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_469),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_546),
.B(n_391),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_535),
.B(n_418),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_475),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_524),
.B(n_410),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_521),
.B(n_226),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_537),
.B(n_420),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_453),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_567),
.B(n_574),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_463),
.B(n_422),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_467),
.B(n_422),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_467),
.B(n_424),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_478),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_538),
.A2(n_397),
.B1(n_182),
.B2(n_235),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_471),
.B(n_424),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_471),
.B(n_424),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_543),
.B(n_406),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_543),
.A2(n_236),
.B1(n_190),
.B2(n_205),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_478),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_473),
.B(n_391),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_480),
.B(n_391),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_480),
.B(n_391),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_543),
.B(n_393),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_453),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_578),
.B(n_460),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_501),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_481),
.B(n_488),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_462),
.B(n_401),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_548),
.B(n_427),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_476),
.B(n_380),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_481),
.B(n_413),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_476),
.B(n_413),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_486),
.A2(n_387),
.B1(n_413),
.B2(n_430),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_450),
.B(n_451),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_482),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_482),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_485),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_485),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_488),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_464),
.A2(n_387),
.B1(n_433),
.B2(n_430),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_585),
.A2(n_259),
.B1(n_280),
.B2(n_246),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_448),
.B(n_439),
.C(n_380),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_493),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_521),
.B(n_409),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_498),
.B(n_387),
.Y(n_713)
);

AOI22x1_ASAP7_75t_L g714 ( 
.A1(n_498),
.A2(n_433),
.B1(n_387),
.B2(n_396),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_465),
.B(n_433),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_500),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_500),
.B(n_387),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_521),
.B(n_389),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_470),
.B(n_250),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_503),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_476),
.B(n_439),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_502),
.B(n_274),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_517),
.B(n_185),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_504),
.B(n_513),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_504),
.B(n_396),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_587),
.B(n_249),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_513),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_514),
.B(n_381),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_514),
.B(n_396),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_487),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_527),
.B(n_396),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_527),
.B(n_257),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_445),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_540),
.A2(n_239),
.B1(n_251),
.B2(n_262),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_531),
.B(n_412),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_531),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_528),
.B(n_412),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_487),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_544),
.B(n_412),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_544),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_528),
.B(n_412),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_540),
.A2(n_224),
.B1(n_190),
.B2(n_211),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_582),
.B(n_279),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_453),
.A2(n_412),
.B1(n_414),
.B2(n_229),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_547),
.B(n_412),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_547),
.B(n_258),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_552),
.B(n_260),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_528),
.B(n_414),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_553),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_553),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_495),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_561),
.B(n_414),
.Y(n_752)
);

O2A1O1Ixp5_ASAP7_75t_L g753 ( 
.A1(n_596),
.A2(n_561),
.B(n_446),
.C(n_444),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_597),
.B(n_453),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_597),
.B(n_453),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_728),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_728),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_626),
.Y(n_758)
);

AO22x1_ASAP7_75t_L g759 ( 
.A1(n_710),
.A2(n_586),
.B1(n_453),
.B2(n_271),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_593),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_642),
.A2(n_565),
.B1(n_586),
.B2(n_454),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_591),
.B(n_528),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_606),
.B(n_443),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_591),
.B(n_558),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_647),
.A2(n_558),
.B(n_456),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_642),
.A2(n_565),
.B1(n_454),
.B2(n_568),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_713),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_606),
.B(n_443),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_602),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_665),
.B(n_444),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_591),
.B(n_558),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_673),
.B(n_446),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_709),
.A2(n_617),
.B(n_616),
.C(n_677),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_618),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_622),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_719),
.A2(n_722),
.B(n_702),
.C(n_636),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_608),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_647),
.A2(n_558),
.B(n_456),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_733),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_737),
.A2(n_456),
.B(n_445),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_658),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_636),
.B(n_447),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_640),
.A2(n_409),
.B(n_447),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_630),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_737),
.A2(n_456),
.B(n_445),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_591),
.B(n_454),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_600),
.B(n_459),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_633),
.B(n_439),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_631),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_595),
.B(n_459),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_619),
.B(n_461),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_741),
.A2(n_456),
.B(n_445),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_591),
.B(n_454),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_696),
.B(n_490),
.C(n_281),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_670),
.B(n_461),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_607),
.A2(n_565),
.B1(n_251),
.B2(n_239),
.Y(n_798)
);

NOR2x1_ASAP7_75t_L g799 ( 
.A(n_635),
.B(n_693),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_613),
.A2(n_219),
.B1(n_492),
.B2(n_235),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_639),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_643),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_702),
.A2(n_507),
.B1(n_530),
.B2(n_495),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_741),
.A2(n_557),
.B(n_445),
.Y(n_804)
);

O2A1O1Ixp5_ASAP7_75t_L g805 ( 
.A1(n_596),
.A2(n_496),
.B(n_530),
.C(n_520),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_591),
.B(n_557),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_748),
.A2(n_557),
.B(n_545),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_609),
.B(n_492),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_748),
.A2(n_601),
.B(n_691),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_691),
.A2(n_557),
.B(n_545),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_675),
.B(n_496),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_649),
.A2(n_409),
.B(n_545),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_719),
.A2(n_505),
.B1(n_507),
.B2(n_525),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_607),
.A2(n_233),
.B1(n_262),
.B2(n_275),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_592),
.B(n_505),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_722),
.A2(n_509),
.B1(n_520),
.B2(n_525),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_651),
.A2(n_557),
.B(n_458),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_625),
.A2(n_409),
.B(n_479),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_612),
.B(n_509),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_608),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_667),
.B(n_219),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_628),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_614),
.A2(n_414),
.B1(n_252),
.B2(n_247),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_740),
.B(n_594),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_628),
.B(n_233),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_SL g826 ( 
.A1(n_598),
.A2(n_275),
.B(n_576),
.C(n_572),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_641),
.B(n_211),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_671),
.B(n_707),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_638),
.B(n_479),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_659),
.A2(n_533),
.B(n_479),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_653),
.B(n_167),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_641),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_650),
.A2(n_564),
.B(n_515),
.Y(n_833)
);

BUFx4f_ASAP7_75t_L g834 ( 
.A(n_661),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_696),
.B(n_219),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_638),
.B(n_512),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_671),
.A2(n_588),
.B(n_576),
.C(n_572),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_650),
.A2(n_512),
.B(n_515),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_711),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_646),
.A2(n_611),
.B(n_605),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_694),
.B(n_269),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_716),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_713),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_654),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_720),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_733),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_669),
.B(n_283),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_709),
.A2(n_407),
.B(n_414),
.C(n_222),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_660),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_733),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_727),
.B(n_523),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_736),
.B(n_523),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_654),
.B(n_414),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_621),
.A2(n_624),
.B(n_623),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_598),
.A2(n_555),
.B(n_571),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_656),
.B(n_286),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_698),
.B(n_407),
.Y(n_857)
);

AO21x1_ASAP7_75t_L g858 ( 
.A1(n_603),
.A2(n_588),
.B(n_566),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_617),
.A2(n_222),
.B(n_276),
.C(n_264),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_700),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_688),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_648),
.A2(n_555),
.B(n_566),
.C(n_563),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_638),
.B(n_529),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_685),
.A2(n_563),
.B(n_556),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_685),
.A2(n_556),
.B(n_551),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_749),
.B(n_534),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_634),
.A2(n_259),
.B(n_276),
.C(n_278),
.Y(n_867)
);

BUFx4f_ASAP7_75t_L g868 ( 
.A(n_721),
.Y(n_868)
);

AOI21x1_ASAP7_75t_L g869 ( 
.A1(n_718),
.A2(n_534),
.B(n_551),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_615),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_603),
.A2(n_536),
.B(n_570),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_750),
.B(n_536),
.Y(n_872)
);

NAND2x1_ASAP7_75t_L g873 ( 
.A(n_599),
.B(n_377),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_689),
.B(n_187),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_718),
.A2(n_570),
.B(n_377),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_690),
.B(n_189),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_715),
.A2(n_246),
.B(n_224),
.C(n_294),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_663),
.A2(n_570),
.B(n_377),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_682),
.B(n_195),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_682),
.B(n_200),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_712),
.A2(n_570),
.B(n_377),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_668),
.B(n_253),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_699),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_726),
.A2(n_236),
.B(n_294),
.C(n_243),
.Y(n_884)
);

AOI21x1_ASAP7_75t_L g885 ( 
.A1(n_674),
.A2(n_243),
.B(n_264),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_678),
.B(n_210),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_751),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_664),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_697),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_627),
.B(n_289),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_695),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_726),
.B(n_230),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_679),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_680),
.B(n_265),
.Y(n_894)
);

AO21x1_ASAP7_75t_L g895 ( 
.A1(n_634),
.A2(n_662),
.B(n_734),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_683),
.B(n_263),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_712),
.A2(n_570),
.B(n_293),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_638),
.B(n_261),
.Y(n_898)
);

AOI33xp33_ASAP7_75t_L g899 ( 
.A1(n_742),
.A2(n_278),
.A3(n_280),
.B1(n_288),
.B2(n_277),
.B3(n_22),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_652),
.A2(n_570),
.B(n_291),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_610),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_620),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_684),
.B(n_241),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_657),
.A2(n_717),
.B(n_638),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_732),
.B(n_240),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_676),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_732),
.B(n_244),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_746),
.B(n_237),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_735),
.A2(n_232),
.B(n_282),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_708),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_664),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_724),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_629),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_739),
.A2(n_273),
.B(n_272),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_729),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_745),
.A2(n_221),
.B(n_220),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_746),
.B(n_216),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_747),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_731),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_752),
.A2(n_288),
.B(n_58),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_701),
.A2(n_277),
.B(n_53),
.Y(n_922)
);

O2A1O1Ixp5_ASAP7_75t_L g923 ( 
.A1(n_747),
.A2(n_277),
.B(n_17),
.C(n_18),
.Y(n_923)
);

OAI321xp33_ASAP7_75t_L g924 ( 
.A1(n_742),
.A2(n_10),
.A3(n_17),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_686),
.B(n_28),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_809),
.A2(n_755),
.B(n_754),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_919),
.B(n_686),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_906),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_776),
.A2(n_723),
.B(n_645),
.C(n_730),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_912),
.B(n_645),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_820),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_892),
.A2(n_604),
.B1(n_632),
.B2(n_744),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_922),
.A2(n_676),
.B(n_692),
.C(n_664),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_888),
.B(n_692),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_808),
.B(n_738),
.C(n_644),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_906),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_820),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_822),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_868),
.B(n_687),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_760),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_835),
.B(n_655),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_844),
.B(n_666),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_891),
.A2(n_714),
.B1(n_706),
.B2(n_705),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_844),
.B(n_704),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_841),
.B(n_703),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_841),
.B(n_681),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_788),
.B(n_672),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_868),
.B(n_68),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_918),
.A2(n_78),
.B1(n_138),
.B2(n_135),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_769),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_779),
.Y(n_951)
);

AO22x1_ASAP7_75t_L g952 ( 
.A1(n_870),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_918),
.A2(n_34),
.B1(n_37),
.B2(n_43),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_822),
.Y(n_954)
);

CKINVDCx16_ASAP7_75t_R g955 ( 
.A(n_775),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_773),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_788),
.B(n_45),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_912),
.B(n_47),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_840),
.A2(n_92),
.B(n_132),
.Y(n_960)
);

AO32x2_ASAP7_75t_L g961 ( 
.A1(n_814),
.A2(n_49),
.A3(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_784),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_834),
.B(n_103),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_906),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_906),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_770),
.A2(n_99),
.B(n_64),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_832),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_781),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_SL g969 ( 
.A1(n_890),
.A2(n_109),
.B(n_65),
.C(n_82),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_849),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_834),
.B(n_83),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_827),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_777),
.B(n_114),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_860),
.A2(n_117),
.B1(n_124),
.B2(n_147),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_800),
.A2(n_895),
.B1(n_860),
.B2(n_925),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_883),
.B(n_861),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_889),
.A2(n_890),
.B(n_856),
.C(n_867),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_883),
.B(n_861),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_832),
.B(n_808),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_893),
.B(n_828),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_772),
.A2(n_854),
.B(n_782),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_910),
.A2(n_758),
.B1(n_766),
.B2(n_761),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_SL g983 ( 
.A(n_796),
.B(n_924),
.C(n_884),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_779),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_827),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_857),
.B(n_767),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_853),
.B(n_799),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_767),
.B(n_843),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_825),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_843),
.B(n_825),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_758),
.A2(n_768),
.B1(n_763),
.B2(n_824),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_821),
.B(n_847),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_798),
.A2(n_905),
.B(n_908),
.Y(n_993)
);

OAI22xp33_ASAP7_75t_L g994 ( 
.A1(n_907),
.A2(n_856),
.B1(n_791),
.B2(n_802),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_756),
.B(n_757),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_904),
.A2(n_762),
.B(n_771),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_839),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_842),
.B(n_882),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_779),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_762),
.A2(n_764),
.B(n_771),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_913),
.B(n_916),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_920),
.B(n_797),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_764),
.A2(n_818),
.B(n_787),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_757),
.B(n_790),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_831),
.Y(n_1005)
);

CKINVDCx6p67_ASAP7_75t_R g1006 ( 
.A(n_779),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_819),
.B(n_845),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_801),
.B(n_899),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_859),
.A2(n_753),
.B(n_848),
.C(n_879),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_789),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_877),
.A2(n_923),
.B(n_811),
.C(n_876),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_880),
.A2(n_888),
.B1(n_911),
.B2(n_874),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_923),
.A2(n_815),
.B(n_793),
.C(n_792),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_783),
.A2(n_806),
.B(n_812),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_759),
.B(n_886),
.Y(n_1015)
);

INVx6_ASAP7_75t_L g1016 ( 
.A(n_789),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_866),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_901),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_894),
.A2(n_896),
.B1(n_903),
.B2(n_902),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_753),
.A2(n_858),
.B(n_898),
.C(n_805),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_837),
.A2(n_872),
.B(n_826),
.C(n_862),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_914),
.B(n_887),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_789),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_806),
.A2(n_898),
.B(n_765),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_887),
.B(n_823),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_805),
.A2(n_921),
.B(n_838),
.C(n_833),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_911),
.A2(n_851),
.B1(n_852),
.B2(n_846),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_SL g1028 ( 
.A1(n_786),
.A2(n_795),
.B(n_871),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_789),
.Y(n_1029)
);

NAND2xp33_ASAP7_75t_L g1030 ( 
.A(n_846),
.B(n_850),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_778),
.A2(n_780),
.B(n_785),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_846),
.B(n_850),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_794),
.A2(n_804),
.B(n_807),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_SL g1034 ( 
.A(n_909),
.B(n_917),
.C(n_915),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_878),
.A2(n_817),
.B(n_881),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_850),
.A2(n_803),
.B1(n_813),
.B2(n_816),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_810),
.A2(n_829),
.B(n_863),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_850),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_864),
.A2(n_865),
.B(n_830),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_869),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_873),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_855),
.B(n_885),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_900),
.Y(n_1043)
);

BUFx12f_ASAP7_75t_L g1044 ( 
.A(n_897),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_875),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_836),
.A2(n_528),
.B(n_521),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_776),
.A2(n_607),
.B(n_627),
.Y(n_1047)
);

AND2x2_ASAP7_75t_SL g1048 ( 
.A(n_868),
.B(n_613),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_857),
.B(n_667),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_774),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_809),
.A2(n_528),
.B(n_521),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_760),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_809),
.A2(n_528),
.B(n_521),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_857),
.B(n_667),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_809),
.A2(n_528),
.B(n_521),
.Y(n_1055)
);

NAND2x1p5_ASAP7_75t_L g1056 ( 
.A(n_888),
.B(n_911),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_777),
.B(n_608),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_776),
.A2(n_606),
.B1(n_597),
.B2(n_892),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_892),
.A2(n_918),
.B1(n_693),
.B2(n_642),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_888),
.B(n_911),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_773),
.A2(n_363),
.B1(n_617),
.B2(n_924),
.C(n_709),
.Y(n_1061)
);

CKINVDCx11_ASAP7_75t_R g1062 ( 
.A(n_955),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1058),
.A2(n_1059),
.B(n_977),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1047),
.A2(n_1009),
.B(n_987),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1048),
.A2(n_1001),
.B1(n_998),
.B2(n_975),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_957),
.A2(n_1061),
.B(n_947),
.C(n_933),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_L g1067 ( 
.A(n_992),
.B(n_1061),
.C(n_953),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_931),
.Y(n_1068)
);

BUFx2_ASAP7_75t_SL g1069 ( 
.A(n_1057),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_981),
.A2(n_926),
.B(n_1051),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_969),
.A2(n_948),
.B(n_963),
.C(n_971),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_983),
.A2(n_1011),
.B(n_929),
.C(n_1015),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_981),
.A2(n_926),
.B(n_1055),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_980),
.A2(n_1054),
.B(n_1049),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_976),
.B(n_978),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_SL g1076 ( 
.A1(n_1012),
.A2(n_929),
.B(n_1011),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1051),
.A2(n_1055),
.B(n_1053),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1053),
.A2(n_1014),
.B(n_1003),
.Y(n_1078)
);

BUFx2_ASAP7_75t_SL g1079 ( 
.A(n_1057),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_945),
.A2(n_946),
.B(n_1002),
.C(n_1013),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_993),
.A2(n_1026),
.A3(n_1035),
.B(n_1014),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1003),
.A2(n_996),
.B(n_1035),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_935),
.B(n_956),
.C(n_927),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1017),
.B(n_941),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_956),
.A2(n_994),
.B(n_958),
.C(n_986),
.Y(n_1085)
);

AO32x2_ASAP7_75t_L g1086 ( 
.A1(n_982),
.A2(n_991),
.A3(n_1036),
.B1(n_943),
.B2(n_961),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_1024),
.A2(n_1037),
.B(n_1033),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_968),
.B(n_937),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1031),
.A2(n_1039),
.B(n_1037),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_997),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_938),
.B(n_967),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1024),
.A2(n_1000),
.B(n_1043),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1040),
.A2(n_1046),
.B(n_1000),
.Y(n_1093)
);

AO31x2_ASAP7_75t_L g1094 ( 
.A1(n_960),
.A2(n_1046),
.A3(n_1027),
.B(n_966),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1040),
.A2(n_1020),
.B(n_1021),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1008),
.B(n_942),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_954),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_1005),
.B(n_970),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1007),
.B(n_930),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1013),
.A2(n_1020),
.B(n_1028),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_1050),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1034),
.A2(n_1019),
.B(n_1030),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_940),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_990),
.B(n_989),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_950),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_962),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1021),
.A2(n_1041),
.B(n_1056),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1034),
.A2(n_1042),
.B(n_939),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_988),
.A2(n_1025),
.B(n_1022),
.Y(n_1109)
);

NOR2x1_ASAP7_75t_R g1110 ( 
.A(n_972),
.B(n_985),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_984),
.A2(n_934),
.B(n_1056),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_965),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1038),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_934),
.A2(n_1060),
.B(n_1041),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_932),
.A2(n_1004),
.B1(n_1052),
.B2(n_973),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_1018),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1032),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1016),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_928),
.A2(n_936),
.B(n_964),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_928),
.B(n_936),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_961),
.A2(n_1045),
.A3(n_1044),
.B(n_949),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_964),
.A2(n_973),
.B(n_1029),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_974),
.A2(n_952),
.B1(n_1006),
.B2(n_1016),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_995),
.A2(n_1016),
.B(n_999),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1023),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_951),
.B(n_999),
.Y(n_1126)
);

AO21x2_ASAP7_75t_L g1127 ( 
.A1(n_951),
.A2(n_926),
.B(n_1014),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_1023),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_959),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1058),
.A2(n_993),
.A3(n_776),
.B(n_1026),
.Y(n_1130)
);

AND4x1_ASAP7_75t_L g1131 ( 
.A(n_957),
.B(n_614),
.C(n_613),
.D(n_499),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_959),
.Y(n_1132)
);

AOI221x1_ASAP7_75t_L g1133 ( 
.A1(n_1058),
.A2(n_776),
.B1(n_977),
.B2(n_957),
.C(n_922),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1035),
.A2(n_1053),
.B(n_1051),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_955),
.B(n_302),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_957),
.A2(n_693),
.B(n_677),
.C(n_696),
.Y(n_1136)
);

NAND3x1_ASAP7_75t_L g1137 ( 
.A(n_957),
.B(n_710),
.C(n_808),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_959),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1059),
.B(n_919),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_955),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_959),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1001),
.B(n_612),
.Y(n_1142)
);

AOI222xp33_ASAP7_75t_L g1143 ( 
.A1(n_957),
.A2(n_439),
.B1(n_380),
.B2(n_1061),
.C1(n_743),
.C2(n_788),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1059),
.B(n_919),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_959),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_955),
.B(n_302),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_SL g1147 ( 
.A1(n_957),
.A2(n_1061),
.B1(n_726),
.B2(n_844),
.C(n_587),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1058),
.A2(n_776),
.B(n_1059),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1058),
.A2(n_776),
.B(n_1059),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1010),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_977),
.A2(n_776),
.B(n_1058),
.C(n_1061),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1035),
.A2(n_1053),
.B(n_1051),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1059),
.B(n_696),
.C(n_892),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_957),
.A2(n_693),
.B(n_677),
.C(n_696),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1001),
.B(n_612),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1057),
.B(n_990),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_981),
.A2(n_528),
.B(n_521),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_981),
.A2(n_528),
.B(n_521),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1058),
.A2(n_993),
.A3(n_776),
.B(n_1026),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_979),
.B(n_693),
.Y(n_1160)
);

CKINVDCx11_ASAP7_75t_R g1161 ( 
.A(n_955),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1058),
.A2(n_993),
.A3(n_776),
.B(n_1026),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1020),
.A2(n_1003),
.B(n_1014),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_957),
.A2(n_710),
.B1(n_892),
.B2(n_800),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1059),
.A2(n_1058),
.B1(n_776),
.B2(n_892),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1010),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1049),
.B(n_1054),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_981),
.A2(n_528),
.B(n_521),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_981),
.A2(n_528),
.B(n_521),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1058),
.A2(n_993),
.A3(n_776),
.B(n_1026),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_SL g1171 ( 
.A1(n_957),
.A2(n_492),
.B(n_800),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1059),
.A2(n_1058),
.B1(n_776),
.B2(n_892),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_981),
.A2(n_528),
.B(n_521),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1059),
.A2(n_892),
.B(n_1058),
.C(n_922),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_937),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_977),
.A2(n_776),
.B(n_1058),
.C(n_1061),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1059),
.A2(n_892),
.B(n_1058),
.C(n_922),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_981),
.A2(n_528),
.B(n_521),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_937),
.Y(n_1179)
);

INVx3_ASAP7_75t_SL g1180 ( 
.A(n_955),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_970),
.Y(n_1181)
);

AOI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1059),
.A2(n_892),
.B(n_696),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_937),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1035),
.A2(n_1053),
.B(n_1051),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1001),
.B(n_612),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_957),
.A2(n_693),
.B(n_677),
.C(n_696),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1001),
.B(n_612),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1001),
.B(n_612),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1057),
.B(n_990),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_SL g1190 ( 
.A(n_1044),
.B(n_888),
.Y(n_1190)
);

NOR2x1_ASAP7_75t_SL g1191 ( 
.A(n_1044),
.B(n_888),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_959),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_937),
.Y(n_1193)
);

OAI22x1_ASAP7_75t_L g1194 ( 
.A1(n_957),
.A2(n_1059),
.B1(n_492),
.B2(n_696),
.Y(n_1194)
);

AOI211x1_ASAP7_75t_L g1195 ( 
.A1(n_1001),
.A2(n_709),
.B(n_895),
.C(n_617),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1164),
.A2(n_1153),
.B1(n_1177),
.B2(n_1174),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1131),
.B(n_1115),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1175),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1143),
.A2(n_1182),
.B1(n_1194),
.B2(n_1067),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1165),
.A2(n_1172),
.B1(n_1149),
.B2(n_1148),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1088),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1063),
.A2(n_1065),
.B1(n_1160),
.B2(n_1171),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_SL g1203 ( 
.A(n_1150),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1133),
.A2(n_1155),
.B1(n_1142),
.B2(n_1187),
.Y(n_1204)
);

OAI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1131),
.A2(n_1115),
.B1(n_1083),
.B2(n_1144),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1083),
.A2(n_1139),
.B1(n_1074),
.B2(n_1096),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1074),
.A2(n_1064),
.B1(n_1185),
.B2(n_1188),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1179),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1135),
.A2(n_1146),
.B1(n_1137),
.B2(n_1100),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1099),
.A2(n_1084),
.B1(n_1101),
.B2(n_1075),
.Y(n_1210)
);

BUFx10_ASAP7_75t_L g1211 ( 
.A(n_1150),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1167),
.A2(n_1102),
.B1(n_1147),
.B2(n_1105),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1151),
.A2(n_1176),
.B1(n_1098),
.B2(n_1066),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1123),
.A2(n_1132),
.B1(n_1141),
.B2(n_1138),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1123),
.A2(n_1145),
.B1(n_1090),
.B2(n_1192),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1136),
.B(n_1154),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1103),
.A2(n_1106),
.B1(n_1183),
.B2(n_1193),
.Y(n_1217)
);

CKINVDCx11_ASAP7_75t_R g1218 ( 
.A(n_1181),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1166),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1091),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1120),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1062),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1068),
.A2(n_1097),
.B1(n_1186),
.B2(n_1180),
.Y(n_1223)
);

BUFx12f_ASAP7_75t_L g1224 ( 
.A(n_1161),
.Y(n_1224)
);

BUFx2_ASAP7_75t_SL g1225 ( 
.A(n_1140),
.Y(n_1225)
);

INVx11_ASAP7_75t_L g1226 ( 
.A(n_1069),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1109),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1080),
.A2(n_1072),
.B1(n_1079),
.B2(n_1116),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1166),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1163),
.A2(n_1113),
.B1(n_1078),
.B2(n_1108),
.Y(n_1230)
);

INVx8_ASAP7_75t_L g1231 ( 
.A(n_1166),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1117),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1163),
.A2(n_1082),
.B1(n_1189),
.B2(n_1156),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1104),
.Y(n_1234)
);

BUFx4_ASAP7_75t_SL g1235 ( 
.A(n_1125),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1189),
.B(n_1195),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1124),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1126),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1127),
.A2(n_1104),
.B1(n_1089),
.B2(n_1195),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1085),
.B(n_1122),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1118),
.Y(n_1241)
);

OAI22x1_ASAP7_75t_SL g1242 ( 
.A1(n_1110),
.A2(n_1112),
.B1(n_1191),
.B2(n_1190),
.Y(n_1242)
);

INVx6_ASAP7_75t_L g1243 ( 
.A(n_1110),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1128),
.B(n_1121),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1127),
.A2(n_1070),
.B1(n_1073),
.B2(n_1095),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1077),
.A2(n_1107),
.B1(n_1086),
.B2(n_1184),
.Y(n_1246)
);

BUFx12f_ASAP7_75t_L g1247 ( 
.A(n_1119),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1076),
.A2(n_1111),
.B1(n_1114),
.B2(n_1092),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1086),
.A2(n_1134),
.B1(n_1152),
.B2(n_1093),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1086),
.A2(n_1121),
.B1(n_1087),
.B2(n_1159),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1071),
.Y(n_1251)
);

BUFx8_ASAP7_75t_SL g1252 ( 
.A(n_1130),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1130),
.A2(n_1159),
.B(n_1170),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1157),
.B(n_1168),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1130),
.A2(n_1170),
.B1(n_1162),
.B2(n_1158),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1162),
.A2(n_1170),
.B(n_1169),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1081),
.Y(n_1257)
);

BUFx8_ASAP7_75t_L g1258 ( 
.A(n_1162),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1081),
.B(n_1094),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1094),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1173),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1178),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1164),
.A2(n_1153),
.B1(n_1177),
.B2(n_1174),
.Y(n_1263)
);

INVx8_ASAP7_75t_L g1264 ( 
.A(n_1150),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1150),
.Y(n_1265)
);

INVx6_ASAP7_75t_L g1266 ( 
.A(n_1150),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1150),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1160),
.B(n_1142),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1129),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1129),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1129),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1160),
.B(n_1142),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1171),
.A2(n_1153),
.B1(n_613),
.B2(n_614),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1150),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1150),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1088),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1150),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1160),
.B(n_1142),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1150),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1113),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1062),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1164),
.A2(n_1153),
.B1(n_1177),
.B2(n_1174),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1062),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1164),
.A2(n_1153),
.B1(n_1177),
.B2(n_1174),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1164),
.A2(n_1153),
.B1(n_1177),
.B2(n_1174),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1150),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1164),
.A2(n_1153),
.B1(n_1177),
.B2(n_1174),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1182),
.B2(n_1153),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1270),
.A2(n_1276),
.B1(n_1296),
.B2(n_1279),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1221),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1268),
.B(n_1275),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1257),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1204),
.B(n_1210),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1227),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1260),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1254),
.A2(n_1245),
.B(n_1261),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1237),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1233),
.B(n_1237),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1254),
.A2(n_1245),
.B(n_1261),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1244),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1259),
.B(n_1200),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1248),
.B(n_1197),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1241),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1204),
.B(n_1210),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1253),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1258),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1258),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1201),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1250),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1250),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1241),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1237),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1246),
.A2(n_1256),
.B(n_1249),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1262),
.A2(n_1249),
.B(n_1246),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1200),
.B(n_1197),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1207),
.B(n_1285),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1220),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1282),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1240),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1230),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1252),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1196),
.A2(n_1263),
.B1(n_1295),
.B2(n_1292),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1270),
.A2(n_1290),
.B1(n_1276),
.B2(n_1283),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1205),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1289),
.A2(n_1293),
.B(n_1216),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1230),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1239),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1233),
.A2(n_1207),
.B(n_1212),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1202),
.B(n_1212),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1198),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1238),
.B(n_1255),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1247),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1243),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1206),
.B(n_1272),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1255),
.B(n_1206),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1228),
.A2(n_1269),
.B(n_1273),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1277),
.A2(n_1215),
.B(n_1214),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1208),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1199),
.B(n_1271),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1214),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1272),
.A2(n_1280),
.B(n_1296),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1243),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1215),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1213),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1213),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1251),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1274),
.B(n_1279),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1274),
.B(n_1290),
.Y(n_1357)
);

INVx5_ASAP7_75t_SL g1358 ( 
.A(n_1226),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1217),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1199),
.B(n_1283),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1232),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1217),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1242),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1209),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1331),
.B(n_1280),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1299),
.B(n_1209),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1308),
.B(n_1223),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1334),
.B(n_1277),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1304),
.A2(n_1307),
.B(n_1334),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1327),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1297),
.B(n_1287),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1332),
.A2(n_1288),
.B1(n_1224),
.B2(n_1291),
.Y(n_1372)
);

OAI31xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1360),
.A2(n_1222),
.A3(n_1225),
.B(n_1203),
.Y(n_1373)
);

AOI221xp5_ASAP7_75t_L g1374 ( 
.A1(n_1356),
.A2(n_1357),
.B1(n_1360),
.B2(n_1297),
.C(n_1338),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1328),
.A2(n_1267),
.B(n_1264),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1338),
.A2(n_1264),
.B(n_1231),
.C(n_1278),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1350),
.A2(n_1234),
.B1(n_1203),
.B2(n_1266),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1322),
.A2(n_1235),
.B(n_1281),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1356),
.A2(n_1264),
.B(n_1231),
.C(n_1286),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1298),
.B(n_1278),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1357),
.A2(n_1343),
.B(n_1301),
.C(n_1312),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1341),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1325),
.B(n_1229),
.Y(n_1383)
);

OR2x6_ASAP7_75t_L g1384 ( 
.A(n_1310),
.B(n_1266),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1364),
.A2(n_1266),
.B(n_1281),
.C(n_1219),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1301),
.A2(n_1294),
.B1(n_1265),
.B2(n_1284),
.C(n_1211),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1328),
.B(n_1211),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1350),
.A2(n_1312),
.B(n_1324),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1324),
.B(n_1219),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1326),
.B(n_1284),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1325),
.B(n_1218),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1322),
.A2(n_1304),
.B(n_1307),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1305),
.B(n_1320),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1323),
.B(n_1333),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1350),
.B(n_1364),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1344),
.A2(n_1349),
.B1(n_1352),
.B2(n_1362),
.C(n_1354),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1350),
.A2(n_1341),
.B1(n_1346),
.B2(n_1363),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1314),
.A2(n_1315),
.B(n_1354),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1316),
.B(n_1359),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1361),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1363),
.A2(n_1315),
.B(n_1314),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1344),
.A2(n_1353),
.B(n_1352),
.C(n_1349),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1348),
.B(n_1341),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1355),
.A2(n_1330),
.B1(n_1353),
.B2(n_1363),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1341),
.B(n_1359),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1304),
.A2(n_1335),
.B(n_1329),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1346),
.A2(n_1355),
.B(n_1339),
.C(n_1310),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1302),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1317),
.A2(n_1318),
.B(n_1345),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1317),
.A2(n_1318),
.B(n_1345),
.Y(n_1410)
);

AOI21xp33_ASAP7_75t_L g1411 ( 
.A1(n_1365),
.A2(n_1346),
.B(n_1337),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1366),
.B(n_1347),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1406),
.B(n_1409),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1378),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1395),
.B(n_1302),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1400),
.Y(n_1416)
);

BUFx2_ASAP7_75t_SL g1417 ( 
.A(n_1398),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1410),
.B(n_1321),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1392),
.Y(n_1419)
);

INVx5_ASAP7_75t_L g1420 ( 
.A(n_1384),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1410),
.B(n_1306),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1410),
.B(n_1313),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1369),
.B(n_1306),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1408),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1395),
.B(n_1313),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1392),
.B(n_1306),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1392),
.B(n_1306),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1365),
.A2(n_1346),
.B1(n_1337),
.B2(n_1310),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1388),
.B(n_1335),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1399),
.B(n_1340),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1378),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1378),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1405),
.B(n_1309),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1414),
.Y(n_1434)
);

OAI211xp5_ASAP7_75t_L g1435 ( 
.A1(n_1411),
.A2(n_1374),
.B(n_1397),
.C(n_1407),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1416),
.Y(n_1436)
);

OAI21xp33_ASAP7_75t_L g1437 ( 
.A1(n_1429),
.A2(n_1368),
.B(n_1371),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1411),
.A2(n_1381),
.B1(n_1396),
.B2(n_1371),
.C(n_1402),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1416),
.B(n_1403),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1421),
.B(n_1394),
.Y(n_1440)
);

NAND4xp25_ASAP7_75t_L g1441 ( 
.A(n_1428),
.B(n_1373),
.C(n_1402),
.D(n_1389),
.Y(n_1441)
);

INVxp67_ASAP7_75t_SL g1442 ( 
.A(n_1422),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1422),
.B(n_1367),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1422),
.B(n_1415),
.Y(n_1444)
);

INVx3_ASAP7_75t_SL g1445 ( 
.A(n_1420),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1426),
.B(n_1393),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1420),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1417),
.B(n_1310),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1426),
.B(n_1383),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1419),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1413),
.A2(n_1303),
.B(n_1300),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1415),
.B(n_1336),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1426),
.B(n_1383),
.Y(n_1453)
);

O2A1O1Ixp5_ASAP7_75t_L g1454 ( 
.A1(n_1429),
.A2(n_1387),
.B(n_1375),
.C(n_1403),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1424),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1424),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1427),
.B(n_1393),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1455),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1455),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1434),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1447),
.B(n_1450),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1434),
.B(n_1414),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1434),
.B(n_1414),
.Y(n_1464)
);

AND2x4_ASAP7_75t_SL g1465 ( 
.A(n_1447),
.B(n_1384),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1440),
.B(n_1423),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1440),
.B(n_1423),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1452),
.B(n_1443),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1440),
.B(n_1423),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1451),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1444),
.B(n_1425),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1446),
.B(n_1431),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1443),
.B(n_1425),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1437),
.B(n_1391),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1446),
.B(n_1431),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1450),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1431),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1446),
.B(n_1431),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1447),
.B(n_1420),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1456),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_1431),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1452),
.B(n_1430),
.Y(n_1482)
);

NAND2x1_ASAP7_75t_L g1483 ( 
.A(n_1447),
.B(n_1432),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1456),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1444),
.B(n_1418),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1437),
.B(n_1430),
.Y(n_1486)
);

NOR2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1441),
.B(n_1447),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1461),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1479),
.B(n_1417),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1461),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1486),
.B(n_1436),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1466),
.B(n_1457),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1486),
.B(n_1436),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1458),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1474),
.B(n_1482),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1471),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1487),
.A2(n_1435),
.B1(n_1438),
.B2(n_1441),
.Y(n_1497)
);

NOR3xp33_ASAP7_75t_L g1498 ( 
.A(n_1462),
.B(n_1435),
.C(n_1438),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1462),
.B(n_1450),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1457),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1466),
.B(n_1457),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1458),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1463),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1479),
.B(n_1417),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1482),
.B(n_1391),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1459),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1463),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1459),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1463),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1467),
.B(n_1449),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1487),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1480),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1433),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1465),
.A2(n_1377),
.B1(n_1448),
.B2(n_1439),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1484),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1468),
.B(n_1433),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1464),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1464),
.Y(n_1519)
);

NAND2x1_ASAP7_75t_L g1520 ( 
.A(n_1476),
.B(n_1448),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1484),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1460),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1467),
.B(n_1469),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1460),
.Y(n_1525)
);

NAND2x2_ASAP7_75t_L g1526 ( 
.A(n_1483),
.B(n_1342),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1467),
.B(n_1453),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1471),
.B(n_1453),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1524),
.B(n_1469),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1533)
);

AOI211xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1497),
.A2(n_1372),
.B(n_1404),
.C(n_1386),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1502),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1495),
.B(n_1469),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1505),
.B(n_1453),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1498),
.B(n_1522),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1511),
.B(n_1370),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1462),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1528),
.B(n_1462),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1489),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1506),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1528),
.B(n_1462),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1464),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1505),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1492),
.B(n_1472),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1472),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1526),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1523),
.B(n_1485),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1508),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1500),
.B(n_1472),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1512),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1526),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1513),
.Y(n_1557)
);

OAI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1491),
.A2(n_1412),
.B(n_1428),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1493),
.B(n_1316),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1516),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1501),
.B(n_1475),
.Y(n_1561)
);

INVxp33_ASAP7_75t_L g1562 ( 
.A(n_1520),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1503),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1488),
.Y(n_1564)
);

AOI21xp33_ASAP7_75t_L g1565 ( 
.A1(n_1562),
.A2(n_1504),
.B(n_1489),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1540),
.B(n_1525),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1490),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1542),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1563),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1541),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1563),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1544),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1534),
.A2(n_1489),
.B(n_1504),
.C(n_1454),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1548),
.B(n_1564),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1563),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_SL g1576 ( 
.A1(n_1534),
.A2(n_1503),
.B(n_1483),
.C(n_1470),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1558),
.A2(n_1515),
.B1(n_1489),
.B2(n_1504),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1558),
.A2(n_1504),
.B(n_1454),
.Y(n_1578)
);

BUFx2_ASAP7_75t_SL g1579 ( 
.A(n_1564),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1537),
.B(n_1527),
.Y(n_1580)
);

INVxp33_ASAP7_75t_L g1581 ( 
.A(n_1559),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1544),
.A2(n_1412),
.B1(n_1330),
.B2(n_1448),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1531),
.B(n_1501),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1530),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1535),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1537),
.B(n_1379),
.C(n_1376),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1535),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1536),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1530),
.A2(n_1476),
.B(n_1385),
.C(n_1450),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1551),
.Y(n_1591)
);

OAI21xp33_ASAP7_75t_L g1592 ( 
.A1(n_1581),
.A2(n_1556),
.B(n_1543),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1572),
.B(n_1532),
.Y(n_1593)
);

AOI222xp33_ASAP7_75t_L g1594 ( 
.A1(n_1574),
.A2(n_1536),
.B1(n_1560),
.B2(n_1557),
.C1(n_1553),
.C2(n_1555),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1579),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1578),
.A2(n_1448),
.B1(n_1476),
.B2(n_1450),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1584),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1574),
.B(n_1556),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1567),
.A2(n_1560),
.B1(n_1557),
.B2(n_1555),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1577),
.A2(n_1539),
.B1(n_1479),
.B2(n_1547),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1566),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1582),
.A2(n_1479),
.B1(n_1547),
.B2(n_1532),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1576),
.A2(n_1545),
.B(n_1553),
.C(n_1470),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1569),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1571),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

NAND2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1586),
.B(n_1476),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1583),
.B(n_1542),
.Y(n_1608)
);

OAI211xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1592),
.A2(n_1576),
.B(n_1573),
.C(n_1565),
.Y(n_1609)
);

OAI31xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1596),
.A2(n_1588),
.A3(n_1587),
.B(n_1585),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1603),
.A2(n_1589),
.B(n_1582),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1601),
.A2(n_1597),
.B1(n_1607),
.B2(n_1595),
.C1(n_1599),
.C2(n_1590),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1593),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1604),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1595),
.B(n_1580),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1605),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1598),
.A2(n_1476),
.B1(n_1499),
.B2(n_1351),
.Y(n_1618)
);

OAI322xp33_ASAP7_75t_L g1619 ( 
.A1(n_1596),
.A2(n_1545),
.A3(n_1552),
.B1(n_1533),
.B2(n_1538),
.C1(n_1518),
.C2(n_1509),
.Y(n_1619)
);

OAI21xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1610),
.A2(n_1594),
.B(n_1599),
.Y(n_1620)
);

NAND4xp25_ASAP7_75t_L g1621 ( 
.A(n_1612),
.B(n_1590),
.C(n_1600),
.D(n_1606),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_SL g1622 ( 
.A(n_1611),
.B(n_1589),
.C(n_1602),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1615),
.Y(n_1623)
);

NAND4xp75_ASAP7_75t_L g1624 ( 
.A(n_1613),
.B(n_1608),
.C(n_1543),
.D(n_1546),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1617),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1610),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_SL g1627 ( 
.A(n_1609),
.B(n_1552),
.C(n_1538),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1618),
.A2(n_1499),
.B(n_1533),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1546),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1499),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1620),
.A2(n_1626),
.B1(n_1627),
.B2(n_1622),
.C(n_1621),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1625),
.B(n_1476),
.C(n_1619),
.Y(n_1632)
);

AOI33xp33_ASAP7_75t_L g1633 ( 
.A1(n_1623),
.A2(n_1509),
.A3(n_1507),
.B1(n_1518),
.B2(n_1519),
.B3(n_1561),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1624),
.B(n_1476),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_SL g1635 ( 
.A(n_1629),
.B(n_1507),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1631),
.A2(n_1630),
.B1(n_1628),
.B2(n_1519),
.C(n_1554),
.Y(n_1636)
);

OAI222xp33_ASAP7_75t_L g1637 ( 
.A1(n_1634),
.A2(n_1450),
.B1(n_1554),
.B2(n_1550),
.C1(n_1549),
.C2(n_1561),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1635),
.Y(n_1638)
);

XNOR2xp5_ASAP7_75t_L g1639 ( 
.A(n_1632),
.B(n_1342),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1633),
.A2(n_1550),
.B1(n_1549),
.B2(n_1347),
.C(n_1521),
.Y(n_1640)
);

AO21x1_ASAP7_75t_L g1641 ( 
.A1(n_1635),
.A2(n_1529),
.B(n_1442),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1638),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1637),
.B(n_1351),
.Y(n_1643)
);

NAND2x1p5_ASAP7_75t_SL g1644 ( 
.A(n_1636),
.B(n_1311),
.Y(n_1644)
);

OA211x2_ASAP7_75t_L g1645 ( 
.A1(n_1640),
.A2(n_1387),
.B(n_1380),
.C(n_1358),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1639),
.A2(n_1465),
.B1(n_1477),
.B2(n_1481),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1643),
.B(n_1641),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_L g1648 ( 
.A(n_1642),
.B(n_1382),
.C(n_1390),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1644),
.B(n_1382),
.C(n_1351),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1649),
.A2(n_1645),
.B1(n_1646),
.B2(n_1478),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1650),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1651),
.B(n_1647),
.Y(n_1652)
);

OAI22x1_ASAP7_75t_L g1653 ( 
.A1(n_1651),
.A2(n_1648),
.B1(n_1382),
.B2(n_1445),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1652),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1653),
.B(n_1358),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1654),
.A2(n_1655),
.B(n_1401),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1654),
.A2(n_1475),
.B1(n_1481),
.B2(n_1478),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1656),
.B(n_1358),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1658),
.Y(n_1659)
);

XNOR2xp5_ASAP7_75t_L g1660 ( 
.A(n_1659),
.B(n_1657),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1660),
.A2(n_1442),
.B1(n_1481),
.B2(n_1478),
.C(n_1477),
.Y(n_1661)
);

AOI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1319),
.B(n_1311),
.C(n_1379),
.Y(n_1662)
);


endmodule