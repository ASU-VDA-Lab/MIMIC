module fake_jpeg_8034_n_81 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_2),
.Y(n_47)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_2),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_3),
.B(n_9),
.Y(n_49)
);

NAND5xp2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_51),
.C(n_52),
.D(n_53),
.E(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_10),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_14),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_16),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_64),
.B1(n_41),
.B2(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_43),
.B1(n_44),
.B2(n_34),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_67),
.B(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_65),
.B1(n_52),
.B2(n_58),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_58),
.B(n_33),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_25),
.B1(n_57),
.B2(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_70),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_25),
.B1(n_38),
.B2(n_42),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_35),
.B(n_37),
.Y(n_76)
);

OAI31xp33_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_77),
.A3(n_24),
.B(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_28),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_18),
.B(n_21),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_35),
.C(n_55),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_35),
.B(n_45),
.Y(n_81)
);


endmodule