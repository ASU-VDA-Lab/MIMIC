module fake_jpeg_26905_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_28),
.B1(n_25),
.B2(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_28),
.B1(n_32),
.B2(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_48),
.B1(n_54),
.B2(n_36),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_17),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_22),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_28),
.B1(n_32),
.B2(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_18),
.B1(n_35),
.B2(n_40),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_39),
.B1(n_38),
.B2(n_34),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_77),
.B1(n_80),
.B2(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_59),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_62),
.Y(n_108)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_65),
.B(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_74),
.B1(n_76),
.B2(n_52),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_34),
.B(n_18),
.C(n_24),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_78),
.B(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_40),
.B1(n_17),
.B2(n_31),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_17),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_101),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_99),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_100),
.B1(n_102),
.B2(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_21),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_52),
.B1(n_21),
.B2(n_19),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_21),
.B1(n_19),
.B2(n_30),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_21),
.B1(n_19),
.B2(n_30),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_30),
.B(n_3),
.C(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_2),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_79),
.C(n_78),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_93),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_71),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_117),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_78),
.C(n_74),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.C(n_89),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_83),
.C(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_132),
.B1(n_128),
.B2(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_91),
.B(n_112),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_85),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_141),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_98),
.B1(n_89),
.B2(n_91),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_109),
.B1(n_123),
.B2(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_147),
.C(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_89),
.B1(n_92),
.B2(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_88),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_122),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_154),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_88),
.A3(n_104),
.B1(n_107),
.B2(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_66),
.B1(n_86),
.B2(n_94),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_158),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_165),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_118),
.A3(n_114),
.B1(n_115),
.B2(n_121),
.C1(n_110),
.C2(n_109),
.Y(n_162)
);

OAI322xp33_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_166),
.A3(n_169),
.B1(n_163),
.B2(n_167),
.C1(n_152),
.C2(n_139),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_113),
.B(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_117),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_94),
.C(n_130),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_149),
.C(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_126),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_141),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_177),
.C(n_178),
.Y(n_189)
);

AOI31xp33_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_164),
.A3(n_158),
.B(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_180),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_153),
.C(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_81),
.C(n_67),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_146),
.B1(n_84),
.B2(n_30),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_165),
.B1(n_168),
.B2(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_146),
.C(n_14),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_190),
.B1(n_13),
.B2(n_11),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_169),
.B1(n_168),
.B2(n_157),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_9),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_170),
.B1(n_161),
.B2(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_176),
.B1(n_181),
.B2(n_183),
.Y(n_191)
);

OAI31xp33_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_192)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_4),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_9),
.B(n_11),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_5),
.B(n_6),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_11),
.C(n_12),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_173),
.C(n_14),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_5),
.C(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_201),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_9),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_193),
.B(n_196),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_188),
.C(n_194),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g205 ( 
.A(n_192),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_12),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_199),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_211),
.B1(n_198),
.B2(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_197),
.C(n_198),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_216),
.B(n_209),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_12),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_215),
.C(n_214),
.Y(n_220)
);

NOR4xp25_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.C(n_219),
.D(n_13),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_13),
.Y(n_223)
);


endmodule