module fake_jpeg_26679_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.Y(n_32)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_26),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_13),
.B(n_18),
.C(n_16),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_40),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_25),
.B(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_20),
.Y(n_43)
);

OA22x2_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_27),
.B1(n_23),
.B2(n_14),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_48),
.B1(n_23),
.B2(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_37),
.C(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_34),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_42),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_57),
.C(n_10),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_45),
.B1(n_48),
.B2(n_39),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_62),
.B1(n_50),
.B2(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_15),
.Y(n_70)
);

NOR4xp25_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.C(n_28),
.D(n_19),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_21),
.B1(n_19),
.B2(n_11),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_15),
.B(n_10),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_20),
.B1(n_17),
.B2(n_15),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_29),
.C(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_19),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_72),
.B(n_75),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_73),
.B(n_58),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_R g80 ( 
.A(n_71),
.B(n_53),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_60),
.B(n_49),
.C(n_55),
.D(n_50),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_66),
.B(n_73),
.C(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_59),
.C(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_1),
.C(n_3),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_64),
.B1(n_81),
.B2(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_84),
.B1(n_68),
.B2(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_82),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_94),
.C(n_7),
.Y(n_99)
);

AOI31xp33_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_3),
.A3(n_6),
.B(n_7),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_87),
.A3(n_88),
.B1(n_5),
.B2(n_6),
.C1(n_1),
.C2(n_8),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_98),
.B(n_6),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_8),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_101),
.C(n_102),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

OA21x2_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_9),
.B(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_101),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_104),
.Y(n_107)
);


endmodule