module fake_jpeg_29388_n_467 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_49),
.Y(n_149)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g154 ( 
.A(n_55),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_7),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_79),
.Y(n_113)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_24),
.B(n_7),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_34),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_89),
.Y(n_140)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_8),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_34),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_95),
.Y(n_122)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_98),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_102),
.B(n_120),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_27),
.B1(n_29),
.B2(n_45),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_104),
.A2(n_110),
.B1(n_142),
.B2(n_147),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_59),
.A2(n_27),
.B1(n_29),
.B2(n_45),
.Y(n_110)
);

BUFx2_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_23),
.B(n_43),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_128),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_60),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_61),
.A2(n_97),
.B1(n_56),
.B2(n_52),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_128),
.B1(n_132),
.B2(n_136),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_41),
.B1(n_27),
.B2(n_46),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_51),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_73),
.A2(n_39),
.B1(n_20),
.B2(n_35),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_18),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_155),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_45),
.B1(n_53),
.B2(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_77),
.A2(n_98),
.B1(n_96),
.B2(n_84),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_78),
.A2(n_39),
.B1(n_35),
.B2(n_33),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_44),
.B1(n_48),
.B2(n_47),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_49),
.B(n_33),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_83),
.B1(n_82),
.B2(n_81),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_157),
.A2(n_174),
.B1(n_141),
.B2(n_100),
.Y(n_239)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_159),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_163),
.Y(n_225)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_183),
.B1(n_201),
.B2(n_110),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_176),
.Y(n_220)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_95),
.B1(n_72),
.B2(n_48),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_113),
.B(n_47),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_177),
.Y(n_227)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_140),
.B(n_44),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_181),
.B(n_198),
.Y(n_221)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_184),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_102),
.A2(n_43),
.B1(n_23),
.B2(n_38),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_187),
.Y(n_243)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_38),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_129),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_154),
.A2(n_45),
.B1(n_43),
.B2(n_38),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_217)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_154),
.A2(n_45),
.B1(n_38),
.B2(n_32),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_103),
.A2(n_38),
.B1(n_32),
.B2(n_9),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_125),
.A2(n_38),
.B1(n_9),
.B2(n_10),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_100),
.B1(n_144),
.B2(n_115),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

OA22x2_ASAP7_75t_SL g201 ( 
.A1(n_104),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_205),
.B1(n_152),
.B2(n_99),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_206),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_208),
.A2(n_218),
.B1(n_158),
.B2(n_182),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_122),
.B(n_143),
.C(n_150),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_233),
.B(n_200),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_108),
.B(n_103),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_173),
.B(n_180),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_214),
.Y(n_252)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_142),
.A3(n_152),
.B1(n_127),
.B2(n_126),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_161),
.B1(n_165),
.B2(n_157),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_126),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_222),
.B(n_185),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_144),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_241),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_124),
.B(n_127),
.C(n_139),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_124),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_203),
.C(n_195),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_141),
.B1(n_107),
.B2(n_160),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_153),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_115),
.B1(n_107),
.B2(n_99),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_187),
.B1(n_204),
.B2(n_162),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_201),
.B(n_183),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_244),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_231),
.A2(n_177),
.B1(n_179),
.B2(n_169),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_248),
.A2(n_258),
.B1(n_217),
.B2(n_229),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_266),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_164),
.B1(n_191),
.B2(n_199),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_251),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_213),
.Y(n_289)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_192),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_263),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_261),
.B(n_262),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_220),
.B(n_10),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_267),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_171),
.B1(n_32),
.B2(n_2),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_0),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_32),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_269),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_6),
.B1(n_14),
.B2(n_12),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_270),
.Y(n_288)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_206),
.B(n_1),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_10),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_216),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_227),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_210),
.B1(n_227),
.B2(n_232),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_210),
.C(n_209),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_287),
.B(n_276),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_247),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_255),
.A2(n_206),
.B1(n_214),
.B2(n_233),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_306),
.Y(n_326)
);

OAI22x1_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_258),
.B1(n_266),
.B2(n_249),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_252),
.A2(n_206),
.B(n_243),
.Y(n_293)
);

AO22x2_ASAP7_75t_L g319 ( 
.A1(n_293),
.A2(n_299),
.B1(n_245),
.B2(n_246),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_264),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_221),
.C(n_215),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_309),
.C(n_254),
.Y(n_311)
);

AOI22x1_ASAP7_75t_L g299 ( 
.A1(n_255),
.A2(n_251),
.B1(n_274),
.B2(n_252),
.Y(n_299)
);

BUFx24_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_301),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_274),
.A2(n_227),
.B1(n_235),
.B2(n_216),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_254),
.B(n_207),
.C(n_224),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_314),
.C(n_321),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_280),
.A2(n_251),
.B(n_257),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_312),
.A2(n_332),
.B(n_334),
.Y(n_362)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_260),
.C(n_247),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_304),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_317),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_267),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_330),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_337),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_300),
.A2(n_256),
.B1(n_258),
.B2(n_245),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_320),
.A2(n_329),
.B1(n_306),
.B2(n_279),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_260),
.C(n_267),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_268),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_336),
.C(n_338),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_225),
.Y(n_323)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_323),
.Y(n_353)
);

OA22x2_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_302),
.B1(n_293),
.B2(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_300),
.A2(n_256),
.B1(n_253),
.B2(n_248),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_263),
.B(n_248),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_278),
.B1(n_305),
.B2(n_303),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_281),
.A2(n_269),
.B(n_253),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_259),
.C(n_271),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_339),
.A2(n_340),
.B1(n_345),
.B2(n_348),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_284),
.B1(n_279),
.B2(n_293),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_302),
.B1(n_308),
.B2(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_342),
.B(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_299),
.B1(n_250),
.B2(n_282),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_304),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_324),
.A2(n_299),
.B1(n_282),
.B2(n_288),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_288),
.B1(n_308),
.B2(n_305),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_350),
.A2(n_321),
.B1(n_319),
.B2(n_310),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_351),
.B(n_356),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_326),
.A2(n_303),
.B1(n_297),
.B2(n_307),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_354),
.A2(n_358),
.B1(n_328),
.B2(n_334),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_265),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_277),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_361),
.Y(n_375)
);

AO22x1_ASAP7_75t_SL g360 ( 
.A1(n_319),
.A2(n_301),
.B1(n_235),
.B2(n_232),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_332),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_275),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_270),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_236),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_347),
.C(n_363),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_370),
.C(n_374),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_369),
.A2(n_371),
.B1(n_340),
.B2(n_344),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_327),
.C(n_314),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_354),
.A2(n_327),
.B1(n_336),
.B2(n_312),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_378),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_338),
.C(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_362),
.A2(n_319),
.B(n_326),
.C(n_337),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_380),
.A2(n_387),
.B(n_360),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_381),
.A2(n_339),
.B1(n_345),
.B2(n_361),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_319),
.C(n_310),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_357),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_388),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_348),
.Y(n_384)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_342),
.B(n_301),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_385),
.B(n_357),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_225),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_386),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_301),
.B(n_212),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_236),
.Y(n_388)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_390),
.A2(n_398),
.B1(n_406),
.B2(n_371),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_393),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_387),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_385),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_374),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_367),
.A2(n_344),
.B1(n_349),
.B2(n_346),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_397),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_344),
.B1(n_365),
.B2(n_232),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_403),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_207),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_224),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_372),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_372),
.B1(n_381),
.B2(n_384),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_408),
.A2(n_396),
.B1(n_400),
.B2(n_392),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_414),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_399),
.B(n_382),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_411),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_368),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_398),
.A2(n_376),
.B1(n_380),
.B2(n_370),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_418),
.B1(n_410),
.B2(n_408),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_390),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_366),
.C(n_375),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_419),
.C(n_421),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_405),
.B(n_375),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_366),
.C(n_212),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_228),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_417),
.C(n_419),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_423),
.B(n_427),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_424),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_413),
.B(n_393),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_426),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_406),
.C(n_396),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_420),
.A2(n_400),
.B(n_401),
.Y(n_428)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_428),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_431),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_401),
.C(n_404),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_389),
.C(n_240),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_238),
.C(n_228),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_420),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_438),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_407),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_443),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_414),
.Y(n_441)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_441),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_238),
.C(n_228),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_6),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_2),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_425),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_451),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_430),
.C(n_12),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_450),
.B(n_449),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_436),
.A2(n_6),
.B(n_14),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_452),
.A2(n_441),
.B(n_442),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_SL g453 ( 
.A1(n_442),
.A2(n_14),
.B(n_15),
.C(n_3),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_455),
.A2(n_456),
.B(n_15),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_435),
.B(n_447),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g460 ( 
.A1(n_458),
.A2(n_453),
.B(n_15),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_SL g459 ( 
.A1(n_457),
.A2(n_453),
.B(n_438),
.C(n_439),
.Y(n_459)
);

AOI321xp33_ASAP7_75t_L g462 ( 
.A1(n_459),
.A2(n_461),
.A3(n_3),
.B1(n_4),
.B2(n_454),
.C(n_333),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_460),
.Y(n_463)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_462),
.A2(n_3),
.B(n_4),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_464),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_463),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_3),
.Y(n_467)
);


endmodule