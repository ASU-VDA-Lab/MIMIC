module fake_netlist_5_138_n_10281 (n_91, n_82, n_122, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_10281);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_10281;

wire n_924;
wire n_6643;
wire n_6122;
wire n_977;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_7981;
wire n_9936;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_9194;
wire n_3241;
wire n_3006;
wire n_6579;
wire n_532;
wire n_9325;
wire n_7164;
wire n_6546;
wire n_5287;
wire n_2327;
wire n_9655;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_8174;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_5207;
wire n_9044;
wire n_2347;
wire n_6786;
wire n_7206;
wire n_7303;
wire n_9083;
wire n_4963;
wire n_8363;
wire n_4508;
wire n_9408;
wire n_4240;
wire n_2021;
wire n_7710;
wire n_8383;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_551;
wire n_3615;
wire n_8328;
wire n_2059;
wire n_7461;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_6649;
wire n_8060;
wire n_9331;
wire n_7154;
wire n_8551;
wire n_3202;
wire n_8002;
wire n_4977;
wire n_3813;
wire n_10108;
wire n_8594;
wire n_6810;
wire n_7660;
wire n_671;
wire n_6276;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_8976;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_8617;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_7686;
wire n_4211;
wire n_10117;
wire n_9846;
wire n_8603;
wire n_7024;
wire n_3448;
wire n_7205;
wire n_9204;
wire n_6742;
wire n_9769;
wire n_3019;
wire n_2096;
wire n_9312;
wire n_8319;
wire n_6694;
wire n_877;
wire n_3776;
wire n_9610;
wire n_7616;
wire n_2530;
wire n_7486;
wire n_1696;
wire n_2483;
wire n_4517;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_8244;
wire n_9273;
wire n_1860;
wire n_4615;
wire n_1107;
wire n_2076;
wire n_1728;
wire n_6090;
wire n_6580;
wire n_7010;
wire n_5480;
wire n_6549;
wire n_8105;
wire n_668;
wire n_6913;
wire n_7867;
wire n_301;
wire n_2147;
wire n_3010;
wire n_7315;
wire n_7004;
wire n_8961;
wire n_2770;
wire n_4131;
wire n_7772;
wire n_5402;
wire n_2584;
wire n_171;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_9773;
wire n_8574;
wire n_3403;
wire n_3624;
wire n_8864;
wire n_3461;
wire n_9173;
wire n_3082;
wire n_7641;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_9363;
wire n_8681;
wire n_7468;
wire n_9796;
wire n_519;
wire n_5469;
wire n_2323;
wire n_6431;
wire n_5744;
wire n_2597;
wire n_9049;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_281;
wire n_7861;
wire n_2052;
wire n_9907;
wire n_4499;
wire n_4927;
wire n_8413;
wire n_9738;
wire n_731;
wire n_5202;
wire n_5648;
wire n_7667;
wire n_1314;
wire n_1512;
wire n_6931;
wire n_9539;
wire n_8114;
wire n_1490;
wire n_317;
wire n_9811;
wire n_6618;
wire n_6408;
wire n_9993;
wire n_569;
wire n_9208;
wire n_3214;
wire n_7523;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_8706;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_8158;
wire n_1449;
wire n_6698;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_297;
wire n_9500;
wire n_2587;
wire n_156;
wire n_8104;
wire n_5848;
wire n_5406;
wire n_219;
wire n_157;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_7421;
wire n_7306;
wire n_600;
wire n_8819;
wire n_223;
wire n_6214;
wire n_7493;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_9420;
wire n_7804;
wire n_8089;
wire n_9557;
wire n_3353;
wire n_264;
wire n_4203;
wire n_3687;
wire n_9382;
wire n_5241;
wire n_6939;
wire n_882;
wire n_2384;
wire n_7528;
wire n_3156;
wire n_8262;
wire n_8290;
wire n_9206;
wire n_696;
wire n_3376;
wire n_7562;
wire n_646;
wire n_5037;
wire n_9388;
wire n_10193;
wire n_436;
wire n_4468;
wire n_8885;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_5661;
wire n_9772;
wire n_3702;
wire n_1040;
wire n_8147;
wire n_6586;
wire n_2202;
wire n_2648;
wire n_4976;
wire n_5008;
wire n_2159;
wire n_10177;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_8310;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_2276;
wire n_6707;
wire n_10175;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_9311;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_9422;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_9040;
wire n_9795;
wire n_521;
wire n_8380;
wire n_845;
wire n_9027;
wire n_8962;
wire n_528;
wire n_7402;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_395;
wire n_553;
wire n_901;
wire n_4484;
wire n_7592;
wire n_3668;
wire n_7152;
wire n_6512;
wire n_9966;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_637;
wire n_8126;
wire n_5689;
wire n_144;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_7801;
wire n_7992;
wire n_1151;
wire n_9161;
wire n_10231;
wire n_1405;
wire n_7463;
wire n_1706;
wire n_3418;
wire n_8556;
wire n_342;
wire n_9369;
wire n_4901;
wire n_9033;
wire n_8305;
wire n_6725;
wire n_7613;
wire n_197;
wire n_2859;
wire n_1075;
wire n_9429;
wire n_3395;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_6464;
wire n_2863;
wire n_2072;
wire n_8317;
wire n_2738;
wire n_8653;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_2968;
wire n_7316;
wire n_1585;
wire n_6820;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_9780;
wire n_10252;
wire n_4421;
wire n_9824;
wire n_6098;
wire n_7019;
wire n_6686;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_10202;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_190;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_7956;
wire n_8939;
wire n_4532;
wire n_3339;
wire n_9489;
wire n_8604;
wire n_228;
wire n_283;
wire n_3349;
wire n_3735;
wire n_7323;
wire n_2248;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_3007;
wire n_1000;
wire n_6769;
wire n_7683;
wire n_6592;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_310;
wire n_3487;
wire n_3310;
wire n_6191;
wire n_6062;
wire n_7903;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_9625;
wire n_8440;
wire n_3983;
wire n_332;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_8525;
wire n_1331;
wire n_4195;
wire n_8416;
wire n_279;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_9570;
wire n_9368;
wire n_8064;
wire n_7575;
wire n_1385;
wire n_440;
wire n_5909;
wire n_793;
wire n_2776;
wire n_8879;
wire n_4408;
wire n_9115;
wire n_2140;
wire n_2385;
wire n_9367;
wire n_9694;
wire n_1819;
wire n_4531;
wire n_6043;
wire n_476;
wire n_2987;
wire n_1527;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_7701;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_345;
wire n_4130;
wire n_8931;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_8214;
wire n_9072;
wire n_6793;
wire n_7873;
wire n_2324;
wire n_9612;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_9971;
wire n_8729;
wire n_7127;
wire n_5397;
wire n_182;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_407;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_7568;
wire n_3208;
wire n_6021;
wire n_9720;
wire n_207;
wire n_3331;
wire n_2379;
wire n_5695;
wire n_7814;
wire n_4983;
wire n_9213;
wire n_2911;
wire n_10187;
wire n_2154;
wire n_4916;
wire n_6926;
wire n_5860;
wire n_3649;
wire n_9607;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_7965;
wire n_2514;
wire n_5862;
wire n_6304;
wire n_8228;
wire n_8210;
wire n_5189;
wire n_6956;
wire n_10040;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_1027;
wire n_326;
wire n_4160;
wire n_6782;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_9554;
wire n_9262;
wire n_2028;
wire n_558;
wire n_3009;
wire n_1276;
wire n_7002;
wire n_8387;
wire n_1412;
wire n_3981;
wire n_8898;
wire n_8410;
wire n_7141;
wire n_5936;
wire n_6126;
wire n_9761;
wire n_1199;
wire n_8795;
wire n_352;
wire n_9649;
wire n_10164;
wire n_10269;
wire n_8501;
wire n_1038;
wire n_520;
wire n_1841;
wire n_6598;
wire n_154;
wire n_6027;
wire n_9254;
wire n_9529;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_870;
wire n_1711;
wire n_6638;
wire n_1891;
wire n_7308;
wire n_5254;
wire n_434;
wire n_3526;
wire n_6900;
wire n_8953;
wire n_2546;
wire n_965;
wire n_9726;
wire n_8823;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_7457;
wire n_4613;
wire n_7718;
wire n_4649;
wire n_7617;
wire n_1888;
wire n_9197;
wire n_6269;
wire n_8843;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_7768;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_7974;
wire n_9106;
wire n_7357;
wire n_6013;
wire n_2449;
wire n_5083;
wire n_8247;
wire n_9564;
wire n_6927;
wire n_9627;
wire n_7975;
wire n_431;
wire n_1194;
wire n_6503;
wire n_5888;
wire n_8172;
wire n_2297;
wire n_4186;
wire n_8940;
wire n_8941;
wire n_7310;
wire n_9739;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_2227;
wire n_4618;
wire n_127;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_7593;
wire n_7716;
wire n_6256;
wire n_2876;
wire n_4099;
wire n_452;
wire n_7406;
wire n_7600;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_10223;
wire n_2479;
wire n_5870;
wire n_9812;
wire n_1464;
wire n_4295;
wire n_649;
wire n_9646;
wire n_5303;
wire n_1444;
wire n_10201;
wire n_7076;
wire n_8780;
wire n_10215;
wire n_9465;
wire n_9928;
wire n_4694;
wire n_8456;
wire n_9970;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_9894;
wire n_10100;
wire n_10278;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_9129;
wire n_3168;
wire n_6982;
wire n_1680;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_9957;
wire n_2607;
wire n_4190;
wire n_3994;
wire n_9558;
wire n_4810;
wire n_7848;
wire n_6727;
wire n_3317;
wire n_8218;
wire n_9267;
wire n_7539;
wire n_1121;
wire n_8769;
wire n_433;
wire n_7229;
wire n_4391;
wire n_949;
wire n_8514;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_8368;
wire n_4681;
wire n_8334;
wire n_1001;
wire n_1503;
wire n_9918;
wire n_4638;
wire n_1468;
wire n_8159;
wire n_3455;
wire n_6097;
wire n_8639;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_1195;
wire n_7797;
wire n_4707;
wire n_2577;
wire n_8216;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_2796;
wire n_757;
wire n_7869;
wire n_6466;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_9956;
wire n_4848;
wire n_9095;
wire n_9715;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_8337;
wire n_8257;
wire n_7983;
wire n_2805;
wire n_7781;
wire n_8125;
wire n_1145;
wire n_524;
wire n_5624;
wire n_394;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_1153;
wire n_3856;
wire n_9246;
wire n_741;
wire n_7624;
wire n_9683;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_1163;
wire n_8063;
wire n_9931;
wire n_6805;
wire n_6185;
wire n_1207;
wire n_5010;
wire n_7762;
wire n_8731;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_8950;
wire n_3918;
wire n_2398;
wire n_6568;
wire n_2857;
wire n_9011;
wire n_9899;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_8295;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_940;
wire n_6351;
wire n_7552;
wire n_8059;
wire n_3516;
wire n_4822;
wire n_8995;
wire n_2155;
wire n_8146;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_6901;
wire n_8082;
wire n_2947;
wire n_123;
wire n_9094;
wire n_978;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_6411;
wire n_3515;
wire n_8339;
wire n_2886;
wire n_267;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_9195;
wire n_3378;
wire n_7746;
wire n_5435;
wire n_1431;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_660;
wire n_8032;
wire n_7139;
wire n_8640;
wire n_4294;
wire n_9332;
wire n_10016;
wire n_1732;
wire n_10070;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_8351;
wire n_4949;
wire n_374;
wire n_10190;
wire n_2941;
wire n_8196;
wire n_6594;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_459;
wire n_7857;
wire n_962;
wire n_9054;
wire n_10150;
wire n_9460;
wire n_9638;
wire n_723;
wire n_2536;
wire n_6387;
wire n_1336;
wire n_7223;
wire n_1758;
wire n_7890;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_9281;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_10134;
wire n_7964;
wire n_5096;
wire n_9740;
wire n_4365;
wire n_9475;
wire n_8865;
wire n_9661;
wire n_1878;
wire n_6019;
wire n_9190;
wire n_6222;
wire n_7165;
wire n_8110;
wire n_3505;
wire n_6223;
wire n_8475;
wire n_8838;
wire n_4610;
wire n_6435;
wire n_9143;
wire n_3730;
wire n_4489;
wire n_7235;
wire n_168;
wire n_974;
wire n_727;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_8488;
wire n_5657;
wire n_957;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_8766;
wire n_6844;
wire n_3001;
wire n_7795;
wire n_8969;
wire n_303;
wire n_7404;
wire n_3945;
wire n_9891;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_6295;
wire n_3597;
wire n_9087;
wire n_9804;
wire n_8087;
wire n_8119;
wire n_1612;
wire n_10135;
wire n_9321;
wire n_7885;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_5857;
wire n_8173;
wire n_4534;
wire n_4500;
wire n_9800;
wire n_7437;
wire n_5014;
wire n_6241;
wire n_8420;
wire n_3185;
wire n_1300;
wire n_6087;
wire n_1127;
wire n_8019;
wire n_9186;
wire n_3523;
wire n_9951;
wire n_1785;
wire n_2829;
wire n_6846;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_9243;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_7822;
wire n_6041;
wire n_2017;
wire n_2604;
wire n_8851;
wire n_6994;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_322;
wire n_7329;
wire n_2390;
wire n_9359;
wire n_5708;
wire n_3213;
wire n_8687;
wire n_6790;
wire n_10001;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_383;
wire n_7194;
wire n_6273;
wire n_3474;
wire n_8740;
wire n_3984;
wire n_6807;
wire n_239;
wire n_630;
wire n_5927;
wire n_2151;
wire n_10189;
wire n_2106;
wire n_9879;
wire n_2716;
wire n_4665;
wire n_8221;
wire n_1913;
wire n_8468;
wire n_7708;
wire n_1823;
wire n_7696;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_9975;
wire n_7115;
wire n_9335;
wire n_4189;
wire n_5670;
wire n_9171;
wire n_1875;
wire n_8815;
wire n_1304;
wire n_9942;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_8952;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_9247;
wire n_9933;
wire n_5965;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_7958;
wire n_10209;
wire n_429;
wire n_8128;
wire n_4687;
wire n_948;
wire n_5751;
wire n_5664;
wire n_9441;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_8667;
wire n_4037;
wire n_6218;
wire n_8863;
wire n_7281;
wire n_10233;
wire n_2922;
wire n_3499;
wire n_3275;
wire n_2645;
wire n_8106;
wire n_9362;
wire n_2727;
wire n_560;
wire n_340;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_6824;
wire n_8717;
wire n_1552;
wire n_6189;
wire n_3618;
wire n_574;
wire n_2593;
wire n_9216;
wire n_8299;
wire n_5262;
wire n_9200;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_824;
wire n_8892;
wire n_359;
wire n_1327;
wire n_10146;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_9067;
wire n_5310;
wire n_366;
wire n_9152;
wire n_8287;
wire n_815;
wire n_4594;
wire n_6153;
wire n_9074;
wire n_7989;
wire n_3424;
wire n_5970;
wire n_1381;
wire n_6418;
wire n_1037;
wire n_6564;
wire n_2301;
wire n_3583;
wire n_8657;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_589;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_9287;
wire n_4102;
wire n_8197;
wire n_9511;
wire n_10052;
wire n_2786;
wire n_8081;
wire n_7192;
wire n_3171;
wire n_6671;
wire n_1437;
wire n_645;
wire n_6591;
wire n_238;
wire n_6266;
wire n_7161;
wire n_7580;
wire n_7153;
wire n_9880;
wire n_10072;
wire n_9843;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_8609;
wire n_3462;
wire n_5441;
wire n_6517;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_222;
wire n_8559;
wire n_7350;
wire n_5690;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_634;
wire n_6967;
wire n_5885;
wire n_9248;
wire n_2254;
wire n_6433;
wire n_1382;
wire n_925;
wire n_3546;
wire n_7535;
wire n_6893;
wire n_424;
wire n_2647;
wire n_9128;
wire n_1311;
wire n_8452;
wire n_1519;
wire n_256;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_10224;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_7632;
wire n_8771;
wire n_380;
wire n_419;
wire n_8140;
wire n_8476;
wire n_9528;
wire n_3244;
wire n_6501;
wire n_8981;
wire n_10157;
wire n_9507;
wire n_6028;
wire n_389;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_136;
wire n_968;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_619;
wire n_9533;
wire n_5362;
wire n_376;
wire n_8137;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_8469;
wire n_515;
wire n_6798;
wire n_351;
wire n_5702;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_7844;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_683;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_9665;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_8423;
wire n_5527;
wire n_6986;
wire n_802;
wire n_8090;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_280;
wire n_1305;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_873;
wire n_9436;
wire n_5355;
wire n_2334;
wire n_9562;
wire n_6745;
wire n_690;
wire n_8260;
wire n_4521;
wire n_8481;
wire n_583;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_2289;
wire n_3051;
wire n_302;
wire n_1343;
wire n_2783;
wire n_6209;
wire n_2263;
wire n_6875;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_7905;
wire n_212;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_5551;
wire n_7766;
wire n_7594;
wire n_3715;
wire n_7803;
wire n_7340;
wire n_6699;
wire n_7747;
wire n_6073;
wire n_972;
wire n_8205;
wire n_5767;
wire n_8401;
wire n_6324;
wire n_3040;
wire n_8651;
wire n_1938;
wire n_5640;
wire n_1200;
wire n_2499;
wire n_10199;
wire n_8284;
wire n_3568;
wire n_9255;
wire n_10039;
wire n_8828;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_6138;
wire n_7603;
wire n_8510;
wire n_1967;
wire n_8810;
wire n_576;
wire n_9034;
wire n_1329;
wire n_3255;
wire n_9203;
wire n_9601;
wire n_5692;
wire n_4856;
wire n_7726;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_8024;
wire n_9946;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_9967;
wire n_6477;
wire n_10274;
wire n_8739;
wire n_3734;
wire n_650;
wire n_8133;
wire n_8373;
wire n_8919;
wire n_4778;
wire n_286;
wire n_2429;
wire n_883;
wire n_6159;
wire n_9647;
wire n_6283;
wire n_7396;
wire n_470;
wire n_9912;
wire n_325;
wire n_132;
wire n_5322;
wire n_856;
wire n_7116;
wire n_1793;
wire n_4352;
wire n_7519;
wire n_4441;
wire n_6943;
wire n_9329;
wire n_918;
wire n_6827;
wire n_4761;
wire n_6173;
wire n_8318;
wire n_942;
wire n_1804;
wire n_189;
wire n_8542;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_8543;
wire n_8846;
wire n_4593;
wire n_6312;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_195;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_7770;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_7664;
wire n_5316;
wire n_9890;
wire n_3831;
wire n_10273;
wire n_3801;
wire n_6300;
wire n_225;
wire n_9609;
wire n_9883;
wire n_10172;
wire n_7815;
wire n_2043;
wire n_9046;
wire n_2751;
wire n_9361;
wire n_8163;
wire n_192;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_6537;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_655;
wire n_9864;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_472;
wire n_7023;
wire n_8972;
wire n_9300;
wire n_1807;
wire n_387;
wire n_2618;
wire n_398;
wire n_7428;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_6783;
wire n_9353;
wire n_4748;
wire n_9766;
wire n_7465;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_8293;
wire n_2840;
wire n_5017;
wire n_9832;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_287;
wire n_555;
wire n_4607;
wire n_5123;
wire n_9954;
wire n_4117;
wire n_8737;
wire n_3636;
wire n_7961;
wire n_1722;
wire n_7847;
wire n_9997;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_9334;
wire n_7149;
wire n_2795;
wire n_8252;
wire n_6459;
wire n_9622;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_8450;
wire n_4817;
wire n_7700;
wire n_9284;
wire n_311;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_9147;
wire n_8367;
wire n_3538;
wire n_10103;
wire n_8834;
wire n_6869;
wire n_8078;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_7914;
wire n_445;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_7967;
wire n_9794;
wire n_4728;
wire n_7117;
wire n_588;
wire n_789;
wire n_9354;
wire n_8471;
wire n_4247;
wire n_4933;
wire n_6977;
wire n_4018;
wire n_8474;
wire n_3900;
wire n_7984;
wire n_1105;
wire n_10185;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_8361;
wire n_6313;
wire n_3872;
wire n_4336;
wire n_6569;
wire n_149;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_9494;
wire n_6555;
wire n_9614;
wire n_9551;
wire n_3877;
wire n_458;
wire n_6639;
wire n_7516;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_9154;
wire n_1102;
wire n_7596;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_8553;
wire n_6490;
wire n_8301;
wire n_2633;
wire n_6961;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_9437;
wire n_1164;
wire n_2097;
wire n_5460;
wire n_7628;
wire n_9276;
wire n_4304;
wire n_6761;
wire n_9346;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_6294;
wire n_6767;
wire n_8518;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_9514;
wire n_4805;
wire n_9402;
wire n_601;
wire n_4885;
wire n_7838;
wire n_8364;
wire n_7786;
wire n_5983;
wire n_9580;
wire n_253;
wire n_9005;
wire n_1661;
wire n_5804;
wire n_7979;
wire n_6376;
wire n_3565;
wire n_172;
wire n_6167;
wire n_8621;
wire n_8993;
wire n_7926;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_9162;
wire n_9921;
wire n_9443;
wire n_861;
wire n_6582;
wire n_1658;
wire n_8910;
wire n_7752;
wire n_1904;
wire n_9897;
wire n_6996;
wire n_9817;
wire n_1345;
wire n_176;
wire n_9301;
wire n_1899;
wire n_6974;
wire n_7731;
wire n_8753;
wire n_6765;
wire n_7577;
wire n_8388;
wire n_9401;
wire n_8321;
wire n_1003;
wire n_6921;
wire n_2067;
wire n_8044;
wire n_8091;
wire n_2219;
wire n_8486;
wire n_7845;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_393;
wire n_7709;
wire n_9689;
wire n_4631;
wire n_1726;
wire n_3035;
wire n_421;
wire n_5194;
wire n_9982;
wire n_6898;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_8508;
wire n_8261;
wire n_1657;
wire n_5886;
wire n_768;
wire n_7080;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_7744;
wire n_1491;
wire n_754;
wire n_9886;
wire n_8034;
wire n_8841;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_10264;
wire n_6960;
wire n_8201;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_1915;
wire n_5610;
wire n_1109;
wire n_5239;
wire n_6836;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_8947;
wire n_1399;
wire n_9671;
wire n_1979;
wire n_6972;
wire n_193;
wire n_2924;
wire n_9297;
wire n_8788;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_5785;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_6093;
wire n_8093;
wire n_435;
wire n_766;
wire n_541;
wire n_6010;
wire n_7247;
wire n_9225;
wire n_8061;
wire n_1117;
wire n_6833;
wire n_2754;
wire n_687;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_536;
wire n_7481;
wire n_10066;
wire n_5204;
wire n_7292;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_8811;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_7687;
wire n_1155;
wire n_1418;
wire n_10184;
wire n_1011;
wire n_8507;
wire n_9662;
wire n_2917;
wire n_9057;
wire n_2425;
wire n_3661;
wire n_3536;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_6265;
wire n_8861;
wire n_1650;
wire n_1137;
wire n_6821;
wire n_8661;
wire n_3934;
wire n_8545;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_8755;
wire n_5788;
wire n_8573;
wire n_8191;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_318;
wire n_5897;
wire n_6887;
wire n_2103;
wire n_653;
wire n_9809;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_8683;
wire n_10081;
wire n_1999;
wire n_8836;
wire n_6676;
wire n_2372;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_9448;
wire n_3943;
wire n_353;
wire n_8136;
wire n_8446;
wire n_9799;
wire n_2430;
wire n_7742;
wire n_9313;
wire n_493;
wire n_8916;
wire n_2433;
wire n_3293;
wire n_7955;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_10037;
wire n_5582;
wire n_10234;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_9989;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_7758;
wire n_7547;
wire n_2528;
wire n_4869;
wire n_9438;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_10036;
wire n_554;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_6648;
wire n_7880;
wire n_4601;
wire n_8075;
wire n_2687;
wire n_1120;
wire n_8857;
wire n_198;
wire n_1890;
wire n_714;
wire n_4220;
wire n_8587;
wire n_9675;
wire n_10030;
wire n_1944;
wire n_909;
wire n_5630;
wire n_1497;
wire n_9667;
wire n_8071;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_7513;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_9537;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_1981;
wire n_7540;
wire n_8646;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_9866;
wire n_5504;
wire n_8630;
wire n_7622;
wire n_9602;
wire n_509;
wire n_7005;
wire n_147;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_7353;
wire n_6219;
wire n_10071;
wire n_9885;
wire n_1889;
wire n_209;
wire n_8315;
wire n_6965;
wire n_9260;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_8314;
wire n_6720;
wire n_1569;
wire n_8149;
wire n_2188;
wire n_6032;
wire n_186;
wire n_8581;
wire n_7174;
wire n_8565;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_756;
wire n_1429;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_7607;
wire n_8209;
wire n_9159;
wire n_399;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_7816;
wire n_9654;
wire n_3170;
wire n_8560;
wire n_7591;
wire n_5775;
wire n_8141;
wire n_2748;
wire n_3311;
wire n_7830;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_8302;
wire n_10015;
wire n_9306;
wire n_2898;
wire n_2717;
wire n_7151;
wire n_6229;
wire n_1861;
wire n_9978;
wire n_760;
wire n_5731;
wire n_8612;
wire n_5581;
wire n_3691;
wire n_3628;
wire n_6668;
wire n_7446;
wire n_220;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_481;
wire n_7053;
wire n_8724;
wire n_5831;
wire n_10171;
wire n_2573;
wire n_7473;
wire n_4435;
wire n_10183;
wire n_2939;
wire n_8070;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_271;
wire n_9279;
wire n_8457;
wire n_2447;
wire n_4764;
wire n_886;
wire n_5653;
wire n_8922;
wire n_8248;
wire n_7966;
wire n_9509;
wire n_6258;
wire n_10095;
wire n_7070;
wire n_1221;
wire n_5394;
wire n_167;
wire n_6755;
wire n_2774;
wire n_9563;
wire n_7276;
wire n_7351;
wire n_1707;
wire n_7942;
wire n_853;
wire n_10057;
wire n_4655;
wire n_3161;
wire n_377;
wire n_4581;
wire n_751;
wire n_6084;
wire n_4827;
wire n_9496;
wire n_8411;
wire n_9644;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_2488;
wire n_7666;
wire n_392;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_8527;
wire n_2476;
wire n_704;
wire n_7211;
wire n_10154;
wire n_4399;
wire n_6531;
wire n_2781;
wire n_5309;
wire n_7901;
wire n_8689;
wire n_9750;
wire n_2778;
wire n_771;
wire n_4782;
wire n_9980;
wire n_8988;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_9251;
wire n_10141;
wire n_2691;
wire n_7368;
wire n_1411;
wire n_8549;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_6771;
wire n_10208;
wire n_2526;
wire n_6389;
wire n_10182;
wire n_9616;
wire n_2703;
wire n_8004;
wire n_2167;
wire n_8658;
wire n_9959;
wire n_8375;
wire n_5764;
wire n_10260;
wire n_6910;
wire n_9291;
wire n_5428;
wire n_9092;
wire n_10261;
wire n_6442;
wire n_3391;
wire n_6102;
wire n_8908;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_6441;
wire n_5543;
wire n_816;
wire n_9818;
wire n_10237;
wire n_9283;
wire n_5678;
wire n_5935;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_7677;
wire n_5085;
wire n_3518;
wire n_8569;
wire n_2956;
wire n_3733;
wire n_328;
wire n_8676;
wire n_10118;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_871;
wire n_7929;
wire n_10028;
wire n_3738;
wire n_685;
wire n_8399;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_6331;
wire n_1555;
wire n_6006;
wire n_8421;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_499;
wire n_6278;
wire n_9304;
wire n_6787;
wire n_402;
wire n_6872;
wire n_6208;
wire n_796;
wire n_4899;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_6632;
wire n_9310;
wire n_1012;
wire n_7754;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_9830;
wire n_9913;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_8001;
wire n_5671;
wire n_3076;
wire n_8322;
wire n_6990;
wire n_8403;
wire n_3535;
wire n_2182;
wire n_6349;
wire n_277;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_7631;
wire n_6830;
wire n_8999;
wire n_8754;
wire n_5185;
wire n_7939;
wire n_8675;
wire n_7898;
wire n_1193;
wire n_6359;
wire n_9375;
wire n_3118;
wire n_8596;
wire n_10073;
wire n_3511;
wire n_8858;
wire n_1226;
wire n_8666;
wire n_3443;
wire n_8313;
wire n_2146;
wire n_7763;
wire n_1487;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_781;
wire n_542;
wire n_3521;
wire n_8555;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_6301;
wire n_2918;
wire n_3232;
wire n_8610;
wire n_1673;
wire n_7945;
wire n_5945;
wire n_2112;
wire n_1739;
wire n_9323;
wire n_2958;
wire n_6744;
wire n_3114;
wire n_3125;
wire n_4981;
wire n_9985;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_8615;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_10026;
wire n_8677;
wire n_9355;
wire n_8602;
wire n_9714;
wire n_7381;
wire n_10041;
wire n_5565;
wire n_4081;
wire n_1103;
wire n_7948;
wire n_3132;
wire n_4407;
wire n_648;
wire n_7291;
wire n_8102;
wire n_312;
wire n_9540;
wire n_3951;
wire n_4894;
wire n_9753;
wire n_5780;
wire n_8460;
wire n_9105;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_10149;
wire n_5846;
wire n_2036;
wire n_7430;
wire n_9700;
wire n_3267;
wire n_4995;
wire n_8871;
wire n_480;
wire n_425;
wire n_9476;
wire n_7870;
wire n_695;
wire n_9875;
wire n_5524;
wire n_8824;
wire n_3964;
wire n_3772;
wire n_229;
wire n_1956;
wire n_9963;
wire n_437;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_6104;
wire n_3884;
wire n_6475;
wire n_8470;
wire n_9582;
wire n_6465;
wire n_10060;
wire n_9574;
wire n_3726;
wire n_6496;
wire n_805;
wire n_2525;
wire n_9732;
wire n_2892;
wire n_2907;
wire n_8238;
wire n_9882;
wire n_6998;
wire n_6145;
wire n_3577;
wire n_8699;
wire n_2820;
wire n_269;
wire n_7305;
wire n_2049;
wire n_10242;
wire n_2273;
wire n_10086;
wire n_9992;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_7980;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_7075;
wire n_7545;
wire n_7846;
wire n_1448;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_8438;
wire n_6194;
wire n_7695;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_8095;
wire n_7537;
wire n_3212;
wire n_666;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_10128;
wire n_7489;
wire n_5106;
wire n_319;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_8112;
wire n_1186;
wire n_5883;
wire n_6985;
wire n_8642;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_7451;
wire n_8624;
wire n_6238;
wire n_713;
wire n_9090;
wire n_1622;
wire n_166;
wire n_1180;
wire n_9149;
wire n_9174;
wire n_3705;
wire n_6548;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_8894;
wire n_2268;
wire n_9226;
wire n_3778;
wire n_6366;
wire n_5706;
wire n_9018;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_7236;
wire n_9835;
wire n_2739;
wire n_469;
wire n_2771;
wire n_4604;
wire n_7269;
wire n_8878;
wire n_549;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_9702;
wire n_3256;
wire n_7560;
wire n_10279;
wire n_667;
wire n_7326;
wire n_7060;
wire n_2386;
wire n_1501;
wire n_7572;
wire n_3086;
wire n_1007;
wire n_6885;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_8807;
wire n_2821;
wire n_9968;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_9924;
wire n_564;
wire n_6529;
wire n_8732;
wire n_8169;
wire n_1738;
wire n_3728;
wire n_8803;
wire n_3064;
wire n_9515;
wire n_3088;
wire n_1021;
wire n_8017;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_8801;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_6423;
wire n_9252;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_7140;
wire n_7233;
wire n_10228;
wire n_819;
wire n_5088;
wire n_2302;
wire n_6558;
wire n_8522;
wire n_5457;
wire n_7352;
wire n_951;
wire n_7986;
wire n_9948;
wire n_7134;
wire n_5532;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_2069;
wire n_6950;
wire n_7246;
wire n_417;
wire n_7650;
wire n_6525;
wire n_3434;
wire n_9871;
wire n_1806;
wire n_933;
wire n_6631;
wire n_6892;
wire n_8203;
wire n_1563;
wire n_7663;
wire n_9423;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_9660;
wire n_9108;
wire n_2024;
wire n_4780;
wire n_8680;
wire n_9631;
wire n_755;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_530;
wire n_4330;
wire n_3695;
wire n_6683;
wire n_556;
wire n_8727;
wire n_2482;
wire n_2677;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_9900;
wire n_7729;
wire n_3987;
wire n_7339;
wire n_902;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_8138;
wire n_6658;
wire n_6264;
wire n_9608;
wire n_9137;
wire n_6925;
wire n_8990;
wire n_5919;
wire n_579;
wire n_1698;
wire n_10077;
wire n_2329;
wire n_8206;
wire n_1098;
wire n_9144;
wire n_2142;
wire n_7767;
wire n_8190;
wire n_6176;
wire n_9778;
wire n_8622;
wire n_320;
wire n_5410;
wire n_3332;
wire n_7146;
wire n_1135;
wire n_8092;
wire n_3048;
wire n_3937;
wire n_10250;
wire n_6124;
wire n_7672;
wire n_2203;
wire n_8242;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_7482;
wire n_9850;
wire n_6864;
wire n_9531;
wire n_7893;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_8331;
wire n_4208;
wire n_7090;
wire n_3786;
wire n_7158;
wire n_371;
wire n_2888;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_8649;
wire n_8684;
wire n_6494;
wire n_5503;
wire n_8323;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_6199;
wire n_8296;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_9139;
wire n_2306;
wire n_9430;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_3022;
wire n_7839;
wire n_4264;
wire n_8882;
wire n_335;
wire n_7504;
wire n_3087;
wire n_9272;
wire n_3489;
wire n_8708;
wire n_2566;
wire n_7360;
wire n_343;
wire n_7681;
wire n_308;
wire n_8448;
wire n_8076;
wire n_7301;
wire n_9041;
wire n_5129;
wire n_9643;
wire n_8904;
wire n_2149;
wire n_1078;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_8277;
wire n_3060;
wire n_4276;
wire n_7794;
wire n_7366;
wire n_8184;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_9944;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_7025;
wire n_8304;
wire n_5320;
wire n_10258;
wire n_1877;
wire n_3049;
wire n_6947;
wire n_1723;
wire n_8586;
wire n_5107;
wire n_9648;
wire n_5999;
wire n_339;
wire n_4485;
wire n_8557;
wire n_9376;
wire n_183;
wire n_8636;
wire n_7309;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_347;
wire n_6863;
wire n_9288;
wire n_6637;
wire n_798;
wire n_6100;
wire n_7860;
wire n_6735;
wire n_2659;
wire n_9521;
wire n_9541;
wire n_1414;
wire n_290;
wire n_8212;
wire n_4975;
wire n_6358;
wire n_9759;
wire n_7911;
wire n_1852;
wire n_578;
wire n_8530;
wire n_9278;
wire n_344;
wire n_9378;
wire n_8665;
wire n_5602;
wire n_9456;
wire n_9086;
wire n_3089;
wire n_7876;
wire n_6050;
wire n_422;
wire n_9711;
wire n_8933;
wire n_2470;
wire n_7244;
wire n_7960;
wire n_5405;
wire n_5253;
wire n_3985;
wire n_496;
wire n_1391;
wire n_9485;
wire n_670;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_9555;
wire n_7610;
wire n_663;
wire n_9999;
wire n_2551;
wire n_9994;
wire n_1587;
wire n_2682;
wire n_6371;
wire n_5903;
wire n_813;
wire n_8690;
wire n_8538;
wire n_1284;
wire n_7043;
wire n_3440;
wire n_6171;
wire n_7751;
wire n_8643;
wire n_6510;
wire n_1748;
wire n_4569;
wire n_6468;
wire n_9142;
wire n_2699;
wire n_9613;
wire n_4897;
wire n_888;
wire n_2769;
wire n_9440;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_8825;
wire n_2615;
wire n_3940;
wire n_7788;
wire n_446;
wire n_1064;
wire n_5842;
wire n_858;
wire n_6352;
wire n_8300;
wire n_2985;
wire n_691;
wire n_5722;
wire n_7534;
wire n_9462;
wire n_5636;
wire n_7719;
wire n_9202;
wire n_7287;
wire n_2753;
wire n_5065;
wire n_363;
wire n_1582;
wire n_7032;
wire n_8451;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_9237;
wire n_3141;
wire n_5084;
wire n_6850;
wire n_8435;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_7119;
wire n_8835;
wire n_4919;
wire n_9788;
wire n_4025;
wire n_461;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_2700;
wire n_7851;
wire n_1211;
wire n_6332;
wire n_9807;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_9573;
wire n_5877;
wire n_8963;
wire n_907;
wire n_3096;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_6434;
wire n_2356;
wire n_8713;
wire n_488;
wire n_6751;
wire n_7068;
wire n_892;
wire n_9392;
wire n_4556;
wire n_6322;
wire n_8353;
wire n_8668;
wire n_5454;
wire n_9390;
wire n_7704;
wire n_2620;
wire n_7773;
wire n_9416;
wire n_6667;
wire n_7526;
wire n_8817;
wire n_1581;
wire n_6530;
wire n_9518;
wire n_4089;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_5621;
wire n_586;
wire n_2919;
wire n_8213;
wire n_8591;
wire n_4327;
wire n_7973;
wire n_230;
wire n_953;
wire n_4218;
wire n_6429;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_7239;
wire n_2757;
wire n_10047;
wire n_963;
wire n_1052;
wire n_954;
wire n_5573;
wire n_6405;
wire n_478;
wire n_8532;
wire n_6613;
wire n_4353;
wire n_8043;
wire n_9196;
wire n_2042;
wire n_534;
wire n_7969;
wire n_6248;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_7821;
wire n_1854;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_10248;
wire n_6894;
wire n_1856;
wire n_7267;
wire n_143;
wire n_4959;
wire n_9589;
wire n_4161;
wire n_5800;
wire n_9898;
wire n_237;
wire n_832;
wire n_1319;
wire n_9373;
wire n_3992;
wire n_2616;
wire n_8606;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_6204;
wire n_2462;
wire n_1532;
wire n_7915;
wire n_3625;
wire n_8121;
wire n_1156;
wire n_8868;
wire n_794;
wire n_7387;
wire n_7431;
wire n_7654;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_686;
wire n_2837;
wire n_847;
wire n_4844;
wire n_6296;
wire n_2979;
wire n_5257;
wire n_9983;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_8276;
wire n_8718;
wire n_702;
wire n_8182;
wire n_2548;
wire n_822;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_6140;
wire n_9039;
wire n_1779;
wire n_8359;
wire n_7441;
wire n_9849;
wire n_8597;
wire n_4738;
wire n_6211;
wire n_8562;
wire n_1369;
wire n_3909;
wire n_8211;
wire n_9962;
wire n_8430;
wire n_6307;
wire n_8007;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_7394;
wire n_8600;
wire n_8311;
wire n_8943;
wire n_809;
wire n_8441;
wire n_4434;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_1942;
wire n_9829;
wire n_6860;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_8978;
wire n_411;
wire n_414;
wire n_5012;
wire n_10121;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_8198;
wire n_9988;
wire n_5697;
wire n_7188;
wire n_8526;
wire n_1810;
wire n_7573;
wire n_2813;
wire n_7879;
wire n_4438;
wire n_2009;
wire n_9848;
wire n_7087;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_7985;
wire n_9045;
wire n_9466;
wire n_6515;
wire n_9348;
wire n_8278;
wire n_6011;
wire n_7722;
wire n_7935;
wire n_8592;
wire n_6645;
wire n_8226;
wire n_3150;
wire n_747;
wire n_6984;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_10235;
wire n_10090;
wire n_615;
wire n_851;
wire n_10153;
wire n_843;
wire n_7193;
wire n_10018;
wire n_8987;
wire n_705;
wire n_3775;
wire n_4133;
wire n_6897;
wire n_7256;
wire n_678;
wire n_4184;
wire n_5203;
wire n_9071;
wire n_2518;
wire n_9356;
wire n_9464;
wire n_2629;
wire n_367;
wire n_4481;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_9239;
wire n_2181;
wire n_10053;
wire n_1829;
wire n_6183;
wire n_10051;
wire n_7522;
wire n_5882;
wire n_9606;
wire n_547;
wire n_4030;
wire n_7881;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_4397;
wire n_1710;
wire n_7502;
wire n_1128;
wire n_9492;
wire n_2928;
wire n_8960;
wire n_7335;
wire n_7103;
wire n_1734;
wire n_4820;
wire n_10151;
wire n_6246;
wire n_590;
wire n_3770;
wire n_8025;
wire n_1308;
wire n_5094;
wire n_6383;
wire n_9031;
wire n_4938;
wire n_9717;
wire n_9516;
wire n_7020;
wire n_8434;
wire n_4179;
wire n_3469;
wire n_8175;
wire n_9693;
wire n_9991;
wire n_5336;
wire n_8850;
wire n_9103;
wire n_372;
wire n_677;
wire n_9477;
wire n_2723;
wire n_314;
wire n_368;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_10253;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_8895;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_295;
wire n_133;
wire n_3113;
wire n_8046;
wire n_6904;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_568;
wire n_8867;
wire n_2856;
wire n_1832;
wire n_8239;
wire n_9599;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_7825;
wire n_8183;
wire n_8924;
wire n_9001;
wire n_3828;
wire n_10218;
wire n_3288;
wire n_5514;
wire n_5091;
wire n_7533;
wire n_4404;
wire n_8578;
wire n_9777;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_8848;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_9222;
wire n_10148;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_9366;
wire n_6611;
wire n_9449;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_906;
wire n_6116;
wire n_919;
wire n_7186;
wire n_4356;
wire n_8230;
wire n_9869;
wire n_6819;
wire n_8725;
wire n_658;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_7936;
wire n_1740;
wire n_6473;
wire n_9741;
wire n_1586;
wire n_4291;
wire n_535;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_8391;
wire n_6310;
wire n_7840;
wire n_592;
wire n_9397;
wire n_1692;
wire n_2982;
wire n_8202;
wire n_2481;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_7906;
wire n_8948;
wire n_2507;
wire n_8678;
wire n_9754;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_9179;
wire n_1614;
wire n_2339;
wire n_457;
wire n_7148;
wire n_6714;
wire n_7017;
wire n_7658;
wire n_8340;
wire n_7250;
wire n_7462;
wire n_7828;
wire n_8905;
wire n_5782;
wire n_4637;
wire n_603;
wire n_4935;
wire n_8691;
wire n_6365;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_10136;
wire n_7401;
wire n_8812;
wire n_9169;
wire n_6828;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_8704;
wire n_6355;
wire n_5596;
wire n_7887;
wire n_396;
wire n_8058;
wire n_1887;
wire n_4413;
wire n_9177;
wire n_10078;
wire n_1073;
wire n_6777;
wire n_5728;
wire n_2346;
wire n_8394;
wire n_662;
wire n_9269;
wire n_3990;
wire n_4493;
wire n_7835;
wire n_218;
wire n_3475;
wire n_1215;
wire n_8181;
wire n_9289;
wire n_8722;
wire n_1592;
wire n_6420;
wire n_6945;
wire n_2882;
wire n_9350;
wire n_1721;
wire n_7356;
wire n_2338;
wire n_7288;
wire n_7637;
wire n_5726;
wire n_7124;
wire n_3672;
wire n_7294;
wire n_5290;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_2721;
wire n_7321;
wire n_1043;
wire n_9166;
wire n_5095;
wire n_10265;
wire n_486;
wire n_8707;
wire n_3002;
wire n_6754;
wire n_337;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_8747;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_7691;
wire n_5928;
wire n_3845;
wire n_8742;
wire n_7108;
wire n_6882;
wire n_2081;
wire n_299;
wire n_7585;
wire n_9125;
wire n_7386;
wire n_4570;
wire n_8552;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7417;
wire n_7888;
wire n_2418;
wire n_9641;
wire n_9960;
wire n_7187;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_9785;
wire n_9923;
wire n_8224;
wire n_7544;
wire n_3458;
wire n_5712;
wire n_1420;
wire n_1132;
wire n_3330;
wire n_4606;
wire n_6166;
wire n_8628;
wire n_4774;
wire n_2477;
wire n_6966;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_9228;
wire n_7255;
wire n_4093;
wire n_1486;
wire n_8037;
wire n_8084;
wire n_7120;
wire n_7218;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_4174;
wire n_8289;
wire n_9801;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_309;
wire n_2367;
wire n_10249;
wire n_9645;
wire n_4766;
wire n_8045;
wire n_5633;
wire n_8697;
wire n_2896;
wire n_652;
wire n_8077;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_1927;
wire n_5583;
wire n_9457;
wire n_1349;
wire n_4460;
wire n_288;
wire n_8026;
wire n_1031;
wire n_3645;
wire n_7889;
wire n_3223;
wire n_3929;
wire n_6110;
wire n_6064;
wire n_6237;
wire n_834;
wire n_7196;
wire n_2255;
wire n_2272;
wire n_893;
wire n_9330;
wire n_6341;
wire n_10012;
wire n_1965;
wire n_9365;
wire n_1902;
wire n_6590;
wire n_1941;
wire n_5501;
wire n_8444;
wire n_9178;
wire n_8654;
wire n_10035;
wire n_9181;
wire n_7923;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_504;
wire n_6697;
wire n_874;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_7559;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_7081;
wire n_9307;
wire n_3189;
wire n_2066;
wire n_10257;
wire n_6449;
wire n_993;
wire n_7832;
wire n_7968;
wire n_3154;
wire n_1551;
wire n_545;
wire n_9238;
wire n_450;
wire n_6141;
wire n_2905;
wire n_10099;
wire n_8449;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_8493;
wire n_628;
wire n_7584;
wire n_9224;
wire n_3788;
wire n_10244;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_6983;
wire n_970;
wire n_7843;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_8958;
wire n_1534;
wire n_8443;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_9756;
wire n_7222;
wire n_3242;
wire n_9624;
wire n_495;
wire n_6071;
wire n_3525;
wire n_8161;
wire n_3486;
wire n_6808;
wire n_8734;
wire n_9547;
wire n_8271;
wire n_9594;
wire n_9901;
wire n_9895;
wire n_2405;
wire n_6724;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_9277;
wire n_4036;
wire n_6571;
wire n_921;
wire n_7470;
wire n_5100;
wire n_9189;
wire n_1795;
wire n_5849;
wire n_8495;
wire n_6251;
wire n_7400;
wire n_9548;
wire n_2578;
wire n_3483;
wire n_128;
wire n_6635;
wire n_10000;
wire n_1821;
wire n_3894;
wire n_9472;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_8994;
wire n_8901;
wire n_8056;
wire n_2656;
wire n_1080;
wire n_9538;
wire n_1274;
wire n_7623;
wire n_8954;
wire n_3524;
wire n_5616;
wire n_7597;
wire n_5034;
wire n_6733;
wire n_1708;
wire n_7071;
wire n_426;
wire n_8840;
wire n_5988;
wire n_6467;
wire n_7859;
wire n_8900;
wire n_6035;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_6522;
wire n_7109;
wire n_2092;
wire n_9434;
wire n_5959;
wire n_2075;
wire n_9052;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_1776;
wire n_4807;
wire n_6562;
wire n_6150;
wire n_9176;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_8157;
wire n_1757;
wire n_890;
wire n_8346;
wire n_1919;
wire n_9697;
wire n_960;
wire n_4230;
wire n_7882;
wire n_8827;
wire n_3419;
wire n_1290;
wire n_8309;
wire n_8344;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_1252;
wire n_9060;
wire n_348;
wire n_5754;
wire n_6016;
wire n_8096;
wire n_8100;
wire n_8822;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_9758;
wire n_3190;
wire n_7212;
wire n_1553;
wire n_3678;
wire n_7908;
wire n_2664;
wire n_8222;
wire n_3456;
wire n_9876;
wire n_5628;
wire n_444;
wire n_1808;
wire n_6726;
wire n_8406;
wire n_316;
wire n_2266;
wire n_10277;
wire n_2650;
wire n_4428;
wire n_146;
wire n_5003;
wire n_5252;
wire n_7009;
wire n_408;
wire n_6554;
wire n_10139;
wire n_10230;
wire n_967;
wire n_6689;
wire n_2731;
wire n_8866;
wire n_6143;
wire n_5614;
wire n_8693;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_10207;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_7777;
wire n_8794;
wire n_2998;
wire n_6277;
wire n_9653;
wire n_7395;
wire n_4684;
wire n_5981;
wire n_6095;
wire n_7671;
wire n_8020;
wire n_6247;
wire n_4840;
wire n_10255;
wire n_9257;
wire n_3162;
wire n_9270;
wire n_983;
wire n_2760;
wire n_6880;
wire n_3377;
wire n_3749;
wire n_10101;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_8736;
wire n_6499;
wire n_6837;
wire n_4423;
wire n_10063;
wire n_4096;
wire n_7393;
wire n_2881;
wire n_8400;
wire n_6616;
wire n_1203;
wire n_9686;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_7871;
wire n_321;
wire n_6946;
wire n_4996;
wire n_621;
wire n_2475;
wire n_8055;
wire n_8333;
wire n_10195;
wire n_9718;
wire n_4598;
wire n_5064;
wire n_9215;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_507;
wire n_8909;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_7484;
wire n_5173;
wire n_6305;
wire n_1228;
wire n_6317;
wire n_3920;
wire n_9762;
wire n_9407;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_828;
wire n_779;
wire n_9964;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_7649;
wire n_1439;
wire n_9953;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_9153;
wire n_945;
wire n_6693;
wire n_8786;
wire n_8541;
wire n_3743;
wire n_6734;
wire n_10173;
wire n_9571;
wire n_7135;
wire n_7014;
wire n_8263;
wire n_1932;
wire n_8884;
wire n_5597;
wire n_4721;
wire n_5635;
wire n_984;
wire n_694;
wire n_6382;
wire n_9019;
wire n_7328;
wire n_1983;
wire n_7635;
wire n_6404;
wire n_10229;
wire n_5975;
wire n_9737;
wire n_4029;
wire n_1594;
wire n_8494;
wire n_900;
wire n_3870;
wire n_6379;
wire n_7703;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_9468;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_6235;
wire n_9870;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_9026;
wire n_3094;
wire n_9710;
wire n_2310;
wire n_3952;
wire n_7265;
wire n_8638;
wire n_2287;
wire n_2860;
wire n_8710;
wire n_2056;
wire n_10019;
wire n_6789;
wire n_7184;
wire n_6440;
wire n_9725;
wire n_6417;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_8177;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_9084;
wire n_7728;
wire n_3442;
wire n_1201;
wire n_7690;
wire n_1114;
wire n_7219;
wire n_7479;
wire n_3998;
wire n_9419;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_669;
wire n_7270;
wire n_1176;
wire n_8170;
wire n_5940;
wire n_8893;
wire n_1149;
wire n_7390;
wire n_1020;
wire n_7805;
wire n_7807;
wire n_211;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_8589;
wire n_9479;
wire n_9820;
wire n_4667;
wire n_2325;
wire n_178;
wire n_8320;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_6272;
wire n_8153;
wire n_7699;
wire n_6484;
wire n_661;
wire n_7674;
wire n_6236;
wire n_8620;
wire n_5576;
wire n_4668;
wire n_8298;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_849;
wire n_6871;
wire n_10270;
wire n_584;
wire n_8235;
wire n_1786;
wire n_430;
wire n_5284;
wire n_9294;
wire n_9126;
wire n_8370;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_6768;
wire n_4759;
wire n_7951;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_7506;
wire n_2340;
wire n_3552;
wire n_875;
wire n_357;
wire n_6717;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_165;
wire n_5578;
wire n_2361;
wire n_8395;
wire n_1173;
wire n_1603;
wire n_969;
wire n_1401;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_8906;
wire n_5530;
wire n_8097;
wire n_304;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_8570;
wire n_5741;
wire n_8902;
wire n_5991;
wire n_3933;
wire n_7330;
wire n_3206;
wire n_7928;
wire n_5506;
wire n_5243;
wire n_3966;
wire n_9819;
wire n_8477;
wire n_5449;
wire n_10236;
wire n_1702;
wire n_6992;
wire n_5221;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_6000;
wire n_9545;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_2649;
wire n_6655;
wire n_7892;
wire n_9165;
wire n_7304;
wire n_10143;
wire n_5792;
wire n_1187;
wire n_6657;
wire n_7756;
wire n_8129;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_8580;
wire n_2542;
wire n_2313;
wire n_7990;
wire n_489;
wire n_1174;
wire n_3914;
wire n_3324;
wire n_4625;
wire n_8122;
wire n_2558;
wire n_8259;
wire n_2063;
wire n_3803;
wire n_8536;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_2252;
wire n_8748;
wire n_7612;
wire n_6113;
wire n_7789;
wire n_4819;
wire n_9056;
wire n_1685;
wire n_917;
wire n_1714;
wire n_8094;
wire n_9341;
wire n_6242;
wire n_7902;
wire n_7088;
wire n_6519;
wire n_8572;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_8120;
wire n_6842;
wire n_7588;
wire n_3390;
wire n_1573;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_2373;
wire n_9172;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_210;
wire n_1737;
wire n_9145;
wire n_6801;
wire n_8099;
wire n_9996;
wire n_10059;
wire n_774;
wire n_2493;
wire n_4930;
wire n_7680;
wire n_8770;
wire n_5276;
wire n_6308;
wire n_1059;
wire n_7398;
wire n_1133;
wire n_6906;
wire n_5078;
wire n_4537;
wire n_7230;
wire n_8700;
wire n_2885;
wire n_9906;
wire n_6629;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_6968;
wire n_9920;
wire n_4282;
wire n_9504;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_665;
wire n_3839;
wire n_1440;
wire n_9482;
wire n_5205;
wire n_9138;
wire n_3333;
wire n_9384;
wire n_8637;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_8757;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_2602;
wire n_5819;
wire n_10147;
wire n_205;
wire n_4579;
wire n_4616;
wire n_8903;
wire n_1496;
wire n_9193;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_6398;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_232;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_9527;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_427;
wire n_3368;
wire n_8585;
wire n_9064;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_8982;
wire n_2765;
wire n_3329;
wire n_6415;
wire n_2994;
wire n_10032;
wire n_6857;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_10200;
wire n_7842;
wire n_2003;
wire n_5856;
wire n_1457;
wire n_8709;
wire n_5446;
wire n_9383;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_9735;
wire n_9943;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_6413;
wire n_7679;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_6361;
wire n_9357;
wire n_3438;
wire n_6231;
wire n_7783;
wire n_4098;
wire n_872;
wire n_594;
wire n_200;
wire n_5684;
wire n_5861;
wire n_8108;
wire n_1297;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_7862;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_5312;
wire n_985;
wire n_5850;
wire n_10014;
wire n_3404;
wire n_3425;
wire n_3217;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_9986;
wire n_626;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_7820;
wire n_7167;
wire n_8692;
wire n_7833;
wire n_2023;
wire n_8820;
wire n_3249;
wire n_2351;
wire n_7643;
wire n_8490;
wire n_676;
wire n_5113;
wire n_4442;
wire n_9491;
wire n_4698;
wire n_642;
wire n_9922;
wire n_6712;
wire n_1602;
wire n_194;
wire n_1178;
wire n_5687;
wire n_4779;
wire n_8062;
wire n_8781;
wire n_2286;
wire n_10203;
wire n_4966;
wire n_503;
wire n_8000;
wire n_2065;
wire n_10061;
wire n_4017;
wire n_8808;
wire n_8233;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_9747;
wire n_620;
wire n_6953;
wire n_1081;
wire n_4418;
wire n_8685;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_9061;
wire n_9168;
wire n_1318;
wire n_780;
wire n_8575;
wire n_8701;
wire n_2977;
wire n_6303;
wire n_6474;
wire n_6182;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_5674;
wire n_3600;
wire n_8670;
wire n_245;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_1388;
wire n_8352;
wire n_7993;
wire n_7930;
wire n_2836;
wire n_5682;
wire n_672;
wire n_8385;
wire n_8875;
wire n_6392;
wire n_8166;
wire n_581;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_8934;
wire n_5117;
wire n_2773;
wire n_9073;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_7999;
wire n_5612;
wire n_265;
wire n_6125;
wire n_443;
wire n_6599;
wire n_7963;
wire n_6685;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_8389;
wire n_9068;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_10158;
wire n_6560;
wire n_1326;
wire n_3176;
wire n_8659;
wire n_8804;
wire n_10043;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_8439;
wire n_9544;
wire n_8814;
wire n_8369;
wire n_5301;
wire n_7800;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_7615;
wire n_9286;
wire n_5898;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_7298;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_7581;
wire n_10131;
wire n_4049;
wire n_6641;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_5563;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_6673;
wire n_8789;
wire n_7172;
wire n_7074;
wire n_5497;
wire n_8790;
wire n_8234;
wire n_4724;
wire n_5832;
wire n_1238;
wire n_7190;
wire n_7112;
wire n_7678;
wire n_10082;
wire n_9265;
wire n_1772;
wire n_282;
wire n_752;
wire n_1476;
wire n_9080;
wire n_1108;
wire n_5526;
wire n_8989;
wire n_10152;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_6195;
wire n_862;
wire n_3584;
wire n_6356;
wire n_8927;
wire n_3756;
wire n_9770;
wire n_381;
wire n_2889;
wire n_9463;
wire n_7001;
wire n_390;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_2772;
wire n_7369;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_7829;
wire n_4382;
wire n_1554;
wire n_9939;
wire n_10159;
wire n_3999;
wire n_8534;
wire n_2844;
wire n_9911;
wire n_9210;
wire n_2138;
wire n_5211;
wire n_6559;
wire n_5230;
wire n_10122;
wire n_7359;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_7144;
wire n_4833;
wire n_8756;
wire n_6841;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_9691;
wire n_5110;
wire n_6653;
wire n_379;
wire n_428;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_8832;
wire n_1973;
wire n_5737;
wire n_786;
wire n_1142;
wire n_9340;
wire n_9351;
wire n_8461;
wire n_8042;
wire n_2579;
wire n_6825;
wire n_6923;
wire n_9950;
wire n_1770;
wire n_138;
wire n_4228;
wire n_4401;
wire n_8021;
wire n_1756;
wire n_8839;
wire n_1716;
wire n_6112;
wire n_2788;
wire n_6547;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_9155;
wire n_6399;
wire n_8623;
wire n_1873;
wire n_3201;
wire n_8758;
wire n_221;
wire n_622;
wire n_6275;
wire n_1087;
wire n_6575;
wire n_5666;
wire n_3472;
wire n_7924;
wire n_7732;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_8511;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_8595;
wire n_1272;
wire n_8873;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7459;
wire n_1247;
wire n_7191;
wire n_9201;
wire n_9823;
wire n_9688;
wire n_7096;
wire n_591;
wire n_3050;
wire n_313;
wire n_8455;
wire n_1478;
wire n_8280;
wire n_3903;
wire n_10102;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_9595;
wire n_5272;
wire n_9530;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_6826;
wire n_9227;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_8372;
wire n_5361;
wire n_8598;
wire n_5683;
wire n_369;
wire n_4171;
wire n_5847;
wire n_7551;
wire n_9400;
wire n_4045;
wire n_598;
wire n_6678;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_9025;
wire n_1460;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_8282;
wire n_7750;
wire n_517;
wire n_413;
wire n_5015;
wire n_2702;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_6748;
wire n_2030;
wire n_903;
wire n_8616;
wire n_3115;
wire n_4749;
wire n_203;
wire n_8336;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_6752;
wire n_9749;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_9285;
wire n_9972;
wire n_10058;
wire n_2209;
wire n_7652;
wire n_8847;
wire n_7808;
wire n_6500;
wire n_4270;
wire n_8135;
wire n_9214;
wire n_2797;
wire n_1255;
wire n_7051;
wire n_9859;
wire n_5152;
wire n_9003;
wire n_2321;
wire n_9271;
wire n_722;
wire n_9258;
wire n_3680;
wire n_6628;
wire n_844;
wire n_201;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_6975;
wire n_1601;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_7536;
wire n_8979;
wire n_8529;
wire n_5688;
wire n_9763;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_9597;
wire n_979;
wire n_2841;
wire n_6293;
wire n_8417;
wire n_9965;
wire n_9076;
wire n_7952;
wire n_3322;
wire n_4576;
wire n_9393;
wire n_8498;
wire n_846;
wire n_2427;
wire n_2505;
wire n_7991;
wire n_7676;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_585;
wire n_7553;
wire n_6905;
wire n_7425;
wire n_270;
wire n_2594;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_8967;
wire n_8355;
wire n_9736;
wire n_4767;
wire n_7998;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_8719;
wire n_3112;
wire n_2349;
wire n_6581;
wire n_10160;
wire n_1379;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_5415;
wire n_4676;
wire n_10241;
wire n_5770;
wire n_7064;
wire n_5892;
wire n_8762;
wire n_4544;
wire n_10180;
wire n_2170;
wire n_8516;
wire n_8880;
wire n_1091;
wire n_6577;
wire n_6899;
wire n_8784;
wire n_641;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_8237;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_9803;
wire n_4429;
wire n_8977;
wire n_575;
wire n_8171;
wire n_4591;
wire n_6370;
wire n_9755;
wire n_3266;
wire n_9805;
wire n_7210;
wire n_4646;
wire n_7899;
wire n_9728;
wire n_5769;
wire n_6065;
wire n_1130;
wire n_7039;
wire n_9659;
wire n_6987;
wire n_4563;
wire n_4725;
wire n_9107;
wire n_2210;
wire n_4169;
wire n_6190;
wire n_6859;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_9917;
wire n_3066;
wire n_6309;
wire n_9520;
wire n_246;
wire n_6623;
wire n_7723;
wire n_2426;
wire n_6527;
wire n_7443;
wire n_9583;
wire n_7811;
wire n_657;
wire n_4320;
wire n_5341;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_9036;
wire n_491;
wire n_9522;
wire n_5979;
wire n_160;
wire n_566;
wire n_565;
wire n_5271;
wire n_5089;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1505;
wire n_1181;
wire n_6929;
wire n_4012;
wire n_5518;
wire n_10125;
wire n_651;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_8279;
wire n_5622;
wire n_807;
wire n_3910;
wire n_4711;
wire n_9723;
wire n_835;
wire n_3319;
wire n_7348;
wire n_10254;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_8912;
wire n_2689;
wire n_3259;
wire n_9488;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_7155;
wire n_8227;
wire n_3688;
wire n_9231;
wire n_8938;
wire n_6865;
wire n_3016;
wire n_1693;
wire n_8787;
wire n_5393;
wire n_10017;
wire n_2599;
wire n_6535;
wire n_904;
wire n_3338;
wire n_7213;
wire n_3414;
wire n_9047;
wire n_1827;
wire n_4671;
wire n_8270;
wire n_4209;
wire n_1271;
wire n_5966;
wire n_1542;
wire n_7456;
wire n_8335;
wire n_5041;
wire n_7420;
wire n_9798;
wire n_9681;
wire n_8054;
wire n_1423;
wire n_9414;
wire n_1166;
wire n_8607;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_9979;
wire n_785;
wire n_9093;
wire n_2200;
wire n_3261;
wire n_6482;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_8150;
wire n_5059;
wire n_9379;
wire n_5505;
wire n_3127;
wire n_7715;
wire n_9486;
wire n_226;
wire n_1780;
wire n_3732;
wire n_6605;
wire n_9134;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_7007;
wire n_8358;
wire n_4699;
wire n_9410;
wire n_3906;
wire n_4127;
wire n_880;
wire n_10045;
wire n_3297;
wire n_544;
wire n_155;
wire n_7909;
wire n_2683;
wire n_1370;
wire n_9151;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_8281;
wire n_9182;
wire n_5908;
wire n_6018;
wire n_4202;
wire n_7168;
wire n_5212;
wire n_9976;
wire n_7736;
wire n_5000;
wire n_8396;
wire n_9591;
wire n_2853;
wire n_1323;
wire n_9838;
wire n_688;
wire n_7177;
wire n_5939;
wire n_10033;
wire n_3766;
wire n_1353;
wire n_800;
wire n_9568;
wire n_7780;
wire n_2880;
wire n_9261;
wire n_9701;
wire n_7379;
wire n_1666;
wire n_4165;
wire n_2389;
wire n_3350;
wire n_4866;
wire n_7444;
wire n_8223;
wire n_5931;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_7813;
wire n_864;
wire n_7030;
wire n_8459;
wire n_5420;
wire n_1264;
wire n_6311;
wire n_447;
wire n_4412;
wire n_3599;
wire n_3407;
wire n_6654;
wire n_6424;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_9752;
wire n_1580;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_497;
wire n_1607;
wire n_8379;
wire n_6879;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_5679;
wire n_947;
wire n_373;
wire n_3710;
wire n_5938;
wire n_9079;
wire n_307;
wire n_6702;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_5098;
wire n_1230;
wire n_4144;
wire n_5724;
wire n_10064;
wire n_5774;
wire n_375;
wire n_2165;
wire n_8793;
wire n_6452;
wire n_929;
wire n_3379;
wire n_4374;
wire n_8975;
wire n_6791;
wire n_3532;
wire n_9170;
wire n_8792;
wire n_1124;
wire n_5131;
wire n_7280;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_8489;
wire n_7110;
wire n_6915;
wire n_8671;
wire n_1104;
wire n_1294;
wire n_7511;
wire n_1257;
wire n_6856;
wire n_1182;
wire n_7941;
wire n_7791;
wire n_9385;
wire n_3531;
wire n_8484;
wire n_2963;
wire n_3834;
wire n_8454;
wire n_10238;
wire n_7232;
wire n_8759;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_8703;
wire n_5790;
wire n_3258;
wire n_10206;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_9670;
wire n_2047;
wire n_6364;
wire n_6451;
wire n_6552;
wire n_1845;
wire n_240;
wire n_2193;
wire n_8325;
wire n_2478;
wire n_5140;
wire n_6328;
wire n_9598;
wire n_4816;
wire n_231;
wire n_8382;
wire n_7827;
wire n_8971;
wire n_1483;
wire n_6363;
wire n_2983;
wire n_7159;
wire n_8127;
wire n_227;
wire n_10079;
wire n_10188;
wire n_3810;
wire n_1289;
wire n_8721;
wire n_9391;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_8889;
wire n_6406;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_9470;
wire n_370;
wire n_5306;
wire n_6978;
wire n_9328;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_9245;
wire n_8232;
wire n_2651;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_7363;
wire n_9833;
wire n_10213;
wire n_6612;
wire n_10107;
wire n_8664;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_9455;
wire n_955;
wire n_5511;
wire n_7863;
wire n_5680;
wire n_9719;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_7295;
wire n_8633;
wire n_9744;
wire n_8842;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_550;
wire n_897;
wire n_8956;
wire n_5280;
wire n_6375;
wire n_6479;
wire n_1428;
wire n_6866;
wire n_7831;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_9698;
wire n_6170;
wire n_1931;
wire n_9124;
wire n_9695;
wire n_4187;
wire n_1070;
wire n_6447;
wire n_4166;
wire n_6263;
wire n_7093;
wire n_9497;
wire n_5206;
wire n_1030;
wire n_8641;
wire n_8479;
wire n_3222;
wire n_1071;
wire n_7466;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_6130;
wire n_1513;
wire n_2970;
wire n_7651;
wire n_2235;
wire n_673;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_680;
wire n_3755;
wire n_8179;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_8973;
wire n_6935;
wire n_1590;
wire n_10194;
wire n_9775;
wire n_7530;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_675;
wire n_4064;
wire n_9038;
wire n_8308;
wire n_4936;
wire n_9630;
wire n_5387;
wire n_1556;
wire n_184;
wire n_1863;
wire n_8378;
wire n_3841;
wire n_8733;
wire n_2118;
wire n_8809;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_468;
wire n_9652;
wire n_10021;
wire n_5058;
wire n_6907;
wire n_129;
wire n_8500;
wire n_6158;
wire n_7661;
wire n_9709;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_8447;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_1322;
wire n_9324;
wire n_3690;
wire n_9934;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_8548;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_8412;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_477;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_9668;
wire n_1971;
wire n_3252;
wire n_7145;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_9877;
wire n_4310;
wire n_9657;
wire n_10111;
wire n_6338;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_9352;
wire n_3954;
wire n_9395;
wire n_8425;
wire n_9349;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_8241;
wire n_7823;
wire n_9209;
wire n_7467;
wire n_736;
wire n_5097;
wire n_10113;
wire n_7932;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_9969;
wire n_3071;
wire n_3739;
wire n_9937;
wire n_593;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_7541;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_7241;
wire n_7717;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_9618;
wire n_10009;
wire n_289;
wire n_4850;
wire n_6625;
wire n_3781;
wire n_4912;
wire n_4813;
wire n_7464;
wire n_9082;
wire n_2590;
wire n_6302;
wire n_9424;
wire n_8274;
wire n_9453;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_8152;
wire n_9637;
wire n_3328;
wire n_6706;
wire n_944;
wire n_8550;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_8264;
wire n_7434;
wire n_7636;
wire n_7054;
wire n_6999;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_8829;
wire n_9183;
wire n_9205;
wire n_9009;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_6228;
wire n_857;
wire n_5650;
wire n_2636;
wire n_10044;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_10221;
wire n_4702;
wire n_6888;
wire n_8266;
wire n_8515;
wire n_10109;
wire n_10169;
wire n_4252;
wire n_4457;
wire n_8648;
wire n_6063;
wire n_971;
wire n_9030;
wire n_9024;
wire n_9523;
wire n_9377;
wire n_8946;
wire n_404;
wire n_6800;
wire n_5139;
wire n_9716;
wire n_1393;
wire n_2319;
wire n_6922;
wire n_596;
wire n_9380;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_8744;
wire n_9000;
wire n_9679;
wire n_9116;
wire n_9742;
wire n_9016;
wire n_7503;
wire n_2808;
wire n_6070;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_9006;
wire n_10091;
wire n_6651;
wire n_7296;
wire n_7091;
wire n_4491;
wire n_7273;
wire n_6647;
wire n_5821;
wire n_266;
wire n_2930;
wire n_5733;
wire n_10029;
wire n_1838;
wire n_9690;
wire n_3514;
wire n_2777;
wire n_8765;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_9852;
wire n_7543;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_9914;
wire n_6184;
wire n_4886;
wire n_8627;
wire n_4090;
wire n_2529;
wire n_7507;
wire n_9451;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_9760;
wire n_1481;
wire n_7555;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_10272;
wire n_868;
wire n_9035;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_9211;
wire n_914;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_9677;
wire n_5048;
wire n_5521;
wire n_7578;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_759;
wire n_8195;
wire n_9070;
wire n_5585;
wire n_6397;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_7033;
wire n_9881;
wire n_324;
wire n_6121;
wire n_1571;
wire n_3119;
wire n_9669;
wire n_7531;
wire n_4142;
wire n_9958;
wire n_1189;
wire n_4082;
wire n_9858;
wire n_8462;
wire n_5561;
wire n_3479;
wire n_9981;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_8377;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_9588;
wire n_6954;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_523;
wire n_1537;
wire n_5875;
wire n_8428;
wire n_8103;
wire n_4262;
wire n_9021;
wire n_2671;
wire n_6646;
wire n_8936;
wire n_8414;
wire n_8362;
wire n_9682;
wire n_1798;
wire n_10137;
wire n_1790;
wire n_4720;
wire n_7131;
wire n_7769;
wire n_6903;
wire n_9050;
wire n_9303;
wire n_9495;
wire n_525;
wire n_1647;
wire n_4685;
wire n_6101;
wire n_9415;
wire n_5968;
wire n_2563;
wire n_10196;
wire n_2387;
wire n_8491;
wire n_9058;
wire n_4334;
wire n_1674;
wire n_6941;
wire n_9845;
wire n_1830;
wire n_2073;
wire n_8831;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_8324;
wire n_139;
wire n_5515;
wire n_6106;
wire n_9822;
wire n_6604;
wire n_4014;
wire n_7418;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_7688;
wire n_2913;
wire n_2336;
wire n_254;
wire n_9640;
wire n_1233;
wire n_8348;
wire n_5607;
wire n_1615;
wire n_4175;
wire n_8288;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_244;
wire n_4648;
wire n_1333;
wire n_8269;
wire n_5006;
wire n_7806;
wire n_10085;
wire n_6566;
wire n_8625;
wire n_1443;
wire n_946;
wire n_1539;
wire n_5734;
wire n_6081;
wire n_8458;
wire n_4892;
wire n_8806;
wire n_7204;
wire n_3823;
wire n_8180;
wire n_1866;
wire n_4173;
wire n_689;
wire n_8601;
wire n_738;
wire n_1624;
wire n_4970;
wire n_8499;
wire n_640;
wire n_9062;
wire n_3816;
wire n_1279;
wire n_8306;
wire n_4108;
wire n_4486;
wire n_610;
wire n_5404;
wire n_9722;
wire n_6047;
wire n_2960;
wire n_8167;
wire n_1090;
wire n_5438;
wire n_9791;
wire n_633;
wire n_9229;
wire n_439;
wire n_4627;
wire n_8613;
wire n_9603;
wire n_758;
wire n_8913;
wire n_7448;
wire n_7354;
wire n_8800;
wire n_6244;
wire n_2290;
wire n_8768;
wire n_6861;
wire n_9099;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_9309;
wire n_7852;
wire n_1049;
wire n_2145;
wire n_5725;
wire n_1639;
wire n_7925;
wire n_1068;
wire n_3030;
wire n_9432;
wire n_2580;
wire n_9454;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_9065;
wire n_331;
wire n_5163;
wire n_2039;
wire n_7748;
wire n_5768;
wire n_4961;
wire n_7556;
wire n_3753;
wire n_7640;
wire n_8187;
wire n_8881;
wire n_2035;
wire n_9704;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_7422;
wire n_7920;
wire n_8433;
wire n_9837;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_9431;
wire n_10167;
wire n_3969;
wire n_9160;
wire n_2459;
wire n_4154;
wire n_9433;
wire n_6588;
wire n_152;
wire n_3396;
wire n_9256;
wire n_9706;
wire n_1445;
wire n_7900;
wire n_7050;
wire n_4023;
wire n_9808;
wire n_9915;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_7136;
wire n_8316;
wire n_7318;
wire n_6055;
wire n_5138;
wire n_1017;
wire n_8397;
wire n_9184;
wire n_5374;
wire n_9133;
wire n_6108;
wire n_8115;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_6165;
wire n_1828;
wire n_6621;
wire n_2320;
wire n_1045;
wire n_7175;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_7810;
wire n_9109;
wire n_4640;
wire n_2583;
wire n_484;
wire n_6323;
wire n_1033;
wire n_8523;
wire n_9207;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_636;
wire n_4367;
wire n_6480;
wire n_2087;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_6597;
wire n_1009;
wire n_454;
wire n_9673;
wire n_8891;
wire n_1989;
wire n_3818;
wire n_7817;
wire n_8294;
wire n_2523;
wire n_255;
wire n_6933;
wire n_4387;
wire n_7878;
wire n_8338;
wire n_4951;
wire n_9010;
wire n_8915;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_1578;
wire n_7289;
wire n_5805;
wire n_7665;
wire n_8131;
wire n_9552;
wire n_3719;
wire n_7855;
wire n_1959;
wire n_3681;
wire n_9841;
wire n_2737;
wire n_1574;
wire n_9230;
wire n_2399;
wire n_7764;
wire n_4308;
wire n_2812;
wire n_473;
wire n_2355;
wire n_2133;
wire n_10198;
wire n_8027;
wire n_6216;
wire n_10096;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_8162;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_2725;
wire n_9132;
wire n_614;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_8855;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_8546;
wire n_9878;
wire n_773;
wire n_208;
wire n_9069;
wire n_8966;
wire n_142;
wire n_7263;
wire n_8487;
wire n_743;
wire n_8844;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_296;
wire n_6911;
wire n_3268;
wire n_9674;
wire n_8533;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_8869;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_9786;
wire n_1237;
wire n_6327;
wire n_8584;
wire n_8932;
wire n_2595;
wire n_9063;
wire n_8998;
wire n_761;
wire n_6607;
wire n_9188;
wire n_9467;
wire n_9372;
wire n_3411;
wire n_4958;
wire n_329;
wire n_9743;
wire n_4271;
wire n_7850;
wire n_7509;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_8480;
wire n_9926;
wire n_7240;
wire n_10094;
wire n_4071;
wire n_4921;
wire n_130;
wire n_1980;
wire n_8911;
wire n_5427;
wire n_5639;
wire n_7725;
wire n_8398;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_8772;
wire n_263;
wire n_4614;
wire n_9480;
wire n_1265;
wire n_8307;
wire n_224;
wire n_8767;
wire n_9113;
wire n_2681;
wire n_9158;
wire n_3103;
wire n_4945;
wire n_765;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_8010;
wire n_1015;
wire n_7278;
wire n_1651;
wire n_9263;
wire n_8347;
wire n_7630;
wire n_2775;
wire n_10162;
wire n_8466;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_9632;
wire n_511;
wire n_8813;
wire n_358;
wire n_1101;
wire n_8354;
wire n_1106;
wire n_4326;
wire n_6695;
wire n_3557;
wire n_8204;
wire n_2230;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_7565;
wire n_9282;
wire n_2851;
wire n_4305;
wire n_174;
wire n_5781;
wire n_7883;
wire n_1455;
wire n_6600;
wire n_767;
wire n_2490;
wire n_1407;
wire n_7410;
wire n_441;
wire n_4213;
wire n_2849;
wire n_7097;
wire n_3692;
wire n_2204;
wire n_9503;
wire n_6421;
wire n_5747;
wire n_7414;
wire n_7495;
wire n_9782;
wire n_5969;
wire n_9114;
wire n_365;
wire n_8312;
wire n_9855;
wire n_4929;
wire n_8040;
wire n_729;
wire n_9347;
wire n_1961;
wire n_4964;
wire n_911;
wire n_9469;
wire n_9680;
wire n_9746;
wire n_1430;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_9633;
wire n_513;
wire n_6458;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_6746;
wire n_8132;
wire n_2508;
wire n_4031;
wire n_7586;
wire n_9501;
wire n_7720;
wire n_6719;
wire n_2416;
wire n_5437;
wire n_623;
wire n_9148;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_2461;
wire n_490;
wire n_6506;
wire n_2243;
wire n_4583;
wire n_6287;
wire n_233;
wire n_6662;
wire n_572;
wire n_8650;
wire n_9585;
wire n_10267;
wire n_8974;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_8688;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_8983;
wire n_2368;
wire n_6851;
wire n_8116;
wire n_9338;
wire n_6687;
wire n_2890;
wire n_6884;
wire n_2554;
wire n_8356;
wire n_8013;
wire n_9075;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_6780;
wire n_6513;
wire n_4891;
wire n_8519;
wire n_7841;
wire n_6619;
wire n_8193;
wire n_391;
wire n_701;
wire n_1023;
wire n_5603;
wire n_539;
wire n_6804;
wire n_803;
wire n_1092;
wire n_3559;
wire n_9370;
wire n_2661;
wire n_2572;
wire n_9409;
wire n_5716;
wire n_3993;
wire n_10138;
wire n_4940;
wire n_6516;
wire n_5208;
wire n_7490;
wire n_1056;
wire n_3588;
wire n_7792;
wire n_6924;
wire n_2308;
wire n_4590;
wire n_7492;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_8329;
wire n_5237;
wire n_7809;
wire n_4664;
wire n_9626;
wire n_3860;
wire n_8154;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_7073;
wire n_2191;
wire n_10007;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_9961;
wire n_1346;
wire n_5727;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_9098;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_1060;
wire n_5347;
wire n_9861;
wire n_3298;
wire n_3033;
wire n_2824;
wire n_248;
wire n_6788;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_6393;
wire n_9536;
wire n_2333;
wire n_8566;
wire n_8086;
wire n_2916;
wire n_8746;
wire n_6249;
wire n_483;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_9593;
wire n_2403;
wire n_9017;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_9703;
wire n_2792;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_378;
wire n_1112;
wire n_3134;
wire n_6572;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_4536;
wire n_7569;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_5967;
wire n_7003;
wire n_9565;
wire n_7897;
wire n_4773;
wire n_7962;
wire n_8942;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_2472;
wire n_4611;
wire n_8113;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_455;
wire n_2993;
wire n_1719;
wire n_8652;
wire n_3864;
wire n_385;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_7419;
wire n_5827;
wire n_1560;
wire n_9337;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_7784;
wire n_1953;
wire n_4422;
wire n_8714;
wire n_6123;
wire n_6934;
wire n_2589;
wire n_7094;
wire n_7500;
wire n_1363;
wire n_1301;
wire n_3482;
wire n_6082;
wire n_8944;
wire n_2233;
wire n_9232;
wire n_1312;
wire n_804;
wire n_9320;
wire n_537;
wire n_4555;
wire n_2827;
wire n_9167;
wire n_5136;
wire n_7864;
wire n_5228;
wire n_153;
wire n_1504;
wire n_10034;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_7790;
wire n_3572;
wire n_250;
wire n_992;
wire n_4215;
wire n_6952;
wire n_7062;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_9526;
wire n_260;
wire n_8107;
wire n_842;
wire n_5471;
wire n_7642;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_9077;
wire n_7045;
wire n_1643;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_9692;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_9141;
wire n_5338;
wire n_7238;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_7126;
wire n_9745;
wire n_5669;
wire n_9787;
wire n_3854;
wire n_8674;
wire n_2468;
wire n_7931;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_540;
wire n_8482;
wire n_8992;
wire n_323;
wire n_6979;
wire n_10024;
wire n_9892;
wire n_6203;
wire n_7405;
wire n_7739;
wire n_894;
wire n_3253;
wire n_8761;
wire n_7207;
wire n_9078;
wire n_8899;
wire n_4027;
wire n_7934;
wire n_831;
wire n_2280;
wire n_9015;
wire n_7454;
wire n_9012;
wire n_4599;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_9233;
wire n_9217;
wire n_1511;
wire n_6368;
wire n_5760;
wire n_234;
wire n_3689;
wire n_6556;
wire n_2020;
wire n_4628;
wire n_9435;
wire n_5668;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_8926;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_9389;
wire n_4458;
wire n_6596;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_6870;
wire n_7639;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_10129;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_635;
wire n_10084;
wire n_7251;
wire n_2303;
wire n_7776;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_7059;
wire n_8561;
wire n_8255;
wire n_7035;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_8029;
wire n_4573;
wire n_6713;
wire n_4118;
wire n_5289;
wire n_5513;
wire n_6747;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_9381;
wire n_4079;
wire n_4091;
wire n_681;
wire n_1638;
wire n_9873;
wire n_5916;
wire n_7029;
wire n_5984;
wire n_7317;
wire n_2002;
wire n_5145;
wire n_9575;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_5132;
wire n_830;
wire n_5191;
wire n_6333;
wire n_6262;
wire n_3085;
wire n_5869;
wire n_8130;
wire n_5925;
wire n_1655;
wire n_9023;
wire n_749;
wire n_6240;
wire n_5359;
wire n_6412;
wire n_9412;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_7782;
wire n_7220;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_482;
wire n_7438;
wire n_1232;
wire n_734;
wire n_9955;
wire n_10161;
wire n_2638;
wire n_7515;
wire n_7574;
wire n_4044;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_8921;
wire n_3971;
wire n_7065;
wire n_10271;
wire n_1338;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_7894;
wire n_1522;
wire n_7868;
wire n_9418;
wire n_6973;
wire n_2949;
wire n_9733;
wire n_2711;
wire n_5363;
wire n_7285;
wire n_8286;
wire n_5200;
wire n_9502;
wire n_338;
wire n_1653;
wire n_5659;
wire n_1506;
wire n_5618;
wire n_6325;
wire n_990;
wire n_2867;
wire n_9765;
wire n_1894;
wire n_975;
wire n_9029;
wire n_2794;
wire n_567;
wire n_3145;
wire n_10163;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_151;
wire n_6721;
wire n_8178;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_9623;
wire n_2392;
wire n_7008;
wire n_711;
wire n_8925;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_8432;
wire n_6111;
wire n_1834;
wire n_10130;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_8047;
wire n_617;
wire n_6260;
wire n_7501;
wire n_1572;
wire n_1968;
wire n_10214;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_6665;
wire n_9783;
wire n_7566;
wire n_7937;
wire n_7055;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_8268;
wire n_8053;
wire n_5858;
wire n_5817;
wire n_6690;
wire n_9840;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_217;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_726;
wire n_9909;
wire n_10192;
wire n_7113;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_8735;
wire n_818;
wire n_7872;
wire n_1970;
wire n_10219;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_8845;
wire n_7242;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_8830;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_7954;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_7819;
wire n_6570;
wire n_1410;
wire n_707;
wire n_8022;
wire n_9532;
wire n_8415;
wire n_9112;
wire n_6498;
wire n_3902;
wire n_10062;
wire n_4730;
wire n_7228;
wire n_9561;
wire n_6692;
wire n_8547;
wire n_937;
wire n_6074;
wire n_2779;
wire n_7561;
wire n_1584;
wire n_487;
wire n_6380;
wire n_3654;
wire n_2164;
wire n_10216;
wire n_9091;
wire n_5996;
wire n_8386;
wire n_8426;
wire n_2115;
wire n_9326;
wire n_8672;
wire n_10049;
wire n_2232;
wire n_5327;
wire n_7994;
wire n_9180;
wire n_8540;
wire n_6045;
wire n_9932;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_9220;
wire n_9834;
wire n_2811;
wire n_3348;
wire n_179;
wire n_7415;
wire n_410;
wire n_9474;
wire n_7793;
wire n_5796;
wire n_7702;
wire n_9542;
wire n_7598;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_895;
wire n_3358;
wire n_8192;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_8791;
wire n_9458;
wire n_4204;
wire n_9642;
wire n_6877;
wire n_6772;
wire n_1543;
wire n_2224;
wire n_1991;
wire n_6823;
wire n_9020;
wire n_732;
wire n_6806;
wire n_7426;
wire n_9910;
wire n_5906;
wire n_8350;
wire n_9100;
wire n_4743;
wire n_500;
wire n_8816;
wire n_1067;
wire n_3805;
wire n_7957;
wire n_3825;
wire n_8712;
wire n_8048;
wire n_6831;
wire n_148;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_9781;
wire n_8663;
wire n_4859;
wire n_7217;
wire n_9940;
wire n_2692;
wire n_538;
wire n_2008;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_799;
wire n_8503;
wire n_6785;
wire n_8254;
wire n_1213;
wire n_6374;
wire n_8959;
wire n_9117;
wire n_6930;
wire n_9198;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_8506;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_7735;
wire n_8265;
wire n_8465;
wire n_1689;
wire n_8049;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_6838;
wire n_869;
wire n_5736;
wire n_401;
wire n_6937;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_1352;
wire n_10080;
wire n_2197;
wire n_7558;
wire n_2199;
wire n_8937;
wire n_5069;
wire n_7442;
wire n_8272;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_9249;
wire n_137;
wire n_294;
wire n_3968;
wire n_9398;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_684;
wire n_124;
wire n_268;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_6674;
wire n_664;
wire n_10155;
wire n_2480;
wire n_235;
wire n_6034;
wire n_7499;
wire n_2363;
wire n_643;
wire n_4072;
wire n_9751;
wire n_916;
wire n_5579;
wire n_1115;
wire n_8381;
wire n_7085;
wire n_4781;
wire n_9579;
wire n_3606;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_2550;
wire n_6762;
wire n_7341;
wire n_467;
wire n_7895;
wire n_4424;
wire n_823;
wire n_8366;
wire n_725;
wire n_8101;
wire n_7611;
wire n_9925;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_8384;
wire n_9889;
wire n_5642;
wire n_3553;
wire n_7224;
wire n_719;
wire n_5880;
wire n_8728;
wire n_6169;
wire n_4746;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_1683;
wire n_10212;
wire n_1530;
wire n_8023;
wire n_8052;
wire n_997;
wire n_7627;
wire n_9998;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_9729;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_8614;
wire n_1268;
wire n_2996;
wire n_5793;
wire n_559;
wire n_5591;
wire n_508;
wire n_7856;
wire n_1320;
wire n_4050;
wire n_9081;
wire n_7496;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_9784;
wire n_2102;
wire n_5623;
wire n_10005;
wire n_1063;
wire n_10217;
wire n_5681;
wire n_4853;
wire n_9856;
wire n_981;
wire n_9101;
wire n_7399;
wire n_867;
wire n_2422;
wire n_6213;
wire n_8656;
wire n_134;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_587;
wire n_2950;
wire n_7605;
wire n_5220;
wire n_5732;
wire n_8897;
wire n_3852;
wire n_9696;
wire n_548;
wire n_5178;
wire n_812;
wire n_6814;
wire n_4520;
wire n_7342;
wire n_518;
wire n_2057;
wire n_9825;
wire n_8014;
wire n_4008;
wire n_5507;
wire n_10093;
wire n_8564;
wire n_905;
wire n_7214;
wire n_7472;
wire n_5077;
wire n_782;
wire n_8371;
wire n_5872;
wire n_3858;
wire n_7408;
wire n_8231;
wire n_9250;
wire n_1901;
wire n_6115;
wire n_4502;
wire n_9572;
wire n_6858;
wire n_8558;
wire n_3032;
wire n_5735;
wire n_4851;
wire n_9483;
wire n_10275;
wire n_9816;
wire n_9253;
wire n_1330;
wire n_8164;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_9136;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_7837;
wire n_8357;
wire n_1745;
wire n_9426;
wire n_3924;
wire n_769;
wire n_8870;
wire n_9831;
wire n_4571;
wire n_2006;
wire n_8143;
wire n_6430;
wire n_6193;
wire n_934;
wire n_6462;
wire n_8422;
wire n_1618;
wire n_5314;
wire n_826;
wire n_2343;
wire n_3439;
wire n_9896;
wire n_9650;
wire n_10002;
wire n_5049;
wire n_6757;
wire n_654;
wire n_6822;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_570;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_6518;
wire n_9767;
wire n_6797;
wire n_2799;
wire n_4454;
wire n_7938;
wire n_8253;
wire n_4229;
wire n_1083;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_9028;
wire n_9055;
wire n_5718;
wire n_10251;
wire n_787;
wire n_6916;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_8563;
wire n_9949;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_522;
wire n_7812;
wire n_4879;
wire n_5051;
wire n_930;
wire n_181;
wire n_9684;
wire n_3926;
wire n_6152;
wire n_10010;
wire n_9724;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_8243;
wire n_1577;
wire n_10226;
wire n_8236;
wire n_8292;
wire n_2854;
wire n_386;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_5777;
wire n_2764;
wire n_7949;
wire n_1498;
wire n_8611;
wire n_7046;
wire n_4225;
wire n_682;
wire n_10020;
wire n_141;
wire n_9826;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_8011;
wire n_9839;
wire n_4300;
wire n_9399;
wire n_3551;
wire n_432;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_6589;
wire n_7579;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_8139;
wire n_140;
wire n_8123;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_7917;
wire n_5951;
wire n_7092;
wire n_2442;
wire n_6197;
wire n_6971;
wire n_9938;
wire n_928;
wire n_8424;
wire n_9776;
wire n_8859;
wire n_1943;
wire n_7460;
wire n_9658;
wire n_3117;
wire n_9605;
wire n_3428;
wire n_9013;
wire n_2961;
wire n_8730;
wire n_9417;
wire n_8156;
wire n_9290;
wire n_9212;
wire n_3351;
wire n_3527;
wire n_236;
wire n_9721;
wire n_7698;
wire n_7886;
wire n_6154;
wire n_7344;
wire n_1396;
wire n_1348;
wire n_6020;
wire n_2883;
wire n_1752;
wire n_9586;
wire n_7904;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_9104;
wire n_7079;
wire n_10225;
wire n_9293;
wire n_462;
wire n_5120;
wire n_8645;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_7774;
wire n_5797;
wire n_7922;
wire n_8189;
wire n_8618;
wire n_6696;
wire n_471;
wire n_4839;
wire n_5222;
wire n_8285;
wire n_5743;
wire n_1028;
wire n_4016;
wire n_9919;
wire n_8826;
wire n_6210;
wire n_10123;
wire n_5772;
wire n_474;
wire n_3435;
wire n_8715;
wire n_3575;
wire n_1546;
wire n_595;
wire n_8782;
wire n_6964;
wire n_10083;
wire n_5801;
wire n_6117;
wire n_632;
wire n_4231;
wire n_8117;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_7670;
wire n_4923;
wire n_3652;
wire n_9445;
wire n_4097;
wire n_170;
wire n_6681;
wire n_161;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_8497;
wire n_745;
wire n_9930;
wire n_2381;
wire n_6661;
wire n_8018;
wire n_3303;
wire n_1654;
wire n_6640;
wire n_3916;
wire n_7940;
wire n_2569;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_6455;
wire n_2196;
wire n_3591;
wire n_7721;
wire n_9727;
wire n_4273;
wire n_3024;
wire n_7606;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_6832;
wire n_8798;
wire n_7836;
wire n_1595;
wire n_2161;
wire n_6160;
wire n_7564;
wire n_2404;
wire n_2083;
wire n_7884;
wire n_8673;
wire n_6718;
wire n_9685;
wire n_2503;
wire n_8502;
wire n_6542;
wire n_10126;
wire n_1540;
wire n_1936;
wire n_6031;
wire n_5568;
wire n_2027;
wire n_5502;
wire n_453;
wire n_403;
wire n_9421;
wire n_2642;
wire n_8577;
wire n_720;
wire n_2500;
wire n_7653;
wire n_10092;
wire n_1918;
wire n_5656;
wire n_863;
wire n_8531;
wire n_8635;
wire n_6763;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_9567;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_9298;
wire n_2414;
wire n_10116;
wire n_6438;
wire n_10048;
wire n_9059;
wire n_1402;
wire n_8485;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_8872;
wire n_644;
wire n_2229;
wire n_8752;
wire n_1397;
wire n_9396;
wire n_4596;
wire n_6758;
wire n_5413;
wire n_2004;
wire n_7976;
wire n_9234;
wire n_9425;
wire n_5412;
wire n_251;
wire n_9620;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_10191;
wire n_6874;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_8341;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_334;
wire n_811;
wire n_6030;
wire n_8521;
wire n_8199;
wire n_6077;
wire n_8005;
wire n_175;
wire n_4119;
wire n_3799;
wire n_7743;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_9280;
wire n_9517;
wire n_4474;
wire n_1089;
wire n_6386;
wire n_9639;
wire n_9192;
wire n_9102;
wire n_5217;
wire n_1004;
wire n_10003;
wire n_10025;
wire n_242;
wire n_8016;
wire n_10156;
wire n_8669;
wire n_5957;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_8283;
wire n_3585;
wire n_2975;
wire n_7655;
wire n_5490;
wire n_438;
wire n_5029;
wire n_8291;
wire n_2704;
wire n_4214;
wire n_8176;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7737;
wire n_10179;
wire n_7433;
wire n_533;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_278;
wire n_7347;
wire n_8145;
wire n_9487;
wire n_10268;
wire n_4580;
wire n_6792;
wire n_7633;
wire n_1263;
wire n_6177;
wire n_5912;
wire n_611;
wire n_1126;
wire n_7798;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_1859;
wire n_9221;
wire n_1677;
wire n_5557;
wire n_7397;
wire n_7389;
wire n_5472;
wire n_7602;
wire n_2955;
wire n_4112;
wire n_8069;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_7554;
wire n_4138;
wire n_5396;
wire n_7693;
wire n_552;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_8888;
wire n_1198;
wire n_6557;
wire n_7300;
wire n_956;
wire n_423;
wire n_9566;
wire n_9578;
wire n_8483;
wire n_8797;
wire n_2134;
wire n_5960;
wire n_8041;
wire n_8605;
wire n_4236;
wire n_2185;
wire n_9868;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_7532;
wire n_9292;
wire n_5143;
wire n_7724;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_6917;
wire n_7510;
wire n_6142;
wire n_1545;
wire n_2374;
wire n_5859;
wire n_173;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_8760;
wire n_854;
wire n_1799;
wire n_2396;
wire n_4734;
wire n_8928;
wire n_10004;
wire n_8374;
wire n_674;
wire n_1939;
wire n_2486;
wire n_8917;
wire n_6163;
wire n_516;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_7118;
wire n_1869;
wire n_8006;
wire n_4013;
wire n_606;
wire n_3039;
wire n_275;
wire n_9884;
wire n_2011;
wire n_6778;
wire n_7946;
wire n_6285;
wire n_8723;
wire n_9857;
wire n_6025;
wire n_8957;
wire n_7257;
wire n_4242;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_10140;
wire n_150;
wire n_3036;
wire n_10013;
wire n_7933;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_8409;
wire n_9815;
wire n_9110;
wire n_7669;
wire n_5268;
wire n_10110;
wire n_6318;
wire n_10133;
wire n_8215;
wire n_8220;
wire n_9471;
wire n_9048;
wire n_191;
wire n_1705;
wire n_659;
wire n_4561;
wire n_2639;
wire n_7927;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_8629;
wire n_3880;
wire n_5122;
wire n_7910;
wire n_1261;
wire n_6315;
wire n_938;
wire n_3186;
wire n_7970;
wire n_4955;
wire n_1154;
wire n_8407;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_406;
wire n_546;
wire n_1280;
wire n_9394;
wire n_3650;
wire n_8991;
wire n_291;
wire n_5840;
wire n_2761;
wire n_257;
wire n_6343;
wire n_10186;
wire n_3157;
wire n_709;
wire n_9191;
wire n_2537;
wire n_9004;
wire n_2144;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_920;
wire n_2515;
wire n_7865;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_6886;
wire n_976;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_8783;
wire n_6912;
wire n_8326;
wire n_5914;
wire n_775;
wire n_8504;
wire n_8445;
wire n_8250;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_9118;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_8408;
wire n_4543;
wire n_2099;
wire n_10120;
wire n_4941;
wire n_7252;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_9051;
wire n_7133;
wire n_1850;
wire n_163;
wire n_6883;
wire n_243;
wire n_5519;
wire n_9908;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_215;
wire n_350;
wire n_196;
wire n_7061;
wire n_8155;
wire n_6009;
wire n_8818;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_7518;
wire n_9123;
wire n_5586;
wire n_580;
wire n_2693;
wire n_10232;
wire n_4065;
wire n_3798;
wire n_6378;
wire n_8660;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_8275;
wire n_1218;
wire n_9327;
wire n_2632;
wire n_6601;
wire n_7216;
wire n_5771;
wire n_475;
wire n_1547;
wire n_777;
wire n_6407;
wire n_9687;
wire n_1755;
wire n_8297;
wire n_9828;
wire n_6749;
wire n_6839;
wire n_415;
wire n_485;
wire n_9519;
wire n_7711;
wire n_958;
wire n_2908;
wire n_10089;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_7705;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_8590;
wire n_4942;
wire n_6217;
wire n_164;
wire n_6680;
wire n_5844;
wire n_2432;
wire n_7972;
wire n_1521;
wire n_6532;
wire n_3405;
wire n_214;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_8072;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7854;
wire n_7614;
wire n_2337;
wire n_7707;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_8050;
wire n_6736;
wire n_5344;
wire n_923;
wire n_6526;
wire n_8142;
wire n_6339;
wire n_4629;
wire n_213;
wire n_2932;
wire n_2980;
wire n_464;
wire n_5225;
wire n_8151;
wire n_6350;
wire n_7013;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_9802;
wire n_9315;
wire n_9296;
wire n_8599;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_10022;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_460;
wire n_4376;
wire n_3986;
wire n_10031;
wire n_5705;
wire n_4753;
wire n_571;
wire n_4552;
wire n_7656;
wire n_3885;
wire n_6845;
wire n_9405;
wire n_9302;
wire n_7105;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_10166;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_5574;
wire n_5126;
wire n_1039;
wire n_6508;
wire n_2214;
wire n_9842;
wire n_9977;
wire n_2055;
wire n_3427;
wire n_9887;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4176;
wire n_4042;
wire n_7570;
wire n_8246;
wire n_9524;
wire n_7771;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_2688;
wire n_5368;
wire n_9322;
wire n_1202;
wire n_10098;
wire n_10042;
wire n_8057;
wire n_9122;
wire n_8349;
wire n_5626;
wire n_9333;
wire n_8743;
wire n_6603;
wire n_6114;
wire n_1463;
wire n_9590;
wire n_6576;
wire n_3651;
wire n_7943;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_8473;
wire n_7208;
wire n_6245;
wire n_2865;
wire n_349;
wire n_2706;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_9676;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_7714;
wire n_9902;
wire n_10054;
wire n_627;
wire n_8535;
wire n_4815;
wire n_9621;
wire n_7202;
wire n_9140;
wire n_9604;
wire n_3580;
wire n_4246;
wire n_7011;
wire n_2139;
wire n_4609;
wire n_7621;
wire n_8068;
wire n_5291;
wire n_9821;
wire n_5876;
wire n_10178;
wire n_6970;
wire n_5114;
wire n_2674;
wire n_6409;
wire n_6704;
wire n_1565;
wire n_4088;
wire n_6876;
wire n_7778;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_9343;
wire n_7028;
wire n_4462;
wire n_4472;
wire n_647;
wire n_3433;
wire n_7320;
wire n_7313;
wire n_6255;
wire n_7343;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_7525;
wire n_2450;
wire n_7875;
wire n_561;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_6938;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_8785;
wire n_9952;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_8327;
wire n_9219;
wire n_7337;
wire n_6989;
wire n_8512;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_3989;
wire n_4475;
wire n_7753;
wire n_10076;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_8168;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_8392;
wire n_7038;
wire n_4683;
wire n_5366;
wire n_728;
wire n_1162;
wire n_272;
wire n_10132;
wire n_9872;
wire n_1847;
wire n_2767;
wire n_6360;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_9553;
wire n_3602;
wire n_2967;
wire n_409;
wire n_6146;
wire n_887;
wire n_9447;
wire n_6270;
wire n_9150;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_300;
wire n_9592;
wire n_5451;
wire n_9984;
wire n_3923;
wire n_931;
wire n_599;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_8419;
wire n_639;
wire n_5086;
wire n_9814;
wire n_1629;
wire n_2801;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_9446;
wire n_4905;
wire n_2763;
wire n_360;
wire n_10023;
wire n_10211;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_9461;
wire n_9793;
wire n_1997;
wire n_6691;
wire n_3748;
wire n_8997;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_187;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_9874;
wire n_7392;
wire n_2215;
wire n_5053;
wire n_7912;
wire n_8245;
wire n_1259;
wire n_6239;
wire n_4553;
wire n_706;
wire n_746;
wire n_6803;
wire n_7919;
wire n_784;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_4809;
wire n_8109;
wire n_5226;
wire n_1244;
wire n_7657;
wire n_1925;
wire n_3660;
wire n_7995;
wire n_1815;
wire n_6048;
wire n_5867;
wire n_8985;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_913;
wire n_6773;
wire n_9403;
wire n_3833;
wire n_5632;
wire n_865;
wire n_8390;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_6336;
wire n_3814;
wire n_8463;
wire n_7041;
wire n_1415;
wire n_2592;
wire n_7802;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_10181;
wire n_10074;
wire n_9731;
wire n_5660;
wire n_4645;
wire n_1191;
wire n_7557;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_6776;
wire n_284;
wire n_3128;
wire n_5426;
wire n_9947;
wire n_6463;
wire n_744;
wire n_629;
wire n_2631;
wire n_7896;
wire n_2178;
wire n_1767;
wire n_9699;
wire n_6372;
wire n_9305;
wire n_7176;
wire n_10220;
wire n_1529;
wire n_8517;
wire n_2469;
wire n_5778;
wire n_5625;
wire n_6396;
wire n_3355;
wire n_9218;
wire n_604;
wire n_2007;
wire n_3917;
wire n_6669;
wire n_9096;
wire n_3942;
wire n_10170;
wire n_10142;
wire n_2736;
wire n_3765;
wire n_498;
wire n_5531;
wire n_9534;
wire n_7826;
wire n_3000;
wire n_252;
wire n_624;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_936;
wire n_1500;
wire n_9164;
wire n_9546;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_7590;
wire n_259;
wire n_448;
wire n_999;
wire n_9358;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_8208;
wire n_1933;
wire n_6995;
wire n_7185;
wire n_1656;
wire n_10127;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_9730;
wire n_6254;
wire n_563;
wire n_6161;
wire n_9066;
wire n_3457;
wire n_9185;
wire n_204;
wire n_1678;
wire n_9318;
wire n_8134;
wire n_7987;
wire n_4324;
wire n_4821;
wire n_8631;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_8694;
wire n_8965;
wire n_8647;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_908;
wire n_6128;
wire n_4086;
wire n_2412;
wire n_7037;
wire n_4814;
wire n_724;
wire n_2084;
wire n_1781;
wire n_3648;
wire n_5749;
wire n_8427;
wire n_3075;
wire n_3173;
wire n_9339;
wire n_5332;
wire n_9596;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_456;
wire n_959;
wire n_3031;
wire n_10006;
wire n_7258;
wire n_7432;
wire n_9156;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_6334;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_8984;
wire n_6848;
wire n_8345;
wire n_2171;
wire n_9973;
wire n_4708;
wire n_6321;
wire n_7765;
wire n_2768;
wire n_2314;
wire n_9708;
wire n_9268;
wire n_8764;
wire n_6794;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_10245;
wire n_514;
wire n_1079;
wire n_7761;
wire n_7197;
wire n_5489;
wire n_1593;
wire n_6400;
wire n_3767;
wire n_442;
wire n_2299;
wire n_131;
wire n_2540;
wire n_2873;
wire n_4589;
wire n_5057;
wire n_9097;
wire n_10280;
wire n_4578;
wire n_1640;
wire n_6705;
wire n_7775;
wire n_9636;
wire n_10256;
wire n_2162;
wire n_7619;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_185;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_8083;
wire n_3502;
wire n_8853;
wire n_3098;
wire n_1383;
wire n_6495;
wire n_5013;
wire n_2312;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_9473;
wire n_3015;
wire n_1171;
wire n_10145;
wire n_9560;
wire n_1920;
wire n_1065;
wire n_5569;
wire n_8038;
wire n_9175;
wire n_8711;
wire n_5439;
wire n_8229;
wire n_8949;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_6481;
wire n_9810;
wire n_3607;
wire n_7548;
wire n_4925;
wire n_9244;
wire n_9584;
wire n_1921;
wire n_1309;
wire n_6534;
wire n_4974;
wire n_8567;
wire n_9439;
wire n_355;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_8655;
wire n_2571;
wire n_1286;
wire n_9235;
wire n_6181;
wire n_1177;
wire n_3276;
wire n_6728;
wire n_8705;
wire n_9043;
wire n_9768;
wire n_3787;
wire n_5119;
wire n_9037;
wire n_2124;
wire n_5715;
wire n_9085;
wire n_8085;
wire n_8777;
wire n_6133;
wire n_8852;
wire n_9264;
wire n_6528;
wire n_10114;
wire n_7604;
wire n_613;
wire n_7407;
wire n_1119;
wire n_1240;
wire n_8185;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_8513;
wire n_6670;
wire n_6774;
wire n_8365;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_361;
wire n_6741;
wire n_7424;
wire n_700;
wire n_6038;
wire n_573;
wire n_4818;
wire n_7727;
wire n_4514;
wire n_388;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_9550;
wire n_9836;
wire n_3248;
wire n_2277;
wire n_6282;
wire n_1568;
wire n_9929;
wire n_2110;
wire n_274;
wire n_8035;
wire n_8505;
wire n_582;
wire n_1332;
wire n_4433;
wire n_8874;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_10008;
wire n_3153;
wire n_6700;
wire n_512;
wire n_7334;
wire n_1591;
wire n_2033;
wire n_7755;
wire n_7684;
wire n_4341;
wire n_8098;
wire n_9187;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_5932;
wire n_6178;
wire n_1111;
wire n_2132;
wire n_6234;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_9406;
wire n_609;
wire n_3838;
wire n_9342;
wire n_1909;
wire n_4277;
wire n_7787;
wire n_4140;
wire n_8067;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_7849;
wire n_5186;
wire n_7367;
wire n_8619;
wire n_9851;
wire n_9559;
wire n_8679;
wire n_9806;
wire n_8644;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_6715;
wire n_5828;
wire n_2831;
wire n_7200;
wire n_1456;
wire n_9860;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_6337;
wire n_261;
wire n_4868;
wire n_8923;
wire n_8970;
wire n_1885;
wire n_8332;
wire n_10119;
wire n_2452;
wire n_8632;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_8876;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_10067;
wire n_4059;
wire n_8856;
wire n_2455;
wire n_9240;
wire n_4595;
wire n_7877;
wire n_1849;
wire n_8945;
wire n_1131;
wire n_8918;
wire n_7799;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_5631;
wire n_8028;
wire n_2467;
wire n_6539;
wire n_1094;
wire n_7243;
wire n_7179;
wire n_2288;
wire n_9345;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_10222;
wire n_346;
wire n_1209;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_602;
wire n_4888;
wire n_7274;
wire n_8774;
wire n_5326;
wire n_1435;
wire n_8779;
wire n_879;
wire n_3394;
wire n_8968;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_8404;
wire n_4669;
wire n_405;
wire n_4339;
wire n_6595;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_7738;
wire n_4060;
wire n_996;
wire n_9223;
wire n_2658;
wire n_9499;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_327;
wire n_8073;
wire n_135;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_7785;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_7373;
wire n_9576;
wire n_9120;
wire n_3589;
wire n_10097;
wire n_952;
wire n_2534;
wire n_1229;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_9651;
wire n_6257;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_9386;
wire n_2989;
wire n_6852;
wire n_2789;
wire n_6346;
wire n_4775;
wire n_9779;
wire n_2216;
wire n_531;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_764;
wire n_1424;
wire n_162;
wire n_5365;
wire n_2933;
wire n_7587;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_7874;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_2328;
wire n_199;
wire n_7760;
wire n_4248;
wire n_9635;
wire n_5915;
wire n_6818;
wire n_9444;
wire n_5452;
wire n_7226;
wire n_8930;
wire n_4754;
wire n_7057;
wire n_7685;
wire n_8031;
wire n_8750;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6815;
wire n_6753;
wire n_9364;
wire n_9581;
wire n_9512;
wire n_3053;
wire n_1299;
wire n_9317;
wire n_3893;
wire n_8593;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_418;
wire n_7730;
wire n_315;
wire n_451;
wire n_8509;
wire n_9314;
wire n_9459;
wire n_8405;
wire n_1699;
wire n_3334;
wire n_9549;
wire n_7913;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_8492;
wire n_6764;
wire n_397;
wire n_5535;
wire n_1432;
wire n_9275;
wire n_3875;
wire n_10210;
wire n_5370;
wire n_7706;
wire n_7891;
wire n_6391;
wire n_4003;
wire n_8088;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_9865;
wire n_6471;
wire n_1844;
wire n_3777;
wire n_6627;
wire n_10027;
wire n_5761;
wire n_10263;
wire n_4784;
wire n_7203;
wire n_8429;
wire n_8854;
wire n_9757;
wire n_2999;
wire n_7512;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_9656;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_7215;
wire n_5209;
wire n_10246;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_7388;
wire n_7694;
wire n_1179;
wire n_6243;
wire n_753;
wire n_6488;
wire n_1048;
wire n_4286;
wire n_9629;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_8686;
wire n_6457;
wire n_4470;
wire n_2236;
wire n_330;
wire n_2816;
wire n_692;
wire n_7982;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_8773;
wire n_8225;
wire n_8583;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_6867;
wire n_8887;
wire n_3417;
wire n_9556;
wire n_1143;
wire n_1579;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_9259;
wire n_9995;
wire n_1688;
wire n_6633;
wire n_9371;
wire n_492;
wire n_8080;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_10050;
wire n_5275;
wire n_4689;
wire n_341;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_2755;
wire n_8964;
wire n_5989;
wire n_543;
wire n_3237;
wire n_9008;
wire n_6574;
wire n_8929;
wire n_8539;
wire n_1992;
wire n_6395;
wire n_4402;
wire n_9484;
wire n_8745;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_7996;
wire n_6233;
wire n_449;
wire n_4550;
wire n_6456;
wire n_1400;
wire n_1214;
wire n_1342;
wire n_8588;
wire n_8554;
wire n_8776;
wire n_9319;
wire n_3382;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_9442;
wire n_10165;
wire n_2169;
wire n_7198;
wire n_1557;
wire n_4201;
wire n_8802;
wire n_9587;
wire n_6784;
wire n_6168;
wire n_9904;
wire n_618;
wire n_9157;
wire n_896;
wire n_8431;
wire n_8453;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_356;
wire n_3099;
wire n_8955;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_8634;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_2192;
wire n_8896;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_7950;
wire n_7249;
wire n_9713;
wire n_2670;
wire n_1646;
wire n_9452;
wire n_10104;
wire n_1307;
wire n_5947;
wire n_7336;
wire n_8837;
wire n_4416;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_814;
wire n_2707;
wire n_8907;
wire n_6799;
wire n_10115;
wire n_8015;
wire n_9974;
wire n_5920;
wire n_6672;
wire n_2471;
wire n_1472;
wire n_6149;
wire n_1671;
wire n_8256;
wire n_10065;
wire n_10243;
wire n_10087;
wire n_7142;
wire n_3230;
wire n_5808;
wire n_1062;
wire n_3342;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_7916;
wire n_6450;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_5353;
wire n_3729;
wire n_8074;
wire n_4978;
wire n_4690;
wire n_10174;
wire n_10266;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_8778;
wire n_783;
wire n_1928;
wire n_8039;
wire n_5244;
wire n_6523;
wire n_5382;
wire n_8065;
wire n_1188;
wire n_6107;
wire n_9634;
wire n_3957;
wire n_6775;
wire n_5274;
wire n_3848;
wire n_8194;
wire n_4284;
wire n_2600;
wire n_8207;
wire n_3919;
wire n_10106;
wire n_9241;
wire n_336;
wire n_6232;
wire n_6445;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_9903;
wire n_3608;
wire n_8582;
wire n_510;
wire n_216;
wire n_6056;
wire n_8537;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_9615;
wire n_3177;
wire n_4053;
wire n_8951;
wire n_7759;
wire n_9600;
wire n_2352;
wire n_7818;
wire n_9748;
wire n_9945;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_9927;
wire n_5587;
wire n_2619;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_8217;
wire n_10046;
wire n_241;
wire n_1110;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_1088;
wire n_8437;
wire n_5249;
wire n_3393;
wire n_8849;
wire n_638;
wire n_7447;
wire n_866;
wire n_7944;
wire n_5198;
wire n_5360;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_9295;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_249;
wire n_6252;
wire n_5866;
wire n_6493;
wire n_8568;
wire n_10239;
wire n_577;
wire n_7947;
wire n_4005;
wire n_9916;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_8980;
wire n_5899;
wire n_7629;
wire n_8051;
wire n_693;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_8716;
wire n_3812;
wire n_9844;
wire n_1886;
wire n_1389;
wire n_7601;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_7757;
wire n_8030;
wire n_9316;
wire n_9663;
wire n_10168;
wire n_306;
wire n_5865;
wire n_10075;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_10068;
wire n_10276;
wire n_3093;
wire n_1843;
wire n_8749;
wire n_3061;
wire n_7138;
wire n_7290;
wire n_8544;
wire n_8249;
wire n_1597;
wire n_9628;
wire n_1659;
wire n_2431;
wire n_6679;
wire n_8496;
wire n_9789;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_7625;
wire n_5822;
wire n_2564;
wire n_9299;
wire n_6259;
wire n_4947;
wire n_876;
wire n_7284;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_6390;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_206;
wire n_7971;
wire n_3174;
wire n_982;
wire n_9022;
wire n_1453;
wire n_2217;
wire n_6630;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_9427;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_6279;
wire n_8698;
wire n_1514;
wire n_8695;
wire n_1771;
wire n_9344;
wire n_557;
wire n_8751;
wire n_1005;
wire n_607;
wire n_679;
wire n_710;
wire n_3090;
wire n_527;
wire n_1168;
wire n_2437;
wire n_3762;
wire n_6813;
wire n_9764;
wire n_5564;
wire n_8273;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_177;
wire n_9242;
wire n_9498;
wire n_8442;
wire n_1988;
wire n_7106;
wire n_8472;
wire n_9535;
wire n_6042;
wire n_7644;
wire n_1853;
wire n_1356;
wire n_6057;
wire n_1787;
wire n_4137;
wire n_7529;
wire n_8986;
wire n_10011;
wire n_6675;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_6476;
wire n_8200;
wire n_3972;
wire n_10055;
wire n_7907;
wire n_125;
wire n_8188;
wire n_8528;
wire n_6207;
wire n_529;
wire n_5539;
wire n_126;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_202;
wire n_9088;
wire n_3308;
wire n_6524;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_8920;
wire n_8267;
wire n_1720;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_159;
wire n_4653;
wire n_9734;
wire n_9505;
wire n_9664;
wire n_2354;
wire n_2246;
wire n_7199;
wire n_5273;
wire n_10262;
wire n_8360;
wire n_4677;
wire n_3901;
wire n_715;
wire n_8036;
wire n_9510;
wire n_1480;
wire n_5261;
wire n_6520;
wire n_7853;
wire n_7648;
wire n_9413;
wire n_9888;
wire n_3757;
wire n_8393;
wire n_8821;
wire n_9863;
wire n_8160;
wire n_9199;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_9014;
wire n_10204;
wire n_9411;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_9336;
wire n_9360;
wire n_9543;
wire n_810;
wire n_2965;
wire n_416;
wire n_3635;
wire n_6024;
wire n_7866;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_1170;
wire n_305;
wire n_2213;
wire n_6425;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_7638;
wire n_8833;
wire n_5703;
wire n_8240;
wire n_4634;
wire n_3337;
wire n_7988;
wire n_2527;
wire n_9404;
wire n_8579;
wire n_855;
wire n_5534;
wire n_6432;
wire n_1461;
wire n_9678;
wire n_3204;
wire n_8258;
wire n_9854;
wire n_7259;
wire n_8626;
wire n_2136;
wire n_6540;
wire n_6955;
wire n_9481;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_9672;
wire n_3129;
wire n_9893;
wire n_4126;
wire n_1282;
wire n_7237;
wire n_1783;
wire n_8935;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_6388;
wire n_10240;
wire n_5904;
wire n_9478;
wire n_4880;
wire n_9266;
wire n_9813;
wire n_6760;
wire n_1907;
wire n_501;
wire n_2686;
wire n_8009;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_5750;
wire n_5572;
wire n_7063;
wire n_10205;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_9042;
wire n_2906;
wire n_4943;
wire n_382;
wire n_2187;
wire n_8012;
wire n_7576;
wire n_9506;
wire n_8608;
wire n_1762;
wire n_1013;
wire n_718;
wire n_8008;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_8079;
wire n_6664;
wire n_5815;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_9666;
wire n_3104;
wire n_10112;
wire n_612;
wire n_6487;
wire n_9146;
wire n_4737;
wire n_7734;
wire n_6729;
wire n_3647;
wire n_10056;
wire n_9862;
wire n_5755;
wire n_825;
wire n_9274;
wire n_2819;
wire n_8702;
wire n_5949;
wire n_506;
wire n_737;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_7858;
wire n_1715;
wire n_9619;
wire n_1952;
wire n_4393;
wire n_7385;
wire n_3720;
wire n_8576;
wire n_9508;
wire n_4535;
wire n_10105;
wire n_7668;
wire n_733;
wire n_8662;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_7476;
wire n_5955;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_792;
wire n_8436;
wire n_9987;
wire n_8124;
wire n_8148;
wire n_8033;
wire n_6843;
wire n_3140;
wire n_7953;
wire n_8343;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_8118;
wire n_298;
wire n_2104;
wire n_505;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_4196;
wire n_6969;
wire n_8741;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5665;
wire n_6485;
wire n_5340;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5783;
wire n_8478;
wire n_5183;
wire n_7082;
wire n_6075;
wire n_9569;
wire n_3084;
wire n_6120;
wire n_1727;
wire n_6659;
wire n_2735;
wire n_6750;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_9935;
wire n_1046;
wire n_9707;
wire n_8376;
wire n_3761;
wire n_9827;
wire n_7689;
wire n_4889;
wire n_7132;
wire n_2014;
wire n_8763;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_7824;
wire n_8996;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_9007;
wire n_4828;
wire n_9797;
wire n_6003;
wire n_5385;
wire n_8726;
wire n_8799;
wire n_4558;
wire n_7796;
wire n_9053;
wire n_6478;
wire n_2172;
wire n_6066;
wire n_9450;
wire n_7034;
wire n_6086;
wire n_9121;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_1129;
wire n_8303;
wire n_8796;
wire n_158;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_10088;
wire n_961;
wire n_2250;
wire n_7084;
wire n_276;
wire n_5845;
wire n_9617;
wire n_9089;
wire n_8883;
wire n_7293;
wire n_1225;
wire n_169;
wire n_8251;
wire n_10247;
wire n_9236;
wire n_400;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_7253;
wire n_2423;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_9493;
wire n_8860;
wire n_994;
wire n_8003;
wire n_6410;
wire n_3344;
wire n_2194;
wire n_848;
wire n_5973;
wire n_4465;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_8524;
wire n_6059;
wire n_5130;
wire n_1567;
wire n_8914;
wire n_7520;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_8520;
wire n_9490;
wire n_3842;
wire n_6103;
wire n_145;
wire n_6809;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_631;
wire n_479;
wire n_6267;
wire n_8165;
wire n_9525;
wire n_1797;
wire n_2957;
wire n_9127;
wire n_9119;
wire n_5855;
wire n_9002;
wire n_10069;
wire n_2357;
wire n_1250;
wire n_8330;
wire n_8682;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_7918;
wire n_6610;
wire n_608;
wire n_10259;
wire n_8467;
wire n_8775;
wire n_8886;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_8696;
wire n_1589;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7514;
wire n_7163;
wire n_7620;
wire n_9867;
wire n_1086;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_5473;
wire n_4612;
wire n_3754;
wire n_1469;
wire n_5946;
wire n_10197;
wire n_2744;
wire n_6711;
wire n_8464;
wire n_4287;
wire n_2397;
wire n_7445;
wire n_384;
wire n_2208;
wire n_6847;
wire n_9131;
wire n_3063;
wire n_9790;
wire n_5177;
wire n_3617;
wire n_7123;
wire n_6384;
wire n_333;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_8720;
wire n_4505;
wire n_7959;
wire n_1676;
wire n_258;
wire n_1113;
wire n_9611;
wire n_7563;
wire n_6298;
wire n_1277;
wire n_2591;
wire n_9032;
wire n_188;
wire n_9428;
wire n_3384;
wire n_9990;
wire n_7361;
wire n_852;
wire n_4602;
wire n_5172;
wire n_8186;
wire n_4449;
wire n_9705;
wire n_1864;
wire n_8890;
wire n_7322;
wire n_8219;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_9774;
wire n_463;
wire n_5070;
wire n_502;
wire n_6377;
wire n_466;
wire n_420;
wire n_1337;
wire n_4445;
wire n_699;
wire n_5566;
wire n_5414;
wire n_8738;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_465;
wire n_2832;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_273;
wire n_3181;
wire n_6348;
wire n_7713;
wire n_616;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_6834;
wire n_10124;
wire n_5313;
wire n_3323;
wire n_9374;
wire n_2734;
wire n_4914;
wire n_9792;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_1076;
wire n_2823;
wire n_1408;
wire n_494;
wire n_1761;
wire n_8066;
wire n_5874;
wire n_7977;
wire n_730;
wire n_8342;
wire n_7508;
wire n_9771;
wire n_9712;
wire n_7021;
wire n_354;
wire n_5270;
wire n_5956;
wire n_7834;
wire n_795;
wire n_4345;
wire n_5188;
wire n_9905;
wire n_180;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_6078;
wire n_7000;
wire n_8571;
wire n_9163;
wire n_9308;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_10038;
wire n_7921;
wire n_8877;
wire n_2655;
wire n_4185;
wire n_8862;
wire n_10144;
wire n_8402;
wire n_4797;
wire n_2366;
wire n_7130;
wire n_1526;
wire n_10176;
wire n_5823;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_9387;
wire n_7538;
wire n_712;
wire n_7517;
wire n_1583;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_7077;
wire n_285;
wire n_412;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_6642;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_7333;
wire n_4364;
wire n_4928;
wire n_4245;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_597;
wire n_3406;
wire n_3604;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_9847;
wire n_5934;
wire n_6942;
wire n_8418;
wire n_2019;
wire n_10227;
wire n_1340;
wire n_1558;
wire n_9577;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_262;
wire n_8805;
wire n_9111;
wire n_1704;
wire n_6511;
wire n_3721;
wire n_1254;
wire n_6507;
wire n_1026;
wire n_2026;
wire n_9513;
wire n_1234;
wire n_2109;
wire n_364;
wire n_2013;
wire n_1990;
wire n_9853;
wire n_1032;
wire n_2614;
wire n_7319;
wire n_7997;
wire n_2991;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_9130;
wire n_2242;
wire n_2752;
wire n_9941;
wire n_2894;
wire n_9135;
wire n_6606;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_8144;
wire n_3699;
wire n_5067;
wire n_7107;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_7469;
wire n_2728;
wire n_3857;
wire n_8111;

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_22),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_53),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_59),
.Y(n_131)
);

INVx4_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_34),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_55),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_29),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_26),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_71),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_10),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_31),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_38),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_17),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_35),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_52),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_92),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_98),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_37),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_3),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_18),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_43),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_39),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_91),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_64),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_16),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_42),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_57),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_46),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_48),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_68),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_14),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_24),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_56),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_0),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_58),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_24),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_51),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_45),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_3),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_110),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_109),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_16),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_108),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_13),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_8),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_10),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_4),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_28),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_30),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_17),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_4),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_65),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_96),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_101),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_100),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_73),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_74),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_90),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_20),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_13),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_118),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_40),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_47),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_25),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_77),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_94),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_22),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_72),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_62),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_113),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_15),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_11),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_1),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_81),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_70),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_7),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_21),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_154),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_154),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_123),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_131),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_135),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_134),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_156),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_187),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_128),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_142),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_175),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_146),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_252),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_259),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_124),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_259),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_267),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_268),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_272),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_273),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_274),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_274),
.Y(n_315)
);

BUFx6f_ASAP7_75t_SL g316 ( 
.A(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_134),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_287),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_203),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_263),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_238),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_160),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_238),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_160),
.Y(n_338)
);

NAND2x1p5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_235),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_303),
.A2(n_201),
.B1(n_125),
.B2(n_242),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_280),
.A2(n_136),
.B1(n_167),
.B2(n_217),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_255),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_302),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_283),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_312),
.A2(n_250),
.B(n_248),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_260),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_314),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_199),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_260),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_263),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_284),
.B(n_261),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_282),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_282),
.B(n_261),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_286),
.B(n_265),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_286),
.Y(n_364)
);

OAI21x1_ASAP7_75t_L g365 ( 
.A1(n_289),
.A2(n_248),
.B(n_250),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_289),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_292),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_279),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_279),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_279),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_279),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_283),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g375 ( 
.A(n_304),
.B(n_199),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_279),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_279),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_279),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_304),
.B(n_275),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_304),
.B(n_265),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_279),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_287),
.B(n_248),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_279),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_290),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_279),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_287),
.B(n_250),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_279),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_290),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_283),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_279),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_283),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_279),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_L g393 ( 
.A(n_300),
.B(n_205),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_279),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_279),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_279),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_283),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_290),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_283),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_304),
.B(n_276),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_279),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_290),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_279),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_291),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_304),
.B(n_276),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_283),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_279),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_283),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g409 ( 
.A(n_304),
.B(n_176),
.Y(n_409)
);

CKINVDCx6p67_ASAP7_75t_R g410 ( 
.A(n_292),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_283),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_287),
.B(n_150),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_301),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_283),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_297),
.B(n_168),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_279),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_279),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_283),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_279),
.Y(n_419)
);

OAI22x1_ASAP7_75t_R g420 ( 
.A1(n_283),
.A2(n_201),
.B1(n_171),
.B2(n_221),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_297),
.B(n_192),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_279),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_299),
.A2(n_195),
.B1(n_200),
.B2(n_237),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_279),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_283),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_304),
.B(n_278),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_279),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_290),
.B(n_278),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_283),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_279),
.Y(n_430)
);

NAND2x1p5_ASAP7_75t_L g431 ( 
.A(n_290),
.B(n_126),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_297),
.A2(n_211),
.B1(n_157),
.B2(n_240),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_279),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_287),
.B(n_139),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_290),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_304),
.B(n_137),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_279),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_382),
.A2(n_266),
.B(n_264),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_319),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_384),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_428),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_319),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_402),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_324),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_324),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_326),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_320),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_326),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g453 ( 
.A1(n_345),
.A2(n_236),
.B1(n_241),
.B2(n_127),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_322),
.B(n_152),
.Y(n_454)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_386),
.A2(n_266),
.B(n_264),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_333),
.Y(n_457)
);

CKINVDCx6p67_ASAP7_75t_R g458 ( 
.A(n_410),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_325),
.Y(n_459)
);

NOR2x1p5_ASAP7_75t_L g460 ( 
.A(n_343),
.B(n_153),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_333),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_320),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_366),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_161),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_337),
.C(n_329),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_362),
.B(n_170),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_320),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_359),
.B(n_264),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_377),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_365),
.A2(n_172),
.B(n_231),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_321),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_380),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_378),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_409),
.B(n_141),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_334),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_345),
.B(n_173),
.Y(n_477)
);

AND3x2_ASAP7_75t_L g478 ( 
.A(n_367),
.B(n_185),
.C(n_143),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_336),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_340),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_318),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_365),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_341),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_318),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_392),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_380),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_379),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_355),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_347),
.B(n_194),
.C(n_186),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_318),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

BUFx6f_ASAP7_75t_SL g497 ( 
.A(n_375),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_322),
.B(n_330),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_355),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_409),
.B(n_145),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_344),
.B(n_147),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_366),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

BUFx6f_ASAP7_75t_SL g506 ( 
.A(n_375),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_407),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_344),
.B(n_151),
.Y(n_511)
);

AND2x2_ASAP7_75t_SL g512 ( 
.A(n_393),
.B(n_344),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_400),
.B(n_191),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_426),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVx8_ASAP7_75t_L g518 ( 
.A(n_355),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_344),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_437),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_370),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_322),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_330),
.B(n_133),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_321),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_330),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_369),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_351),
.B(n_158),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_351),
.B(n_159),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_364),
.B(n_169),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_369),
.Y(n_531)
);

AO21x2_ASAP7_75t_L g532 ( 
.A1(n_393),
.A2(n_196),
.B(n_225),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_369),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_355),
.B(n_205),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_371),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_318),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_376),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_356),
.B(n_197),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_376),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_376),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_144),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_422),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_351),
.B(n_162),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_372),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_331),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_373),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_356),
.B(n_198),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_398),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_381),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_383),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_390),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_394),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_395),
.B(n_148),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_396),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_403),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_343),
.B(n_206),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_351),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_331),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_416),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_417),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_348),
.B(n_163),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_331),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_331),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_398),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_398),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_359),
.B(n_266),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_398),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_353),
.B(n_149),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_435),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_327),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_327),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_355),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_388),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_357),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_350),
.B(n_354),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_338),
.A2(n_204),
.B(n_202),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_388),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_348),
.B(n_165),
.Y(n_584)
);

AO22x2_ASAP7_75t_L g585 ( 
.A1(n_346),
.A2(n_155),
.B1(n_164),
.B2(n_180),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_363),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_363),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_355),
.B(n_205),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_412),
.B(n_233),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_360),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_360),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_360),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_400),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_388),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_388),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_405),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_388),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_323),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_431),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_405),
.B(n_232),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_434),
.B(n_209),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_323),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_413),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_323),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_436),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_332),
.B(n_183),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_431),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_397),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_339),
.B(n_218),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_432),
.B(n_208),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_339),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_361),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_361),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_343),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_358),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_335),
.B(n_229),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_358),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_358),
.A2(n_210),
.B1(n_177),
.B2(n_178),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_364),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_423),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_364),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_328),
.B(n_222),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_404),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_368),
.B(n_207),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_368),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_349),
.B(n_226),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_420),
.A2(n_216),
.B(n_224),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_349),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_374),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_410),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_342),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_374),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_389),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_389),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_391),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_391),
.B(n_205),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_429),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_399),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_399),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_406),
.B(n_193),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_406),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_411),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_411),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_418),
.Y(n_644)
);

AO21x2_ASAP7_75t_L g645 ( 
.A1(n_418),
.A2(n_132),
.B(n_184),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_397),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_429),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_425),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_425),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_408),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_408),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_414),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_414),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_415),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_322),
.B(n_212),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_352),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_352),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_352),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_352),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_428),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_320),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_320),
.Y(n_662)
);

INVx8_ASAP7_75t_L g663 ( 
.A(n_355),
.Y(n_663)
);

INVxp33_ASAP7_75t_SL g664 ( 
.A(n_366),
.Y(n_664)
);

AOI21x1_ASAP7_75t_L g665 ( 
.A1(n_382),
.A2(n_176),
.B(n_234),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_352),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_428),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_352),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_415),
.B(n_190),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_359),
.B(n_239),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_352),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_318),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_366),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_352),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_319),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_L g676 ( 
.A(n_364),
.B(n_166),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_352),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_352),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_319),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_409),
.B(n_214),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_319),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_322),
.B(n_215),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_319),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_352),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_365),
.A2(n_188),
.B(n_181),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_352),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_319),
.Y(n_687)
);

AND3x2_ASAP7_75t_L g688 ( 
.A(n_415),
.B(n_239),
.C(n_230),
.Y(n_688)
);

CKINVDCx11_ASAP7_75t_R g689 ( 
.A(n_397),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_352),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_409),
.B(n_223),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_322),
.B(n_227),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_352),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_352),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_352),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_352),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_322),
.B(n_228),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_352),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_355),
.B(n_234),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_320),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_352),
.Y(n_701)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_382),
.A2(n_234),
.B(n_184),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_352),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_361),
.B(n_234),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_397),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_352),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_415),
.B(n_230),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_352),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_352),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_352),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_355),
.B(n_184),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_322),
.B(n_184),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_352),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_322),
.B(n_176),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_322),
.B(n_176),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_352),
.Y(n_716)
);

AO21x2_ASAP7_75t_L g717 ( 
.A1(n_365),
.A2(n_44),
.B(n_112),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_428),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_352),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_415),
.B(n_174),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_428),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_415),
.B(n_174),
.C(n_169),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_319),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_352),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_409),
.B(n_5),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_320),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_473),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_536),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_440),
.B(n_33),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_646),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_646),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_473),
.B(n_6),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_608),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_449),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_512),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_580),
.B(n_469),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_491),
.B(n_12),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_449),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_461),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_523),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_526),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_630),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_526),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_461),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_580),
.B(n_61),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_486),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_523),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_558),
.B(n_49),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_527),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_558),
.B(n_63),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_520),
.B(n_36),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_526),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_520),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_527),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_531),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_531),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_486),
.Y(n_757)
);

AND2x6_ASAP7_75t_L g758 ( 
.A(n_440),
.B(n_66),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_539),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_496),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_520),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_539),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_496),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_539),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_491),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_593),
.B(n_15),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_536),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_536),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_525),
.B(n_79),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_536),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_536),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_725),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_512),
.A2(n_87),
.B1(n_97),
.B2(n_95),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_533),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_469),
.B(n_86),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_533),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_608),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_593),
.B(n_596),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_499),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_596),
.B(n_21),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_499),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_508),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_625),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_569),
.B(n_88),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_472),
.B(n_23),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_537),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_569),
.B(n_102),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_439),
.B(n_23),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_439),
.B(n_26),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_508),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_439),
.B(n_27),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_707),
.B(n_720),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_464),
.B(n_465),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_705),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_549),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_640),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_625),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_439),
.B(n_577),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_675),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_675),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_689),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_525),
.B(n_590),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_492),
.B(n_515),
.Y(n_804)
);

OAI221xp5_ASAP7_75t_L g805 ( 
.A1(n_576),
.A2(n_577),
.B1(n_586),
.B2(n_587),
.C(n_592),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_537),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_679),
.Y(n_807)
);

BUFx10_ASAP7_75t_L g808 ( 
.A(n_626),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_705),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_598),
.B(n_602),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_598),
.B(n_602),
.Y(n_811)
);

AND3x2_ASAP7_75t_L g812 ( 
.A(n_530),
.B(n_648),
.C(n_610),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_654),
.B(n_492),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_439),
.B(n_442),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_578),
.B(n_607),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_679),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_549),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_630),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_515),
.B(n_472),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_549),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_681),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_681),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_540),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_549),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_683),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_683),
.Y(n_826)
);

OR2x6_ASAP7_75t_L g827 ( 
.A(n_630),
.B(n_633),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_442),
.B(n_656),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_549),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_687),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_567),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_687),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_463),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_654),
.B(n_467),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_540),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_723),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_723),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_689),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_654),
.B(n_581),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_443),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_443),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_542),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_542),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_543),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_656),
.B(n_657),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_485),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_485),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_513),
.B(n_616),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_604),
.B(n_590),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_489),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_446),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_630),
.B(n_633),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_543),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_591),
.B(n_621),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_489),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_657),
.B(n_658),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_446),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_670),
.B(n_576),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_591),
.B(n_621),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_567),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_630),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_633),
.B(n_648),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_670),
.B(n_605),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_669),
.B(n_612),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_495),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_463),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_673),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_589),
.B(n_603),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_448),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_448),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_450),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_620),
.A2(n_631),
.B1(n_604),
.B2(n_613),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_495),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_450),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_568),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_452),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_452),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_444),
.B(n_447),
.Y(n_878)
);

INVx5_ASAP7_75t_L g879 ( 
.A(n_493),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_457),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_457),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_658),
.B(n_659),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_659),
.B(n_666),
.Y(n_883)
);

INVx4_ASAP7_75t_SL g884 ( 
.A(n_487),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_513),
.B(n_650),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_672),
.Y(n_886)
);

AND3x2_ASAP7_75t_L g887 ( 
.A(n_609),
.B(n_629),
.C(n_628),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_619),
.B(n_607),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_466),
.Y(n_889)
);

CKINVDCx8_ASAP7_75t_R g890 ( 
.A(n_673),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_666),
.B(n_668),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_668),
.B(n_671),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_466),
.Y(n_893)
);

AND2x2_ASAP7_75t_SL g894 ( 
.A(n_633),
.B(n_650),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_470),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_671),
.A2(n_696),
.B1(n_674),
.B2(n_677),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_470),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_477),
.B(n_538),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_633),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_637),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_474),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_619),
.B(n_607),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_474),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_480),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_652),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_622),
.B(n_548),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_585),
.A2(n_453),
.B1(n_695),
.B2(n_710),
.Y(n_907)
);

INVx8_ASAP7_75t_L g908 ( 
.A(n_607),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_674),
.B(n_677),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_SL g910 ( 
.A(n_497),
.B(n_506),
.Y(n_910)
);

NAND3x1_ASAP7_75t_L g911 ( 
.A(n_627),
.B(n_651),
.C(n_649),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_664),
.B(n_611),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_568),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_637),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_619),
.B(n_607),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_637),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_480),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_481),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_451),
.B(n_462),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_623),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_570),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_611),
.B(n_451),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_481),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_482),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_609),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_672),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_585),
.A2(n_453),
.B1(n_695),
.B2(n_698),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_462),
.Y(n_928)
);

AND2x6_ASAP7_75t_L g929 ( 
.A(n_684),
.B(n_686),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_441),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_664),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_482),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_458),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_504),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_484),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_684),
.B(n_686),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_468),
.B(n_661),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_484),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_546),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_504),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_652),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_490),
.Y(n_942)
);

AND2x2_ASAP7_75t_SL g943 ( 
.A(n_653),
.B(n_636),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_468),
.B(n_661),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_662),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_546),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_690),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_662),
.B(n_700),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_700),
.B(n_726),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_585),
.A2(n_453),
.B1(n_693),
.B2(n_713),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_490),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_600),
.B(n_638),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_501),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_504),
.B(n_628),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_690),
.B(n_693),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_653),
.B(n_636),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_694),
.B(n_696),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_642),
.B(n_629),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_458),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_501),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_632),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_632),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_694),
.B(n_698),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_445),
.Y(n_964)
);

AND2x6_ASAP7_75t_L g965 ( 
.A(n_701),
.B(n_703),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_634),
.B(n_635),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_505),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_634),
.B(n_635),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_456),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_726),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_497),
.A2(n_506),
.B1(n_517),
.B2(n_514),
.Y(n_971)
);

BUFx10_ASAP7_75t_L g972 ( 
.A(n_497),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_701),
.B(n_724),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_505),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_599),
.B(n_578),
.Y(n_975)
);

AND2x4_ASAP7_75t_SL g976 ( 
.A(n_599),
.B(n_639),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_639),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_507),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_571),
.B(n_551),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_641),
.B(n_643),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_660),
.B(n_667),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_641),
.B(n_643),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_644),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_718),
.B(n_721),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_507),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_644),
.B(n_647),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_647),
.B(n_494),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_570),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_509),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_509),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_551),
.B(n_552),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_614),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_510),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_510),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_614),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_704),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_724),
.B(n_703),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_546),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_615),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_599),
.B(n_578),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_514),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_552),
.B(n_553),
.Y(n_1002)
);

NOR2x1p5_ASAP7_75t_L g1003 ( 
.A(n_627),
.B(n_722),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_553),
.B(n_547),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_SL g1005 ( 
.A(n_506),
.B(n_493),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_706),
.B(n_709),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_547),
.B(n_550),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_534),
.B(n_588),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_550),
.B(n_555),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_460),
.B(n_557),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_706),
.B(n_709),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_516),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_572),
.Y(n_1013)
);

OAI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_555),
.A2(n_565),
.B1(n_556),
.B2(n_561),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_585),
.A2(n_453),
.B1(n_716),
.B2(n_713),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_516),
.Y(n_1016)
);

OAI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_556),
.A2(n_561),
.B1(n_565),
.B2(n_560),
.Y(n_1017)
);

INVxp67_ASAP7_75t_SL g1018 ( 
.A(n_710),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_562),
.B(n_584),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_475),
.B(n_502),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_559),
.Y(n_1021)
);

INVxp33_ASAP7_75t_L g1022 ( 
.A(n_624),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_716),
.B(n_678),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_680),
.B(n_691),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_517),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_678),
.B(n_708),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_572),
.Y(n_1027)
);

INVx5_ASAP7_75t_L g1028 ( 
.A(n_493),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_459),
.A2(n_545),
.B(n_566),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_519),
.Y(n_1030)
);

XOR2xp5_ASAP7_75t_L g1031 ( 
.A(n_618),
.B(n_503),
.Y(n_1031)
);

NAND2xp33_ASAP7_75t_L g1032 ( 
.A(n_578),
.B(n_493),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_476),
.B(n_479),
.Y(n_1033)
);

AND2x6_ASAP7_75t_L g1034 ( 
.A(n_678),
.B(n_719),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_519),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_615),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_483),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_578),
.B(n_676),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_708),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_617),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_521),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_521),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_488),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_522),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_708),
.B(n_719),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_535),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_582),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_573),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_498),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_573),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_574),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_559),
.Y(n_1052)
);

XNOR2xp5_ASAP7_75t_L g1053 ( 
.A(n_511),
.B(n_528),
.Y(n_1053)
);

OR2x2_ASAP7_75t_SL g1054 ( 
.A(n_688),
.B(n_617),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_529),
.B(n_544),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_500),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_645),
.B(n_704),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_574),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_575),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_575),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_559),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_563),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_719),
.B(n_601),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_563),
.B(n_564),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_563),
.B(n_564),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_564),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_487),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_454),
.B(n_606),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_487),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_655),
.B(n_692),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_554),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_682),
.B(n_697),
.Y(n_1072)
);

AND2x6_ASAP7_75t_L g1073 ( 
.A(n_487),
.B(n_594),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_487),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_594),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_524),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_500),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_SL g1078 ( 
.A(n_704),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_645),
.B(n_704),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_582),
.B(n_541),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_645),
.B(n_582),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_438),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_478),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_597),
.B(n_532),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_685),
.B(n_579),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_438),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_597),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_579),
.B(n_595),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_455),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_532),
.B(n_595),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_717),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_500),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_455),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_717),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_500),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_728),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_792),
.B(n_532),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_898),
.B(n_712),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_906),
.B(n_714),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1007),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_858),
.B(n_471),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_857),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_991),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_863),
.B(n_471),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_920),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_734),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_793),
.B(n_534),
.C(n_588),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_839),
.B(n_715),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_839),
.B(n_471),
.Y(n_1109)
);

AOI22x1_ASAP7_75t_L g1110 ( 
.A1(n_1076),
.A2(n_583),
.B1(n_595),
.B2(n_579),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_864),
.B(n_583),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_738),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_739),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_869),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_819),
.B(n_717),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_864),
.B(n_583),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_977),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1008),
.B(n_518),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_979),
.B(n_518),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_979),
.B(n_518),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_744),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_871),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_746),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_736),
.B(n_518),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_736),
.B(n_663),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_757),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_868),
.B(n_663),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_961),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_947),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_728),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_876),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_745),
.B(n_663),
.Y(n_1132)
);

NOR2x1p5_ASAP7_75t_L g1133 ( 
.A(n_959),
.B(n_665),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_834),
.B(n_1071),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_745),
.B(n_663),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1020),
.A2(n_699),
.B1(n_711),
.B2(n_702),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_894),
.B(n_665),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_947),
.B(n_699),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_881),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1018),
.B(n_1068),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1024),
.A2(n_702),
.B1(n_711),
.B2(n_925),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_893),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_943),
.B(n_956),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_L g1144 ( 
.A(n_879),
.B(n_1028),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1018),
.B(n_1068),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_772),
.A2(n_785),
.B(n_773),
.C(n_1033),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_918),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_799),
.A2(n_1095),
.B1(n_805),
.B2(n_925),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1002),
.A2(n_981),
.B1(n_984),
.B2(n_1004),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_961),
.B(n_983),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_783),
.B(n_798),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_982),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_814),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_986),
.Y(n_1154)
);

INVxp67_ASAP7_75t_L g1155 ( 
.A(n_968),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_962),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_742),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_760),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_905),
.Y(n_1159)
);

AND2x4_ASAP7_75t_SL g1160 ( 
.A(n_827),
.B(n_852),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_1067),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1002),
.B(n_748),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_966),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_763),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_L g1165 ( 
.A(n_753),
.B(n_761),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_938),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1004),
.B(n_778),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_799),
.B(n_1049),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_872),
.B(n_1039),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1009),
.B(n_775),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_983),
.B(n_794),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_742),
.B(n_827),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_SL g1173 ( 
.A1(n_910),
.A2(n_952),
.B1(n_1019),
.B2(n_797),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_872),
.B(n_1039),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1009),
.B(n_814),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_775),
.B(n_784),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_742),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_779),
.Y(n_1178)
);

AND2x6_ASAP7_75t_L g1179 ( 
.A(n_1067),
.B(n_1069),
.Y(n_1179)
);

BUFx4f_ASAP7_75t_L g1180 ( 
.A(n_827),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_966),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_784),
.B(n_787),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_914),
.B(n_916),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_953),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_727),
.B(n_765),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_978),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_914),
.B(n_916),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_727),
.B(n_765),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_748),
.B(n_750),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_989),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_964),
.B(n_969),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_910),
.A2(n_971),
.B1(n_980),
.B2(n_966),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_993),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_994),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_964),
.B(n_969),
.Y(n_1195)
);

NOR2x1p5_ASAP7_75t_L g1196 ( 
.A(n_818),
.B(n_861),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1025),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_781),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_728),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_878),
.B(n_1043),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_787),
.B(n_1067),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1046),
.B(n_804),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_941),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1035),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1044),
.B(n_849),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_777),
.B(n_795),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_840),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_954),
.B(n_958),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_R g1209 ( 
.A(n_866),
.B(n_867),
.Y(n_1209)
);

OAI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_772),
.A2(n_1029),
.B(n_785),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1069),
.B(n_750),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1069),
.B(n_741),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_849),
.B(n_1063),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1063),
.B(n_1029),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_930),
.B(n_1037),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_796),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_841),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_981),
.A2(n_984),
.B1(n_1031),
.B2(n_810),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_809),
.B(n_730),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_930),
.B(n_810),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_899),
.B(n_811),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_SL g1222 ( 
.A(n_890),
.B(n_931),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_899),
.B(n_811),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_782),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_790),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_987),
.A2(n_1057),
.B1(n_1079),
.B2(n_735),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_852),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_851),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_800),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_741),
.B(n_743),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1055),
.B(n_732),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_980),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_735),
.A2(n_919),
.B1(n_937),
.B2(n_803),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_743),
.B(n_752),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_980),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_870),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_805),
.A2(n_1017),
.B(n_1014),
.C(n_766),
.Y(n_1237)
);

BUFx8_ASAP7_75t_L g1238 ( 
.A(n_1078),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_773),
.A2(n_737),
.B(n_780),
.C(n_813),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_852),
.B(n_862),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_801),
.B(n_807),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_816),
.B(n_821),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_862),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_752),
.B(n_759),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_759),
.B(n_762),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_R g1246 ( 
.A(n_733),
.B(n_802),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_822),
.B(n_825),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_826),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_830),
.Y(n_1249)
);

NOR3xp33_ASAP7_75t_L g1250 ( 
.A(n_912),
.B(n_1083),
.C(n_922),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1022),
.B(n_808),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_832),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_731),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_862),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_836),
.B(n_837),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_762),
.B(n_764),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_919),
.B(n_937),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_808),
.B(n_797),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1060),
.B(n_828),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_874),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1060),
.B(n_828),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_796),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_845),
.B(n_882),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_SL g1264 ( 
.A(n_833),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_907),
.A2(n_950),
.B1(n_1015),
.B2(n_927),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_764),
.B(n_1017),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_877),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_812),
.B(n_788),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1053),
.A2(n_971),
.B1(n_1003),
.B2(n_1005),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_880),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_900),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_788),
.A2(n_789),
.B1(n_791),
.B2(n_769),
.Y(n_1272)
);

NAND2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1077),
.B(n_1092),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1014),
.A2(n_789),
.B(n_791),
.C(n_751),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1083),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_883),
.B(n_891),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_892),
.B(n_909),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_892),
.B(n_909),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_936),
.B(n_955),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_L g1280 ( 
.A(n_908),
.B(n_879),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_889),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_895),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_812),
.B(n_887),
.C(n_944),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_936),
.B(n_955),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1005),
.A2(n_1072),
.B1(n_1070),
.B2(n_948),
.Y(n_1285)
);

BUFx8_ASAP7_75t_L g1286 ( 
.A(n_1078),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_897),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_928),
.B(n_945),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_928),
.B(n_945),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_901),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_939),
.Y(n_1291)
);

AO221x1_ASAP7_75t_L g1292 ( 
.A1(n_1094),
.A2(n_771),
.B1(n_995),
.B2(n_1040),
.C(n_992),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_963),
.B(n_973),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_903),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_904),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_928),
.B(n_945),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_917),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_923),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_924),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_963),
.B(n_973),
.Y(n_1300)
);

OAI22x1_ASAP7_75t_R g1301 ( 
.A1(n_838),
.A2(n_933),
.B1(n_833),
.B2(n_972),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_970),
.B(n_879),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_932),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_935),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_976),
.B(n_934),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_970),
.B(n_879),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_997),
.B(n_1006),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_942),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_970),
.B(n_1028),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_951),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_960),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_911),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_887),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_967),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_997),
.B(n_1006),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_L g1316 ( 
.A1(n_1085),
.A2(n_1094),
.B(n_888),
.C(n_902),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1023),
.B(n_856),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1047),
.A2(n_949),
.B1(n_1081),
.B2(n_1050),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_974),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_985),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_972),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_940),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_990),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1032),
.A2(n_915),
.B(n_1056),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1010),
.A2(n_753),
.B1(n_761),
.B2(n_996),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1001),
.Y(n_1326)
);

AO22x2_ASAP7_75t_L g1327 ( 
.A1(n_1047),
.A2(n_1091),
.B1(n_884),
.B2(n_896),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_740),
.A2(n_853),
.B1(n_747),
.B2(n_749),
.Y(n_1328)
);

NAND2xp33_ASAP7_75t_L g1329 ( 
.A(n_908),
.B(n_1028),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_847),
.B(n_850),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1023),
.B(n_856),
.Y(n_1331)
);

INVxp33_ASAP7_75t_L g1332 ( 
.A(n_847),
.Y(n_1332)
);

BUFx5_ASAP7_75t_L g1333 ( 
.A(n_1034),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_856),
.B(n_929),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1054),
.B(n_1010),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1012),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1010),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_856),
.B(n_929),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1016),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_929),
.B(n_957),
.Y(n_1340)
);

OAI221xp5_ASAP7_75t_L g1341 ( 
.A1(n_907),
.A2(n_927),
.B1(n_950),
.B2(n_1015),
.C(n_859),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_929),
.B(n_957),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_847),
.B(n_850),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_854),
.A2(n_1080),
.B1(n_1041),
.B2(n_1030),
.C(n_1042),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_957),
.B(n_965),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1028),
.B(n_1056),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_957),
.B(n_965),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_965),
.B(n_1011),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_754),
.B(n_755),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_965),
.B(n_1011),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_756),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1056),
.B(n_992),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_774),
.A2(n_844),
.B1(n_843),
.B2(n_823),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1056),
.B(n_992),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_776),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_939),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1011),
.B(n_1026),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_786),
.A2(n_842),
.B1(n_835),
.B2(n_806),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1077),
.B(n_1092),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1011),
.B(n_1026),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_850),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_855),
.B(n_926),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1051),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1045),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_855),
.B(n_926),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1045),
.B(n_1034),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_855),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1065),
.A2(n_846),
.B1(n_926),
.B2(n_886),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_995),
.B(n_1036),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_865),
.B(n_886),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_995),
.B(n_1036),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1034),
.B(n_1065),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1058),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1066),
.A2(n_886),
.B1(n_873),
.B2(n_865),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1074),
.A2(n_815),
.B1(n_1090),
.B2(n_896),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1034),
.B(n_908),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_865),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_873),
.A2(n_729),
.B1(n_758),
.B2(n_1036),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_999),
.B(n_1040),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1061),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_831),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_873),
.Y(n_1382)
);

NAND2xp33_ASAP7_75t_L g1383 ( 
.A(n_815),
.B(n_729),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1062),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_831),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_846),
.B(n_988),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_860),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_875),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_875),
.B(n_1013),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_913),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_913),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_921),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1080),
.B(n_999),
.C(n_1040),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_884),
.B(n_771),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1090),
.C(n_1084),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1059),
.B(n_1048),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_999),
.B(n_884),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_921),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1013),
.B(n_1027),
.Y(n_1399)
);

INVx8_ASAP7_75t_L g1400 ( 
.A(n_1073),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_796),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1027),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1048),
.B(n_1059),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1059),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_946),
.B(n_1021),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_946),
.B(n_1021),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1084),
.A2(n_1000),
.B1(n_975),
.B2(n_729),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1075),
.B(n_1087),
.Y(n_1408)
);

NAND2x1_ASAP7_75t_L g1409 ( 
.A(n_767),
.B(n_829),
.Y(n_1409)
);

CKINVDCx16_ASAP7_75t_R g1410 ( 
.A(n_1075),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_817),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1064),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1064),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_998),
.A2(n_1052),
.B1(n_829),
.B2(n_767),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_729),
.A2(n_758),
.B1(n_1075),
.B2(n_1087),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_817),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_817),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1087),
.B(n_820),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1082),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_820),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_820),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_998),
.B(n_1052),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_768),
.B(n_770),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_768),
.Y(n_1424)
);

NAND2xp33_ASAP7_75t_L g1425 ( 
.A(n_758),
.B(n_1073),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1086),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_770),
.B(n_824),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_824),
.B(n_1038),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1088),
.B(n_1073),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_L g1430 ( 
.A(n_758),
.B(n_1073),
.Y(n_1430)
);

NOR3xp33_ASAP7_75t_L g1431 ( 
.A(n_792),
.B(n_906),
.C(n_346),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1007),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_792),
.B(n_906),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_792),
.A2(n_906),
.B1(n_793),
.B2(n_898),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_858),
.B(n_472),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1007),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_858),
.B(n_472),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_920),
.Y(n_1438)
);

NOR3xp33_ASAP7_75t_L g1439 ( 
.A(n_792),
.B(n_906),
.C(n_346),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_920),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_862),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_857),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_792),
.B(n_898),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_906),
.B(n_512),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_792),
.B(n_898),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_858),
.B(n_472),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1007),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1007),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_792),
.B(n_898),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_857),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_906),
.B(n_512),
.Y(n_1451)
);

AND2x6_ASAP7_75t_L g1452 ( 
.A(n_1067),
.B(n_1069),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_857),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_857),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_857),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_858),
.B(n_472),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_792),
.B(n_906),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_792),
.B(n_906),
.Y(n_1458)
);

NAND2xp33_ASAP7_75t_L g1459 ( 
.A(n_898),
.B(n_607),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_968),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_857),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_792),
.B(n_898),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_742),
.B(n_827),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_857),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1007),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_792),
.B(n_898),
.Y(n_1466)
);

AO221x1_ASAP7_75t_L g1467 ( 
.A1(n_735),
.A2(n_585),
.B1(n_344),
.B2(n_351),
.C(n_872),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_SL g1468 ( 
.A(n_833),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_728),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1007),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1007),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1007),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_792),
.B(n_898),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_792),
.B(n_898),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_SL g1475 ( 
.A(n_833),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_792),
.A2(n_906),
.B(n_793),
.C(n_720),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_792),
.B(n_898),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_792),
.B(n_906),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_792),
.B(n_898),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_742),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_792),
.B(n_898),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_792),
.B(n_898),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1007),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_857),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_906),
.B(n_512),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1032),
.A2(n_578),
.B(n_500),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_792),
.B(n_898),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_858),
.B(n_472),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_906),
.B(n_512),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_920),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_857),
.Y(n_1491)
);

NOR2xp67_ASAP7_75t_L g1492 ( 
.A(n_866),
.B(n_364),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1007),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_906),
.B(n_512),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_792),
.B(n_898),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_947),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_792),
.B(n_898),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_906),
.B(n_512),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_858),
.B(n_472),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1007),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_857),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_857),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_728),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_792),
.B(n_898),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_792),
.A2(n_906),
.B1(n_707),
.B2(n_720),
.C(n_793),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1007),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_792),
.B(n_898),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_792),
.B(n_898),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_SL g1509 ( 
.A(n_833),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_906),
.B(n_512),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1007),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_906),
.B(n_512),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_792),
.B(n_906),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_857),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_792),
.B(n_898),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_906),
.B(n_512),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1007),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_858),
.B(n_472),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_866),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1007),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_792),
.B(n_898),
.Y(n_1521)
);

NAND2xp33_ASAP7_75t_L g1522 ( 
.A(n_898),
.B(n_607),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_792),
.B(n_898),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_792),
.B(n_898),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_792),
.A2(n_906),
.B1(n_707),
.B2(n_720),
.C(n_793),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_920),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_792),
.B(n_898),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_792),
.B(n_898),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_792),
.A2(n_906),
.B1(n_793),
.B2(n_898),
.Y(n_1529)
);

NAND2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1095),
.B(n_1067),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_792),
.B(n_898),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1007),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_857),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_906),
.B(n_512),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_792),
.A2(n_793),
.B1(n_906),
.B2(n_898),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1007),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_906),
.B(n_512),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_906),
.B(n_512),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1007),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_906),
.B(n_512),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_857),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_968),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_792),
.B(n_906),
.C(n_720),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1007),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1007),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_939),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_857),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_857),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_857),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_792),
.B(n_906),
.C(n_346),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_792),
.B(n_906),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1007),
.Y(n_1552)
);

NOR2xp67_ASAP7_75t_L g1553 ( 
.A(n_866),
.B(n_364),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_792),
.B(n_898),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_968),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_792),
.A2(n_793),
.B1(n_906),
.B2(n_898),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_792),
.A2(n_906),
.B1(n_707),
.B2(n_720),
.C(n_793),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_906),
.B(n_512),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_728),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_L g1560 ( 
.A(n_792),
.B(n_906),
.C(n_346),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_857),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1007),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_848),
.B(n_885),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_906),
.B(n_512),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_857),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_848),
.B(n_885),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_857),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_848),
.B(n_885),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_792),
.B(n_898),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_906),
.B(n_512),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_792),
.B(n_906),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_906),
.A2(n_792),
.B1(n_848),
.B2(n_344),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_792),
.A2(n_906),
.B1(n_793),
.B2(n_898),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_792),
.A2(n_906),
.B1(n_793),
.B2(n_898),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_862),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1007),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_792),
.B(n_898),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_792),
.B(n_898),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_968),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_792),
.B(n_898),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_857),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1032),
.A2(n_578),
.B(n_500),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_792),
.B(n_898),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1007),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_792),
.B(n_898),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_792),
.B(n_898),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1007),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_857),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_792),
.A2(n_906),
.B1(n_793),
.B2(n_898),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_906),
.B(n_512),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_906),
.B(n_512),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1007),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_792),
.B(n_906),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_858),
.B(n_472),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1007),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1007),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_792),
.B(n_906),
.C(n_720),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_L g1598 ( 
.A(n_792),
.B(n_906),
.C(n_346),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1007),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_920),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_857),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_742),
.B(n_827),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_858),
.B(n_472),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_792),
.B(n_906),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_968),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_906),
.B(n_512),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_792),
.B(n_898),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_858),
.B(n_472),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_792),
.B(n_898),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1007),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_792),
.B(n_906),
.Y(n_1611)
);

NOR2x1p5_ASAP7_75t_L g1612 ( 
.A(n_959),
.B(n_458),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_908),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_857),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_792),
.B(n_898),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_857),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_792),
.B(n_898),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_920),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_906),
.A2(n_792),
.B1(n_848),
.B2(n_344),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_792),
.B(n_906),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1426),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1419),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1400),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1419),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1433),
.B(n_1457),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1209),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1433),
.B(n_1457),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1364),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1444),
.B(n_1451),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1458),
.B(n_1478),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1364),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1189),
.B(n_1162),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1476),
.A2(n_1525),
.B(n_1505),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1259),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1478),
.A2(n_1513),
.B1(n_1571),
.B2(n_1551),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_R g1636 ( 
.A(n_1519),
.B(n_1530),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1619),
.B(n_1572),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1434),
.B(n_1529),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1189),
.B(n_1162),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1400),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1458),
.B(n_1513),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_R g1642 ( 
.A(n_1530),
.B(n_1410),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1207),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1159),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1180),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1180),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1551),
.B(n_1571),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1261),
.Y(n_1648)
);

O2A1O1Ixp5_ASAP7_75t_L g1649 ( 
.A1(n_1543),
.A2(n_1597),
.B(n_1604),
.C(n_1593),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1207),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1217),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1400),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1160),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1573),
.B(n_1574),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1217),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1593),
.A2(n_1611),
.B1(n_1620),
.B2(n_1604),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1228),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1129),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1611),
.B(n_1620),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1333),
.Y(n_1660)
);

AO22x1_ASAP7_75t_L g1661 ( 
.A1(n_1431),
.A2(n_1550),
.B1(n_1560),
.B2(n_1439),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1228),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1179),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1160),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1189),
.B(n_1162),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1236),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1557),
.B(n_1589),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1240),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1236),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1333),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1267),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1146),
.A2(n_1210),
.B1(n_1556),
.B2(n_1535),
.C(n_1265),
.Y(n_1673)
);

BUFx8_ASAP7_75t_L g1674 ( 
.A(n_1264),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1240),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1146),
.A2(n_1462),
.B1(n_1466),
.B2(n_1449),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1598),
.A2(n_1474),
.B1(n_1477),
.B2(n_1473),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1208),
.B(n_1444),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1128),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1479),
.B(n_1481),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1282),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1482),
.B(n_1487),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1134),
.B(n_1173),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1294),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1495),
.B(n_1497),
.Y(n_1686)
);

XOR2xp5_ASAP7_75t_L g1687 ( 
.A(n_1206),
.B(n_1335),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1504),
.A2(n_1508),
.B1(n_1515),
.B2(n_1507),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1333),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1239),
.A2(n_1107),
.B(n_1099),
.C(n_1521),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1523),
.B(n_1524),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1239),
.A2(n_1099),
.B(n_1528),
.C(n_1527),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1531),
.B(n_1554),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1294),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1569),
.B(n_1577),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1297),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1451),
.A2(n_1485),
.B1(n_1494),
.B2(n_1489),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1209),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1246),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1578),
.B(n_1580),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1221),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1583),
.B(n_1585),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1586),
.B(n_1607),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1609),
.B(n_1615),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1617),
.B(n_1168),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1156),
.Y(n_1706)
);

O2A1O1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1485),
.A2(n_1494),
.B(n_1498),
.C(n_1489),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1240),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1297),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1303),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1171),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1498),
.B(n_1510),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1510),
.B(n_1512),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1512),
.B(n_1516),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1516),
.B(n_1534),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1534),
.B(n_1537),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1537),
.A2(n_1540),
.B1(n_1558),
.B2(n_1538),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1538),
.A2(n_1558),
.B1(n_1564),
.B2(n_1540),
.Y(n_1718)
);

INVxp67_ASAP7_75t_SL g1719 ( 
.A(n_1496),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1564),
.A2(n_1590),
.B1(n_1591),
.B2(n_1570),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1570),
.B(n_1590),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1120),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1563),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1591),
.A2(n_1606),
.B1(n_1467),
.B2(n_1218),
.Y(n_1724)
);

OAI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1155),
.A2(n_1542),
.B1(n_1579),
.B2(n_1555),
.C(n_1460),
.Y(n_1725)
);

AO22x1_ASAP7_75t_L g1726 ( 
.A1(n_1312),
.A2(n_1268),
.B1(n_1250),
.B2(n_1313),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1606),
.B(n_1435),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1333),
.Y(n_1728)
);

BUFx12f_ASAP7_75t_SL g1729 ( 
.A(n_1172),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1153),
.B(n_1169),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1303),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1304),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1566),
.B(n_1568),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1174),
.B(n_1175),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1605),
.B(n_1150),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1304),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1308),
.Y(n_1737)
);

AND3x1_ASAP7_75t_L g1738 ( 
.A(n_1269),
.B(n_1251),
.C(n_1268),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1437),
.B(n_1446),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1161),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1150),
.B(n_1213),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1308),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1203),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1221),
.B(n_1223),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1492),
.B(n_1553),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1183),
.B(n_1187),
.Y(n_1746)
);

NAND2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1118),
.B(n_1346),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1456),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1314),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1226),
.A2(n_1251),
.B1(n_1337),
.B2(n_1258),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1161),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1314),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1320),
.Y(n_1753)
);

OR2x2_ASAP7_75t_SL g1754 ( 
.A(n_1283),
.B(n_1231),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1149),
.B(n_1488),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1183),
.B(n_1187),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1119),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1143),
.B(n_1214),
.Y(n_1758)
);

BUFx12f_ASAP7_75t_L g1759 ( 
.A(n_1238),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1143),
.B(n_1263),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1325),
.B(n_1258),
.C(n_1192),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1320),
.Y(n_1762)
);

AO22x1_ASAP7_75t_L g1763 ( 
.A1(n_1200),
.A2(n_1109),
.B1(n_1127),
.B2(n_1148),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1367),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1323),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1104),
.B(n_1097),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1341),
.A2(n_1415),
.B1(n_1233),
.B2(n_1378),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1499),
.A2(n_1594),
.B1(n_1603),
.B2(n_1518),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1161),
.Y(n_1770)
);

OAI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1608),
.A2(n_1195),
.B(n_1191),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1323),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1326),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1246),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1161),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1326),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1100),
.B(n_1432),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1339),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1339),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1394),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1275),
.A2(n_1103),
.B1(n_1109),
.B2(n_1215),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1102),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1284),
.B(n_1293),
.Y(n_1784)
);

BUFx4f_ASAP7_75t_L g1785 ( 
.A(n_1172),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1393),
.B(n_1459),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1105),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1300),
.B(n_1307),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1152),
.B(n_1154),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1221),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1441),
.A2(n_1575),
.B1(n_1243),
.B2(n_1223),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1102),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1223),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1114),
.Y(n_1794)
);

NOR2x2_ASAP7_75t_L g1795 ( 
.A(n_1172),
.B(n_1463),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1438),
.B(n_1440),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1114),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1315),
.B(n_1108),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1122),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1522),
.A2(n_1582),
.B(n_1486),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1490),
.B(n_1526),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1463),
.B(n_1602),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1122),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1101),
.A2(n_1436),
.B1(n_1448),
.B2(n_1447),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1292),
.Y(n_1805)
);

NOR2x2_ASAP7_75t_L g1806 ( 
.A(n_1463),
.B(n_1602),
.Y(n_1806)
);

OR2x6_ASAP7_75t_SL g1807 ( 
.A(n_1321),
.B(n_1420),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1465),
.A2(n_1470),
.B1(n_1472),
.B2(n_1471),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1483),
.A2(n_1493),
.B1(n_1506),
.B2(n_1500),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1108),
.B(n_1098),
.Y(n_1810)
);

INVx5_ASAP7_75t_L g1811 ( 
.A(n_1179),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1167),
.B(n_1111),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1253),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1257),
.B(n_1219),
.C(n_1254),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1116),
.B(n_1511),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1600),
.B(n_1618),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1131),
.B(n_1139),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1253),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1517),
.B(n_1520),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1131),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_R g1821 ( 
.A(n_1222),
.B(n_1157),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1602),
.B(n_1227),
.Y(n_1822)
);

OR2x6_ASAP7_75t_L g1823 ( 
.A(n_1237),
.B(n_1211),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1139),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1394),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1117),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1142),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1227),
.B(n_1211),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1142),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1532),
.B(n_1536),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1118),
.B(n_1346),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1185),
.B(n_1188),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1539),
.B(n_1544),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1202),
.B(n_1545),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1147),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1552),
.A2(n_1576),
.B1(n_1584),
.B2(n_1562),
.Y(n_1836)
);

AND2x6_ASAP7_75t_L g1837 ( 
.A(n_1291),
.B(n_1356),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1147),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1587),
.B(n_1592),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1166),
.Y(n_1840)
);

OR2x4_ASAP7_75t_L g1841 ( 
.A(n_1330),
.B(n_1343),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1333),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1595),
.B(n_1596),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1184),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1599),
.B(n_1610),
.Y(n_1845)
);

BUFx4f_ASAP7_75t_L g1846 ( 
.A(n_1424),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1327),
.A2(n_1395),
.B1(n_1242),
.B2(n_1247),
.Y(n_1847)
);

INVx5_ASAP7_75t_L g1848 ( 
.A(n_1179),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1238),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1333),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1220),
.B(n_1205),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1186),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1186),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1332),
.B(n_1232),
.Y(n_1854)
);

INVx3_ASAP7_75t_L g1855 ( 
.A(n_1333),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1190),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1291),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1179),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1613),
.B(n_1394),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1285),
.B(n_1163),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1241),
.B(n_1255),
.Y(n_1861)
);

NOR3xp33_ASAP7_75t_SL g1862 ( 
.A(n_1330),
.B(n_1362),
.C(n_1343),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1106),
.B(n_1112),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1190),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1238),
.A2(n_1286),
.B1(n_1327),
.B2(n_1383),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1235),
.A2(n_1272),
.B1(n_1181),
.B2(n_1322),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1170),
.A2(n_1115),
.B1(n_1121),
.B2(n_1113),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1193),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1194),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1194),
.B(n_1197),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1170),
.A2(n_1123),
.B1(n_1158),
.B2(n_1126),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1197),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1204),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1164),
.B(n_1178),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1271),
.B(n_1367),
.Y(n_1875)
);

INVx4_ASAP7_75t_L g1876 ( 
.A(n_1179),
.Y(n_1876)
);

NAND2xp33_ASAP7_75t_L g1877 ( 
.A(n_1424),
.B(n_1165),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1198),
.B(n_1224),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1332),
.B(n_1424),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1424),
.B(n_1305),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1452),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1266),
.A2(n_1252),
.B1(n_1249),
.B2(n_1248),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1204),
.Y(n_1883)
);

INVx4_ASAP7_75t_L g1884 ( 
.A(n_1452),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1442),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1411),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1225),
.B(n_1229),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1442),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1356),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1260),
.B(n_1270),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1382),
.B(n_1361),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_SL g1892 ( 
.A(n_1274),
.B(n_1141),
.C(n_1125),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1450),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1452),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1450),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1281),
.B(n_1287),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1613),
.B(n_1372),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1452),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1452),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1377),
.B(n_1151),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1362),
.B(n_1365),
.Y(n_1901)
);

INVx4_ASAP7_75t_L g1902 ( 
.A(n_1096),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1368),
.B(n_1365),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1290),
.B(n_1295),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1351),
.A2(n_1355),
.B1(n_1373),
.B2(n_1363),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1411),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1370),
.B(n_1157),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1298),
.A2(n_1319),
.B1(n_1336),
.B2(n_1311),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1357),
.B(n_1360),
.Y(n_1909)
);

NAND2x1p5_ASAP7_75t_L g1910 ( 
.A(n_1266),
.B(n_1302),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1096),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1454),
.B(n_1455),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_R g1914 ( 
.A(n_1177),
.B(n_1480),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1455),
.B(n_1461),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1464),
.B(n_1484),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1230),
.B(n_1234),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1546),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_1286),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1484),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_R g1923 ( 
.A(n_1480),
.B(n_1264),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1491),
.B(n_1501),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1491),
.B(n_1501),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1502),
.B(n_1514),
.Y(n_1926)
);

A2O1A1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1316),
.A2(n_1395),
.B(n_1407),
.C(n_1124),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1502),
.B(n_1514),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1546),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1359),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1096),
.Y(n_1931)
);

OR2x4_ASAP7_75t_L g1932 ( 
.A(n_1423),
.B(n_1396),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1533),
.B(n_1541),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1533),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1468),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1541),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1547),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1286),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1359),
.Y(n_1939)
);

AND2x6_ASAP7_75t_L g1940 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1940)
);

INVxp67_ASAP7_75t_L g1941 ( 
.A(n_1468),
.Y(n_1941)
);

NAND3xp33_ASAP7_75t_L g1942 ( 
.A(n_1318),
.B(n_1344),
.C(n_1328),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1096),
.Y(n_1943)
);

NOR2x1_ASAP7_75t_L g1944 ( 
.A(n_1144),
.B(n_1280),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1547),
.B(n_1548),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1374),
.B(n_1386),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1548),
.Y(n_1947)
);

AND2x6_ASAP7_75t_SL g1948 ( 
.A(n_1301),
.B(n_1396),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1404),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1327),
.A2(n_1138),
.B1(n_1136),
.B2(n_1406),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1549),
.B(n_1561),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1549),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1561),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1349),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1565),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1565),
.A2(n_1616),
.B1(n_1614),
.B2(n_1601),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1130),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1567),
.B(n_1581),
.Y(n_1958)
);

INVx5_ASAP7_75t_L g1959 ( 
.A(n_1130),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1567),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1475),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1581),
.A2(n_1616),
.B1(n_1614),
.B2(n_1601),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1588),
.B(n_1317),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1588),
.B(n_1331),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1381),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1381),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1390),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1475),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1144),
.A2(n_1132),
.B(n_1135),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1130),
.Y(n_1970)
);

BUFx2_ASAP7_75t_L g1971 ( 
.A(n_1130),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1390),
.B(n_1392),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1406),
.A2(n_1375),
.B1(n_1405),
.B2(n_1422),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1399),
.B(n_1392),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1398),
.B(n_1403),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1230),
.B(n_1234),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1509),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1398),
.Y(n_1978)
);

OAI21xp33_ASAP7_75t_L g1979 ( 
.A1(n_1380),
.A2(n_1384),
.B(n_1353),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1199),
.B(n_1216),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1288),
.A2(n_1296),
.B1(n_1289),
.B2(n_1244),
.Y(n_1981)
);

NOR2xp67_ASAP7_75t_L g1982 ( 
.A(n_1376),
.B(n_1412),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1199),
.B(n_1401),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1385),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1389),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1199),
.B(n_1469),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1340),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1199),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1366),
.B(n_1358),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1509),
.Y(n_1991)
);

A2O1A1Ixp33_ASAP7_75t_SL g1992 ( 
.A1(n_1423),
.A2(n_1425),
.B(n_1430),
.C(n_1324),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1342),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1345),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1347),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1196),
.A2(n_1288),
.B1(n_1296),
.B2(n_1289),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1413),
.B(n_1402),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1391),
.B(n_1369),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1348),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1350),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1369),
.B(n_1379),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1371),
.B(n_1379),
.Y(n_2002)
);

NOR2x2_ASAP7_75t_L g2003 ( 
.A(n_1612),
.B(n_1421),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1216),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1244),
.B(n_1256),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1371),
.B(n_1408),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1245),
.Y(n_2007)
);

INVx6_ASAP7_75t_L g2008 ( 
.A(n_1216),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1216),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1408),
.B(n_1418),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_1262),
.Y(n_2012)
);

CKINVDCx20_ASAP7_75t_R g2013 ( 
.A(n_1262),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1212),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1201),
.A2(n_1429),
.B1(n_1212),
.B2(n_1137),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1418),
.B(n_1201),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1262),
.B(n_1559),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_R g2018 ( 
.A(n_1329),
.B(n_1559),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1262),
.B(n_1559),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1429),
.B(n_1397),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1401),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1397),
.B(n_1559),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1401),
.B(n_1503),
.Y(n_2023)
);

INVxp33_ASAP7_75t_L g2024 ( 
.A(n_1401),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1110),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1132),
.A2(n_1135),
.B(n_1137),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1469),
.Y(n_2027)
);

NOR2xp67_ASAP7_75t_L g2028 ( 
.A(n_1416),
.B(n_1417),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1469),
.B(n_1503),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1469),
.B(n_1503),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1428),
.B(n_1427),
.Y(n_2031)
);

NOR2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1409),
.B(n_1417),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1428),
.B(n_1302),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1503),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1352),
.Y(n_2035)
);

NAND2xp33_ASAP7_75t_L g2036 ( 
.A(n_1273),
.B(n_1306),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1416),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1306),
.B(n_1309),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1133),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1309),
.A2(n_1352),
.B1(n_1354),
.B2(n_1414),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1354),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1273),
.B(n_858),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1426),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2044)
);

BUFx3_ASAP7_75t_L g2045 ( 
.A(n_1180),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1159),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1209),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_1159),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1159),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_R g2052 ( 
.A(n_1519),
.B(n_397),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1180),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1209),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1400),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1426),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1400),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1426),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1426),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1208),
.B(n_858),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1419),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1419),
.Y(n_2067)
);

INVxp67_ASAP7_75t_L g2068 ( 
.A(n_1159),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1180),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1159),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1209),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1419),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_1159),
.Y(n_2075)
);

INVxp67_ASAP7_75t_L g2076 ( 
.A(n_1159),
.Y(n_2076)
);

CKINVDCx20_ASAP7_75t_R g2077 ( 
.A(n_1209),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_1161),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1400),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2081)
);

NOR2x1p5_ASAP7_75t_L g2082 ( 
.A(n_1335),
.B(n_458),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2083)
);

NAND2x1p5_ASAP7_75t_L g2084 ( 
.A(n_1180),
.B(n_1067),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1426),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1419),
.Y(n_2089)
);

NOR3xp33_ASAP7_75t_SL g2090 ( 
.A(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1400),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_SL g2093 ( 
.A1(n_1433),
.A2(n_1457),
.B1(n_1478),
.B2(n_1458),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1419),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2095)
);

INVx5_ASAP7_75t_L g2096 ( 
.A(n_1179),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2100)
);

BUFx3_ASAP7_75t_L g2101 ( 
.A(n_1180),
.Y(n_2101)
);

INVx5_ASAP7_75t_L g2102 ( 
.A(n_1179),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1400),
.Y(n_2103)
);

AOI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_1476),
.A2(n_792),
.B(n_1505),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1426),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1426),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1426),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1419),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1419),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_1400),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1161),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1400),
.Y(n_2116)
);

OAI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1159),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1426),
.Y(n_2122)
);

BUFx4f_ASAP7_75t_L g2123 ( 
.A(n_1400),
.Y(n_2123)
);

XNOR2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1519),
.B(n_342),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2126)
);

INVx3_ASAP7_75t_L g2127 ( 
.A(n_1400),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1426),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1159),
.Y(n_2130)
);

INVxp67_ASAP7_75t_L g2131 ( 
.A(n_1159),
.Y(n_2131)
);

BUFx8_ASAP7_75t_L g2132 ( 
.A(n_1264),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1419),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1419),
.Y(n_2135)
);

NOR3xp33_ASAP7_75t_SL g2136 ( 
.A(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1180),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2138)
);

BUFx4f_ASAP7_75t_L g2139 ( 
.A(n_1400),
.Y(n_2139)
);

BUFx8_ASAP7_75t_L g2140 ( 
.A(n_1264),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2141)
);

O2A1O1Ixp33_ASAP7_75t_L g2142 ( 
.A1(n_1505),
.A2(n_1525),
.B(n_1557),
.C(n_1476),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1208),
.B(n_858),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_1128),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1426),
.Y(n_2151)
);

OR2x6_ASAP7_75t_L g2152 ( 
.A(n_1240),
.B(n_1189),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1209),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1419),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_1400),
.Y(n_2155)
);

INVx5_ASAP7_75t_L g2156 ( 
.A(n_1179),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1426),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1209),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1426),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2162)
);

NAND2xp33_ASAP7_75t_L g2163 ( 
.A(n_1146),
.B(n_1431),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1419),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1419),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1419),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1426),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1426),
.Y(n_2170)
);

NOR3xp33_ASAP7_75t_L g2171 ( 
.A(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_1444),
.B(n_1451),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1008),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1419),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_1159),
.Y(n_2176)
);

O2A1O1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_1505),
.A2(n_1525),
.B(n_1557),
.C(n_1476),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1180),
.Y(n_2178)
);

OR2x6_ASAP7_75t_L g2179 ( 
.A(n_1240),
.B(n_1189),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1419),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1209),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1419),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1426),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1208),
.B(n_858),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1208),
.B(n_858),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1426),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1400),
.Y(n_2194)
);

OAI221xp5_ASAP7_75t_L g2195 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1513),
.B2(n_1478),
.C(n_1457),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1426),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1426),
.Y(n_2197)
);

NOR2x2_ASAP7_75t_L g2198 ( 
.A(n_1240),
.B(n_650),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1400),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2200)
);

A2O1A1Ixp33_ASAP7_75t_L g2201 ( 
.A1(n_1433),
.A2(n_1457),
.B(n_1478),
.C(n_1458),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_1159),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1426),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1400),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_1159),
.Y(n_2206)
);

AND2x6_ASAP7_75t_SL g2207 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_SL g2208 ( 
.A(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_SL g2209 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1426),
.Y(n_2213)
);

AOI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1426),
.Y(n_2215)
);

NAND2x1p5_ASAP7_75t_L g2216 ( 
.A(n_1180),
.B(n_1067),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2217)
);

INVx3_ASAP7_75t_L g2218 ( 
.A(n_1400),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1400),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1209),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1426),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1426),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2225)
);

INVx2_ASAP7_75t_SL g2226 ( 
.A(n_1367),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1419),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1419),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1208),
.B(n_858),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1180),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1426),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1419),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2237)
);

NOR3xp33_ASAP7_75t_SL g2238 ( 
.A(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1426),
.Y(n_2239)
);

INVx5_ASAP7_75t_L g2240 ( 
.A(n_1179),
.Y(n_2240)
);

NAND2x1p5_ASAP7_75t_L g2241 ( 
.A(n_1180),
.B(n_1067),
.Y(n_2241)
);

NAND2x1p5_ASAP7_75t_L g2242 ( 
.A(n_1180),
.B(n_1067),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_1180),
.Y(n_2244)
);

INVx5_ASAP7_75t_L g2245 ( 
.A(n_1179),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_1161),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_1159),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2248)
);

INVx2_ASAP7_75t_SL g2249 ( 
.A(n_1161),
.Y(n_2249)
);

AND2x6_ASAP7_75t_SL g2250 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1426),
.Y(n_2251)
);

BUFx12f_ASAP7_75t_L g2252 ( 
.A(n_1238),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1208),
.B(n_858),
.Y(n_2254)
);

INVx5_ASAP7_75t_L g2255 ( 
.A(n_1179),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2256)
);

INVx4_ASAP7_75t_SL g2257 ( 
.A(n_1179),
.Y(n_2257)
);

BUFx3_ASAP7_75t_L g2258 ( 
.A(n_1180),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_SL g2259 ( 
.A(n_1476),
.B(n_1525),
.C(n_1505),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1426),
.Y(n_2260)
);

INVx2_ASAP7_75t_SL g2261 ( 
.A(n_1367),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1419),
.Y(n_2262)
);

BUFx4f_ASAP7_75t_L g2263 ( 
.A(n_1400),
.Y(n_2263)
);

OR2x6_ASAP7_75t_L g2264 ( 
.A(n_1240),
.B(n_1189),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1426),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1426),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1208),
.B(n_858),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2269)
);

INVx1_ASAP7_75t_SL g2270 ( 
.A(n_1128),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_1128),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_1209),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1426),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1426),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1426),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1426),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2281)
);

OAI21xp33_ASAP7_75t_SL g2282 ( 
.A1(n_1140),
.A2(n_1008),
.B(n_1145),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1426),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1419),
.Y(n_2284)
);

OAI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_1433),
.A2(n_1457),
.B1(n_1478),
.B2(n_1458),
.Y(n_2285)
);

INVx3_ASAP7_75t_L g2286 ( 
.A(n_1400),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_1400),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1419),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1419),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_1400),
.Y(n_2293)
);

NOR3xp33_ASAP7_75t_SL g2294 ( 
.A(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1426),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1208),
.B(n_858),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1426),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1008),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_1161),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_L g2303 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1426),
.Y(n_2304)
);

AOI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1426),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_L g2307 ( 
.A(n_1146),
.B(n_1431),
.Y(n_2307)
);

NOR2x1_ASAP7_75t_L g2308 ( 
.A(n_1140),
.B(n_1145),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_1400),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1426),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_1400),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_SL g2313 ( 
.A1(n_1433),
.A2(n_1457),
.B1(n_1478),
.B2(n_1458),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_L g2314 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_1159),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1189),
.B(n_1162),
.Y(n_2316)
);

INVx2_ASAP7_75t_SL g2317 ( 
.A(n_1161),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1426),
.Y(n_2318)
);

NOR2xp67_ASAP7_75t_L g2319 ( 
.A(n_1283),
.B(n_621),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1426),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1426),
.Y(n_2325)
);

NOR2xp67_ASAP7_75t_L g2326 ( 
.A(n_1283),
.B(n_621),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2328)
);

AOI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_1208),
.B(n_858),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_1208),
.B(n_858),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2332)
);

NOR2xp67_ASAP7_75t_L g2333 ( 
.A(n_1283),
.B(n_621),
.Y(n_2333)
);

AOI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1426),
.Y(n_2335)
);

AOI22xp33_ASAP7_75t_L g2336 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_1400),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_1572),
.B(n_1619),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1433),
.B(n_1457),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.Y(n_2341)
);

AND2x6_ASAP7_75t_SL g2342 ( 
.A(n_1647),
.B(n_2111),
.Y(n_2342)
);

AOI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2171),
.A2(n_1667),
.B1(n_2259),
.B2(n_2209),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_1790),
.B(n_2152),
.Y(n_2344)
);

INVxp67_ASAP7_75t_SL g2345 ( 
.A(n_1658),
.Y(n_2345)
);

NOR2xp33_ASAP7_75t_L g2346 ( 
.A(n_2195),
.B(n_2119),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2285),
.B(n_1635),
.Y(n_2347)
);

NAND2x1_ASAP7_75t_L g2348 ( 
.A(n_1837),
.B(n_1858),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1702),
.B(n_2165),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2212),
.B(n_2234),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2195),
.B(n_2269),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2281),
.B(n_2289),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_1727),
.B(n_1679),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2259),
.A2(n_2209),
.B1(n_2208),
.B2(n_2090),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_1635),
.B(n_2058),
.Y(n_2355)
);

AOI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_1767),
.A2(n_1784),
.B(n_1780),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_1727),
.B(n_1679),
.Y(n_2357)
);

AO21x1_ASAP7_75t_L g2358 ( 
.A1(n_1633),
.A2(n_2177),
.B(n_2142),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_1660),
.Y(n_2359)
);

AOI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_1767),
.A2(n_1784),
.B(n_1780),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_1766),
.B(n_1629),
.Y(n_2361)
);

OAI21x1_ASAP7_75t_L g2362 ( 
.A1(n_1969),
.A2(n_2026),
.B(n_1757),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1625),
.B(n_1627),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_1680),
.Y(n_2364)
);

AOI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_1788),
.A2(n_2307),
.B(n_2163),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2013),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2058),
.B(n_2097),
.Y(n_2367)
);

OAI21xp33_ASAP7_75t_L g2368 ( 
.A1(n_2136),
.A2(n_2294),
.B(n_2238),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_1625),
.B(n_1627),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_1788),
.A2(n_1798),
.B(n_1730),
.Y(n_2370)
);

BUFx2_ASAP7_75t_L g2371 ( 
.A(n_1701),
.Y(n_2371)
);

O2A1O1Ixp33_ASAP7_75t_L g2372 ( 
.A1(n_2104),
.A2(n_2177),
.B(n_2142),
.C(n_1633),
.Y(n_2372)
);

OAI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2104),
.A2(n_1690),
.B(n_1692),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_1630),
.B(n_1641),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1630),
.B(n_1641),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1673),
.B(n_1712),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_1798),
.A2(n_1730),
.B(n_1722),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1659),
.B(n_2048),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1659),
.B(n_2048),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2050),
.B(n_2056),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1628),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_2123),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_1673),
.B(n_1712),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1628),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2050),
.B(n_2056),
.Y(n_2385)
);

NOR2x1_ASAP7_75t_L g2386 ( 
.A(n_1942),
.B(n_2308),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_1722),
.A2(n_1757),
.B(n_1892),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1643),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_1892),
.A2(n_2308),
.B(n_2044),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2097),
.B(n_2148),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2064),
.B(n_2066),
.Y(n_2391)
);

NOR3xp33_ASAP7_75t_L g2392 ( 
.A(n_1661),
.B(n_1649),
.C(n_1638),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2064),
.B(n_2066),
.Y(n_2393)
);

AO22x1_ASAP7_75t_L g2394 ( 
.A1(n_2117),
.A2(n_1944),
.B1(n_1810),
.B2(n_1814),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_1637),
.A2(n_2088),
.B(n_2078),
.Y(n_2395)
);

BUFx12f_ASAP7_75t_L g2396 ( 
.A(n_1759),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2099),
.A2(n_2120),
.B(n_2118),
.Y(n_2397)
);

AOI33xp33_ASAP7_75t_L g2398 ( 
.A1(n_2093),
.A2(n_2313),
.A3(n_1656),
.B1(n_2129),
.B2(n_2138),
.B3(n_2134),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2072),
.B(n_2081),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1643),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2146),
.A2(n_2167),
.B(n_2159),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1643),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_1790),
.B(n_2152),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2117),
.A2(n_2148),
.B1(n_2214),
.B2(n_2193),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2072),
.B(n_2081),
.Y(n_2405)
);

OAI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2282),
.A2(n_1649),
.B(n_2181),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_1644),
.Y(n_2407)
);

INVxp67_ASAP7_75t_L g2408 ( 
.A(n_2051),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_1714),
.B(n_1716),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2341),
.A2(n_2214),
.B1(n_2217),
.B2(n_2193),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2189),
.A2(n_2229),
.B(n_2225),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2083),
.B(n_2085),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2217),
.B(n_2280),
.Y(n_2413)
);

AOI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_1654),
.A2(n_2313),
.B1(n_2093),
.B2(n_1684),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_1813),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2310),
.A2(n_2337),
.B(n_2321),
.Y(n_2416)
);

OR2x6_ASAP7_75t_L g2417 ( 
.A(n_1969),
.B(n_1823),
.Y(n_2417)
);

AOI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2339),
.A2(n_2036),
.B(n_2173),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2280),
.B(n_2287),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1650),
.Y(n_2420)
);

AOI21x1_ASAP7_75t_L g2421 ( 
.A1(n_1661),
.A2(n_1763),
.B(n_2025),
.Y(n_2421)
);

OAI21xp33_ASAP7_75t_L g2422 ( 
.A1(n_2070),
.A2(n_2221),
.B(n_2192),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2233),
.A2(n_2277),
.B1(n_2303),
.B2(n_2256),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1650),
.Y(n_2424)
);

AOI21xp5_ASAP7_75t_L g2425 ( 
.A1(n_2300),
.A2(n_1927),
.B(n_1861),
.Y(n_2425)
);

OA22x2_ASAP7_75t_L g2426 ( 
.A1(n_2287),
.A2(n_2305),
.B1(n_2334),
.B2(n_2329),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_1714),
.B(n_1716),
.Y(n_2427)
);

O2A1O1Ixp33_ASAP7_75t_L g2428 ( 
.A1(n_2201),
.A2(n_1703),
.B(n_1695),
.C(n_1677),
.Y(n_2428)
);

OAI22xp5_ASAP7_75t_SL g2429 ( 
.A1(n_2314),
.A2(n_2328),
.B1(n_2336),
.B2(n_2332),
.Y(n_2429)
);

CKINVDCx10_ASAP7_75t_R g2430 ( 
.A(n_2124),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2083),
.B(n_2085),
.Y(n_2431)
);

BUFx8_ASAP7_75t_L g2432 ( 
.A(n_1759),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_SL g2433 ( 
.A(n_2305),
.B(n_2329),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_1701),
.Y(n_2434)
);

NOR3xp33_ASAP7_75t_L g2435 ( 
.A(n_1677),
.B(n_1726),
.C(n_1782),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_1660),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2123),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1650),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_1631),
.Y(n_2439)
);

AOI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_1861),
.A2(n_2282),
.B(n_1734),
.Y(n_2440)
);

OAI21xp33_ASAP7_75t_L g2441 ( 
.A1(n_2334),
.A2(n_2341),
.B(n_2098),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2095),
.B(n_2098),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2095),
.B(n_2108),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1631),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_1734),
.A2(n_1973),
.B(n_1705),
.Y(n_2445)
);

OA22x2_ASAP7_75t_L g2446 ( 
.A1(n_1678),
.A2(n_1688),
.B1(n_1782),
.B2(n_1750),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2108),
.B(n_2109),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2109),
.B(n_2113),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2113),
.B(n_2125),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_1973),
.A2(n_1705),
.B(n_1950),
.Y(n_2450)
);

NOR2xp67_ASAP7_75t_L g2451 ( 
.A(n_1678),
.B(n_1811),
.Y(n_2451)
);

NAND3xp33_ASAP7_75t_L g2452 ( 
.A(n_1688),
.B(n_2126),
.C(n_2125),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2123),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_1950),
.A2(n_1810),
.B(n_1992),
.Y(n_2454)
);

AOI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2320),
.A2(n_2323),
.B1(n_2327),
.B2(n_2322),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2126),
.B(n_2141),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1655),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_1744),
.B(n_1766),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_1944),
.A2(n_1763),
.B(n_1719),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_SL g2460 ( 
.A(n_1858),
.B(n_1876),
.Y(n_2460)
);

NOR2x1p5_ASAP7_75t_L g2461 ( 
.A(n_1921),
.B(n_1938),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_1676),
.B(n_1681),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_1942),
.A2(n_2026),
.B(n_1847),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_1847),
.A2(n_1768),
.B(n_1786),
.Y(n_2464)
);

AOI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_1768),
.A2(n_1786),
.B(n_1812),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_2123),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2141),
.B(n_2144),
.Y(n_2467)
);

OA22x2_ASAP7_75t_L g2468 ( 
.A1(n_1750),
.A2(n_1866),
.B1(n_1805),
.B2(n_2149),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2144),
.B(n_2149),
.Y(n_2469)
);

O2A1O1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_2150),
.A2(n_2162),
.B(n_2175),
.C(n_2160),
.Y(n_2470)
);

A2O1A1Ixp33_ASAP7_75t_L g2471 ( 
.A1(n_1771),
.A2(n_2322),
.B(n_2323),
.C(n_2320),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2150),
.B(n_2160),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2162),
.B(n_2175),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_1622),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2180),
.B(n_2182),
.Y(n_2475)
);

NAND3xp33_ASAP7_75t_SL g2476 ( 
.A(n_2180),
.B(n_2183),
.C(n_2182),
.Y(n_2476)
);

OAI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2183),
.A2(n_2210),
.B1(n_2211),
.B2(n_2205),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2205),
.B(n_2210),
.Y(n_2478)
);

OAI21xp33_ASAP7_75t_L g2479 ( 
.A1(n_2211),
.A2(n_2237),
.B(n_2236),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_1744),
.B(n_1793),
.Y(n_2480)
);

O2A1O1Ixp33_ASAP7_75t_L g2481 ( 
.A1(n_2236),
.A2(n_2243),
.B(n_2248),
.C(n_2237),
.Y(n_2481)
);

NOR3xp33_ASAP7_75t_L g2482 ( 
.A(n_1726),
.B(n_2248),
.C(n_2243),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_2327),
.A2(n_2340),
.B1(n_2253),
.B2(n_2275),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1622),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_1812),
.A2(n_1760),
.B(n_2031),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2253),
.B(n_2268),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2268),
.B(n_2275),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_1744),
.B(n_1793),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_1760),
.A2(n_1707),
.B(n_1877),
.Y(n_2489)
);

O2A1O1Ixp33_ASAP7_75t_L g2490 ( 
.A1(n_2278),
.A2(n_2298),
.B(n_2299),
.C(n_2288),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_1707),
.A2(n_1823),
.B(n_1785),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_1676),
.B(n_1681),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_1744),
.B(n_1972),
.Y(n_2493)
);

O2A1O1Ixp33_ASAP7_75t_L g2494 ( 
.A1(n_2278),
.A2(n_2298),
.B(n_2299),
.C(n_2288),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_2302),
.B(n_2340),
.Y(n_2495)
);

OR2x4_ASAP7_75t_L g2496 ( 
.A(n_1901),
.B(n_2033),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_SL g2497 ( 
.A(n_1683),
.B(n_1686),
.Y(n_2497)
);

O2A1O1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_2302),
.A2(n_1686),
.B(n_1691),
.C(n_1683),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_1691),
.B(n_1693),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_1693),
.B(n_1700),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2139),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_1672),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_1940),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_1682),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_1700),
.B(n_1704),
.Y(n_2505)
);

OAI22xp5_ASAP7_75t_L g2506 ( 
.A1(n_1704),
.A2(n_1769),
.B1(n_1648),
.B2(n_1634),
.Y(n_2506)
);

CKINVDCx16_ASAP7_75t_R g2507 ( 
.A(n_2052),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_1823),
.A2(n_1785),
.B(n_2025),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_1823),
.A2(n_1785),
.B(n_2025),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_1823),
.A2(n_1785),
.B(n_1989),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_1741),
.B(n_1746),
.Y(n_2511)
);

INVxp67_ASAP7_75t_L g2512 ( 
.A(n_2075),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2139),
.Y(n_2513)
);

AOI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_1738),
.A2(n_1771),
.B1(n_1755),
.B2(n_1866),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_1741),
.B(n_1746),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_1682),
.Y(n_2516)
);

OAI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_1634),
.A2(n_1648),
.B1(n_1865),
.B2(n_1882),
.Y(n_2517)
);

O2A1O1Ixp5_ASAP7_75t_L g2518 ( 
.A1(n_1860),
.A2(n_1946),
.B(n_1903),
.C(n_2039),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_1865),
.A2(n_1882),
.B1(n_1804),
.B2(n_1756),
.Y(n_2519)
);

INVx4_ASAP7_75t_L g2520 ( 
.A(n_1811),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_1756),
.B(n_2063),
.Y(n_2521)
);

OAI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_1735),
.A2(n_1754),
.B1(n_1834),
.B2(n_1863),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_1811),
.A2(n_2096),
.B(n_1848),
.Y(n_2523)
);

BUFx4f_ASAP7_75t_L g2524 ( 
.A(n_1640),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_1761),
.A2(n_2326),
.B(n_2333),
.C(n_2319),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2207),
.B(n_2250),
.Y(n_2526)
);

AOI21x1_ASAP7_75t_L g2527 ( 
.A1(n_2319),
.A2(n_2333),
.B(n_2326),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2139),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_2130),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_L g2530 ( 
.A(n_1724),
.B(n_1738),
.C(n_1867),
.Y(n_2530)
);

NAND2x1p5_ASAP7_75t_L g2531 ( 
.A(n_1811),
.B(n_1848),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2063),
.B(n_2143),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_1624),
.Y(n_2533)
);

BUFx12f_ASAP7_75t_L g2534 ( 
.A(n_1759),
.Y(n_2534)
);

AOI21xp5_ASAP7_75t_L g2535 ( 
.A1(n_1811),
.A2(n_2096),
.B(n_1848),
.Y(n_2535)
);

OAI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_1717),
.A2(n_1720),
.B(n_1910),
.Y(n_2536)
);

A2O1A1Ixp33_ASAP7_75t_L g2537 ( 
.A1(n_1919),
.A2(n_2005),
.B(n_1976),
.C(n_1996),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2143),
.B(n_2188),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_1754),
.A2(n_1863),
.B1(n_1878),
.B2(n_1874),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2207),
.B(n_2250),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_SL g2541 ( 
.A(n_1921),
.Y(n_2541)
);

NOR2x1_ASAP7_75t_L g2542 ( 
.A(n_1930),
.B(n_1939),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_1624),
.Y(n_2543)
);

OAI22xp5_ASAP7_75t_L g2544 ( 
.A1(n_1874),
.A2(n_1878),
.B1(n_1887),
.B2(n_1815),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1685),
.Y(n_2545)
);

NOR2x1_ASAP7_75t_R g2546 ( 
.A(n_2252),
.B(n_1626),
.Y(n_2546)
);

NOR2x1_ASAP7_75t_L g2547 ( 
.A(n_1930),
.B(n_1939),
.Y(n_2547)
);

A2O1A1Ixp33_ASAP7_75t_L g2548 ( 
.A1(n_1996),
.A2(n_1720),
.B(n_1717),
.C(n_2042),
.Y(n_2548)
);

OAI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_1887),
.A2(n_1815),
.B1(n_1711),
.B2(n_1809),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_1723),
.B(n_1733),
.Y(n_2550)
);

BUFx3_ASAP7_75t_L g2551 ( 
.A(n_1813),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_1725),
.A2(n_1932),
.B1(n_1841),
.B2(n_1718),
.Y(n_2552)
);

NAND2x1_ASAP7_75t_L g2553 ( 
.A(n_1837),
.B(n_1858),
.Y(n_2553)
);

A2O1A1Ixp33_ASAP7_75t_L g2554 ( 
.A1(n_2042),
.A2(n_1982),
.B(n_2040),
.C(n_1862),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_1972),
.B(n_1694),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2188),
.B(n_2190),
.Y(n_2556)
);

NOR2xp33_ASAP7_75t_SL g2557 ( 
.A(n_1858),
.B(n_1876),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2102),
.A2(n_2240),
.B(n_2156),
.Y(n_2558)
);

BUFx4f_ASAP7_75t_L g2559 ( 
.A(n_1640),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_1629),
.B(n_2172),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2190),
.B(n_2230),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2230),
.B(n_2254),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2065),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2156),
.A2(n_2245),
.B(n_2240),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2202),
.Y(n_2565)
);

XNOR2xp5_ASAP7_75t_L g2566 ( 
.A(n_1687),
.B(n_2124),
.Y(n_2566)
);

AND2x2_ASAP7_75t_SL g2567 ( 
.A(n_2139),
.B(n_2263),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2156),
.A2(n_2245),
.B(n_2240),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_1680),
.Y(n_2569)
);

NAND2x1p5_ASAP7_75t_L g2570 ( 
.A(n_2240),
.B(n_2245),
.Y(n_2570)
);

AOI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2245),
.A2(n_2255),
.B(n_1846),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2254),
.B(n_2267),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2267),
.B(n_2296),
.Y(n_2573)
);

AO21x1_ASAP7_75t_L g2574 ( 
.A1(n_1910),
.A2(n_2016),
.B(n_1715),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2245),
.A2(n_2255),
.B(n_1846),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_1694),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2296),
.B(n_2330),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2330),
.B(n_2331),
.Y(n_2578)
);

OA22x2_ASAP7_75t_L g2579 ( 
.A1(n_1805),
.A2(n_1687),
.B1(n_2179),
.B2(n_2152),
.Y(n_2579)
);

OAI21xp5_ASAP7_75t_L g2580 ( 
.A1(n_1910),
.A2(n_1697),
.B(n_2015),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2245),
.A2(n_2255),
.B(n_1846),
.Y(n_2581)
);

OAI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_1808),
.A2(n_1836),
.B1(n_1725),
.B2(n_1890),
.Y(n_2582)
);

AOI22xp33_ASAP7_75t_L g2583 ( 
.A1(n_2172),
.A2(n_1715),
.B1(n_1721),
.B2(n_1713),
.Y(n_2583)
);

A2O1A1Ixp33_ASAP7_75t_L g2584 ( 
.A1(n_1982),
.A2(n_2040),
.B(n_1832),
.C(n_1979),
.Y(n_2584)
);

AOI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2255),
.A2(n_1846),
.B(n_1721),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2331),
.B(n_1739),
.Y(n_2586)
);

BUFx2_ASAP7_75t_L g2587 ( 
.A(n_1940),
.Y(n_2587)
);

BUFx12f_ASAP7_75t_L g2588 ( 
.A(n_2252),
.Y(n_2588)
);

OAI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_1987),
.A2(n_1994),
.B(n_1993),
.Y(n_2589)
);

OAI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_1987),
.A2(n_1994),
.B(n_1993),
.Y(n_2590)
);

INVx2_ASAP7_75t_SL g2591 ( 
.A(n_1818),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_1739),
.B(n_1954),
.Y(n_2592)
);

INVxp67_ASAP7_75t_L g2593 ( 
.A(n_2315),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_1954),
.B(n_1748),
.Y(n_2594)
);

BUFx6f_ASAP7_75t_L g2595 ( 
.A(n_2263),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_1819),
.B(n_1833),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_1857),
.A2(n_1889),
.B(n_1884),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_1940),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_1889),
.A2(n_1884),
.B(n_1876),
.Y(n_2599)
);

OAI21x1_ASAP7_75t_L g2600 ( 
.A1(n_1660),
.A2(n_1689),
.B(n_1671),
.Y(n_2600)
);

OAI21xp33_ASAP7_75t_L g2601 ( 
.A1(n_1819),
.A2(n_1839),
.B(n_1833),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_1884),
.A2(n_1964),
.B(n_1963),
.Y(n_2602)
);

O2A1O1Ixp33_ASAP7_75t_L g2603 ( 
.A1(n_1789),
.A2(n_1830),
.B(n_1891),
.C(n_1743),
.Y(n_2603)
);

BUFx12f_ASAP7_75t_L g2604 ( 
.A(n_2252),
.Y(n_2604)
);

NOR2x1_ASAP7_75t_L g2605 ( 
.A(n_1930),
.B(n_1939),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2147),
.B(n_2270),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_1710),
.Y(n_2607)
);

NAND2x1_ASAP7_75t_L g2608 ( 
.A(n_1837),
.B(n_1930),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_1839),
.B(n_1843),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_1843),
.B(n_1845),
.Y(n_2610)
);

NAND2xp33_ASAP7_75t_L g2611 ( 
.A(n_1698),
.B(n_2047),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1710),
.Y(n_2612)
);

A2O1A1Ixp33_ASAP7_75t_L g2613 ( 
.A1(n_1979),
.A2(n_2039),
.B(n_1999),
.C(n_2000),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_1671),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_1710),
.Y(n_2615)
);

A2O1A1Ixp33_ASAP7_75t_L g2616 ( 
.A1(n_1995),
.A2(n_2000),
.B(n_1999),
.C(n_2035),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2147),
.B(n_2270),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_1845),
.B(n_1758),
.Y(n_2618)
);

O2A1O1Ixp33_ASAP7_75t_L g2619 ( 
.A1(n_2068),
.A2(n_2076),
.B(n_2176),
.C(n_2131),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_1890),
.A2(n_1904),
.B1(n_1915),
.B2(n_1896),
.Y(n_2620)
);

A2O1A1Ixp33_ASAP7_75t_L g2621 ( 
.A1(n_1995),
.A2(n_2035),
.B(n_1871),
.C(n_2020),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2271),
.B(n_1636),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_2271),
.B(n_1642),
.Y(n_2623)
);

BUFx6f_ASAP7_75t_L g2624 ( 
.A(n_2263),
.Y(n_2624)
);

OAI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_1896),
.A2(n_1904),
.B1(n_1915),
.B2(n_1758),
.Y(n_2625)
);

INVxp67_ASAP7_75t_L g2626 ( 
.A(n_2046),
.Y(n_2626)
);

AOI21xp5_ASAP7_75t_L g2627 ( 
.A1(n_1728),
.A2(n_1850),
.B(n_1842),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_1752),
.Y(n_2628)
);

AOI21xp5_ASAP7_75t_L g2629 ( 
.A1(n_1842),
.A2(n_1855),
.B(n_1850),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_1851),
.B(n_1909),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_1855),
.A2(n_2263),
.B(n_1985),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2067),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_1821),
.B(n_1900),
.Y(n_2633)
);

O2A1O1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2206),
.A2(n_2247),
.B(n_1706),
.C(n_1880),
.Y(n_2634)
);

AOI21x1_ASAP7_75t_L g2635 ( 
.A1(n_2001),
.A2(n_2006),
.B(n_2002),
.Y(n_2635)
);

INVx2_ASAP7_75t_SL g2636 ( 
.A(n_1818),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_1837),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_1909),
.B(n_1777),
.Y(n_2638)
);

AOI21x1_ASAP7_75t_L g2639 ( 
.A1(n_2002),
.A2(n_2006),
.B(n_2041),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_1777),
.B(n_2046),
.Y(n_2640)
);

AOI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_1932),
.A2(n_2011),
.B(n_2152),
.Y(n_2641)
);

OAI21xp33_ASAP7_75t_L g2642 ( 
.A1(n_1908),
.A2(n_1791),
.B(n_1905),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_1826),
.B(n_1787),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2049),
.B(n_2071),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_1752),
.B(n_1762),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_1640),
.Y(n_2646)
);

OAI21x1_ASAP7_75t_L g2647 ( 
.A1(n_1747),
.A2(n_1831),
.B(n_2011),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_1762),
.Y(n_2648)
);

NOR2x1_ASAP7_75t_R g2649 ( 
.A(n_2054),
.B(n_2073),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2067),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_1645),
.A2(n_1646),
.B1(n_2053),
.B2(n_2045),
.Y(n_2651)
);

INVx4_ASAP7_75t_L g2652 ( 
.A(n_2257),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2077),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2153),
.Y(n_2654)
);

BUFx6f_ASAP7_75t_L g2655 ( 
.A(n_1640),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2152),
.A2(n_2264),
.B(n_2179),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2049),
.B(n_2071),
.Y(n_2657)
);

AOI221xp5_ASAP7_75t_L g2658 ( 
.A1(n_1854),
.A2(n_2121),
.B1(n_1961),
.B2(n_1941),
.C(n_1816),
.Y(n_2658)
);

AOI33xp33_ASAP7_75t_L g2659 ( 
.A1(n_1981),
.A2(n_2014),
.A3(n_1662),
.B1(n_1657),
.B2(n_1670),
.B3(n_1666),
.Y(n_2659)
);

A2O1A1Ixp33_ASAP7_75t_L g2660 ( 
.A1(n_2035),
.A2(n_1828),
.B(n_2041),
.C(n_2038),
.Y(n_2660)
);

OAI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2014),
.A2(n_2007),
.B(n_2010),
.Y(n_2661)
);

O2A1O1Ixp5_ASAP7_75t_L g2662 ( 
.A1(n_1907),
.A2(n_1745),
.B(n_1879),
.C(n_2038),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2179),
.A2(n_2264),
.B(n_1959),
.Y(n_2663)
);

NAND2xp33_ASAP7_75t_L g2664 ( 
.A(n_2158),
.B(n_2185),
.Y(n_2664)
);

INVx4_ASAP7_75t_L g2665 ( 
.A(n_2257),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_SL g2666 ( 
.A(n_2121),
.B(n_1828),
.Y(n_2666)
);

AND2x6_ASAP7_75t_L g2667 ( 
.A(n_1663),
.B(n_1802),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_1762),
.B(n_1772),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_1828),
.B(n_1699),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_1632),
.B(n_1639),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_1828),
.B(n_1774),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_1632),
.B(n_1639),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_1632),
.B(n_1639),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_SL g2674 ( 
.A(n_1729),
.B(n_1770),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2264),
.A2(n_1959),
.B(n_1929),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_1632),
.B(n_1639),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_1665),
.B(n_2057),
.Y(n_2677)
);

INVx2_ASAP7_75t_SL g2678 ( 
.A(n_1959),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_1665),
.B(n_2057),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2074),
.Y(n_2680)
);

AOI21x1_ASAP7_75t_L g2681 ( 
.A1(n_2007),
.A2(n_2010),
.B(n_2038),
.Y(n_2681)
);

AOI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_1959),
.A2(n_1929),
.B(n_1920),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_1665),
.B(n_2057),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_1665),
.B(n_2057),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2074),
.Y(n_2685)
);

OAI21xp33_ASAP7_75t_L g2686 ( 
.A1(n_1645),
.A2(n_2045),
.B(n_1646),
.Y(n_2686)
);

A2O1A1Ixp33_ASAP7_75t_L g2687 ( 
.A1(n_2038),
.A2(n_1805),
.B(n_1790),
.C(n_1675),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2087),
.B(n_2092),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_1920),
.A2(n_1929),
.B(n_1775),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_1940),
.A2(n_1675),
.B1(n_1708),
.B2(n_1668),
.Y(n_2690)
);

BUFx12f_ASAP7_75t_L g2691 ( 
.A(n_1674),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_1940),
.A2(n_1675),
.B1(n_1708),
.B2(n_1668),
.Y(n_2692)
);

AOI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_1920),
.A2(n_1775),
.B(n_1770),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_1645),
.A2(n_1646),
.B1(n_2053),
.B2(n_2045),
.Y(n_2694)
);

AOI21xp5_ASAP7_75t_L g2695 ( 
.A1(n_1770),
.A2(n_1775),
.B(n_1939),
.Y(n_2695)
);

OAI21xp5_ASAP7_75t_L g2696 ( 
.A1(n_1747),
.A2(n_1831),
.B(n_1974),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_1770),
.A2(n_1775),
.B(n_1802),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2087),
.B(n_2092),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2087),
.B(n_2092),
.Y(n_2699)
);

INVxp67_ASAP7_75t_L g2700 ( 
.A(n_1796),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2087),
.B(n_2092),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_1975),
.B(n_1772),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_1802),
.A2(n_1924),
.B(n_1916),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2100),
.B(n_2145),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_1802),
.A2(n_1924),
.B(n_1916),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_1772),
.B(n_1778),
.Y(n_2706)
);

AOI21x1_ASAP7_75t_L g2707 ( 
.A1(n_1621),
.A2(n_2059),
.B(n_2043),
.Y(n_2707)
);

BUFx12f_ASAP7_75t_L g2708 ( 
.A(n_1674),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2100),
.B(n_2145),
.Y(n_2709)
);

NAND3xp33_ASAP7_75t_L g2710 ( 
.A(n_1956),
.B(n_1962),
.C(n_1674),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2100),
.B(n_2145),
.Y(n_2711)
);

CKINVDCx16_ASAP7_75t_R g2712 ( 
.A(n_1807),
.Y(n_2712)
);

AOI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_1925),
.A2(n_1928),
.B(n_1926),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2074),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_1778),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_1925),
.A2(n_1928),
.B(n_1926),
.Y(n_2716)
);

O2A1O1Ixp33_ASAP7_75t_L g2717 ( 
.A1(n_1875),
.A2(n_1801),
.B(n_1949),
.C(n_2053),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_1640),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2100),
.B(n_2145),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_1778),
.B(n_1817),
.Y(n_2720)
);

NOR2x1_ASAP7_75t_L g2721 ( 
.A(n_1668),
.B(n_1708),
.Y(n_2721)
);

INVx1_ASAP7_75t_SL g2722 ( 
.A(n_1906),
.Y(n_2722)
);

AOI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_1933),
.A2(n_1951),
.B(n_1945),
.Y(n_2723)
);

BUFx2_ASAP7_75t_L g2724 ( 
.A(n_1940),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2200),
.B(n_2223),
.Y(n_2725)
);

NAND2x1_ASAP7_75t_L g2726 ( 
.A(n_1837),
.B(n_1940),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2200),
.B(n_2223),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_1817),
.B(n_1870),
.Y(n_2728)
);

AOI21x1_ASAP7_75t_L g2729 ( 
.A1(n_1621),
.A2(n_2059),
.B(n_2043),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_1841),
.B(n_2220),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2200),
.B(n_2223),
.Y(n_2731)
);

O2A1O1Ixp33_ASAP7_75t_L g2732 ( 
.A1(n_2069),
.A2(n_2101),
.B(n_2178),
.C(n_2137),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_1933),
.A2(n_1951),
.B(n_1945),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_1870),
.B(n_1912),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2069),
.A2(n_2137),
.B(n_2178),
.C(n_2101),
.Y(n_2735)
);

AOI21x1_ASAP7_75t_L g2736 ( 
.A1(n_2061),
.A2(n_2086),
.B(n_2062),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_1651),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_1837),
.Y(n_2738)
);

AOI21xp5_ASAP7_75t_L g2739 ( 
.A1(n_1958),
.A2(n_1975),
.B(n_1751),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2200),
.B(n_2223),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_1912),
.B(n_1913),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_1841),
.B(n_2272),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2316),
.B(n_1913),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_1917),
.B(n_1918),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2316),
.B(n_1917),
.Y(n_2745)
);

AOI33xp33_ASAP7_75t_L g2746 ( 
.A1(n_1651),
.A2(n_1779),
.A3(n_1776),
.B1(n_1773),
.B2(n_1765),
.B3(n_1657),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2089),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2316),
.B(n_1918),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2316),
.B(n_1662),
.Y(n_2749)
);

OAI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2069),
.A2(n_2137),
.B1(n_2178),
.B2(n_2101),
.Y(n_2750)
);

A2O1A1Ixp33_ASAP7_75t_L g2751 ( 
.A1(n_2231),
.A2(n_2258),
.B(n_2244),
.C(n_2061),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_1948),
.B(n_2231),
.Y(n_2752)
);

NOR2x1_ASAP7_75t_L g2753 ( 
.A(n_1623),
.B(n_2060),
.Y(n_2753)
);

A2O1A1Ixp33_ASAP7_75t_L g2754 ( 
.A1(n_2231),
.A2(n_2258),
.B(n_2244),
.C(n_2062),
.Y(n_2754)
);

OAI321xp33_ASAP7_75t_L g2755 ( 
.A1(n_1998),
.A2(n_2122),
.A3(n_2335),
.B1(n_2325),
.B2(n_2324),
.C(n_2107),
.Y(n_2755)
);

A2O1A1Ixp33_ASAP7_75t_L g2756 ( 
.A1(n_2244),
.A2(n_2258),
.B(n_2086),
.C(n_2106),
.Y(n_2756)
);

OAI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2105),
.A2(n_2106),
.B1(n_2122),
.B2(n_2107),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_1897),
.B(n_1822),
.Y(n_2758)
);

CKINVDCx8_ASAP7_75t_R g2759 ( 
.A(n_1948),
.Y(n_2759)
);

A2O1A1Ixp33_ASAP7_75t_L g2760 ( 
.A1(n_2105),
.A2(n_2128),
.B(n_2157),
.C(n_2151),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_1740),
.A2(n_2079),
.B(n_1751),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_1740),
.A2(n_2079),
.B(n_1751),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_1837),
.Y(n_2763)
);

CKINVDCx14_ASAP7_75t_R g2764 ( 
.A(n_1849),
.Y(n_2764)
);

OAI21xp33_ASAP7_75t_L g2765 ( 
.A1(n_2128),
.A2(n_2157),
.B(n_2151),
.Y(n_2765)
);

O2A1O1Ixp33_ASAP7_75t_L g2766 ( 
.A1(n_2022),
.A2(n_1990),
.B(n_1998),
.C(n_1906),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2089),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_1696),
.B(n_1709),
.Y(n_2768)
);

NOR2xp33_ASAP7_75t_L g2769 ( 
.A(n_1807),
.B(n_1822),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_1740),
.A2(n_2115),
.B(n_2079),
.Y(n_2770)
);

OAI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_2161),
.A2(n_2169),
.B1(n_2187),
.B2(n_2170),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_1640),
.Y(n_2772)
);

CKINVDCx20_ASAP7_75t_R g2773 ( 
.A(n_1674),
.Y(n_2773)
);

A2O1A1Ixp33_ASAP7_75t_L g2774 ( 
.A1(n_2161),
.A2(n_2169),
.B(n_2187),
.C(n_2170),
.Y(n_2774)
);

O2A1O1Ixp33_ASAP7_75t_L g2775 ( 
.A1(n_2022),
.A2(n_1990),
.B(n_1653),
.C(n_1664),
.Y(n_2775)
);

OAI21x1_ASAP7_75t_L g2776 ( 
.A1(n_2089),
.A2(n_2110),
.B(n_2094),
.Y(n_2776)
);

NAND3xp33_ASAP7_75t_L g2777 ( 
.A(n_2132),
.B(n_2140),
.C(n_1732),
.Y(n_2777)
);

O2A1O1Ixp33_ASAP7_75t_L g2778 ( 
.A1(n_1653),
.A2(n_1664),
.B(n_1822),
.C(n_1974),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_1731),
.B(n_1736),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_1736),
.Y(n_2780)
);

NOR2xp67_ASAP7_75t_L g2781 ( 
.A(n_1623),
.B(n_2060),
.Y(n_2781)
);

O2A1O1Ixp5_ASAP7_75t_L g2782 ( 
.A1(n_1980),
.A2(n_1986),
.B(n_2017),
.C(n_1983),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_1737),
.B(n_1742),
.Y(n_2783)
);

OR2x2_ASAP7_75t_L g2784 ( 
.A(n_1749),
.B(n_1753),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_1749),
.B(n_1753),
.Y(n_2785)
);

A2O1A1Ixp33_ASAP7_75t_L g2786 ( 
.A1(n_2191),
.A2(n_2196),
.B(n_2335),
.C(n_2325),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2094),
.Y(n_2787)
);

A2O1A1Ixp33_ASAP7_75t_L g2788 ( 
.A1(n_2191),
.A2(n_2265),
.B(n_2324),
.C(n_2318),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2196),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2197),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_1729),
.B(n_1664),
.Y(n_2791)
);

AOI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2246),
.A2(n_2301),
.B(n_2249),
.Y(n_2792)
);

INVxp67_ASAP7_75t_L g2793 ( 
.A(n_1997),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_1897),
.B(n_1623),
.Y(n_2794)
);

CKINVDCx5p33_ASAP7_75t_R g2795 ( 
.A(n_2132),
.Y(n_2795)
);

AOI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2249),
.A2(n_2317),
.B(n_2301),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2317),
.A2(n_2216),
.B(n_2084),
.Y(n_2797)
);

NOR2xp67_ASAP7_75t_L g2798 ( 
.A(n_1623),
.B(n_2060),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_1764),
.B(n_2226),
.Y(n_2799)
);

AND2x2_ASAP7_75t_SL g2800 ( 
.A(n_1663),
.B(n_2338),
.Y(n_2800)
);

NAND2x1p5_ASAP7_75t_L g2801 ( 
.A(n_2060),
.B(n_2080),
.Y(n_2801)
);

OAI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_1940),
.A2(n_1792),
.B(n_1783),
.Y(n_2802)
);

O2A1O1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_1764),
.A2(n_2261),
.B(n_2226),
.C(n_2318),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_SL g2804 ( 
.A(n_2261),
.B(n_2027),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2197),
.B(n_2203),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2317),
.A2(n_2216),
.B(n_2084),
.Y(n_2806)
);

NOR2xp67_ASAP7_75t_L g2807 ( 
.A(n_2080),
.B(n_2114),
.Y(n_2807)
);

A2O1A1Ixp33_ASAP7_75t_L g2808 ( 
.A1(n_2203),
.A2(n_2215),
.B(n_2213),
.C(n_2306),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2084),
.A2(n_2241),
.B(n_2216),
.Y(n_2809)
);

AOI221xp5_ASAP7_75t_L g2810 ( 
.A1(n_1921),
.A2(n_1938),
.B1(n_2213),
.B2(n_2311),
.C(n_2215),
.Y(n_2810)
);

NAND3xp33_ASAP7_75t_L g2811 ( 
.A(n_2132),
.B(n_2140),
.C(n_1997),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2222),
.A2(n_2265),
.B1(n_2283),
.B2(n_2224),
.Y(n_2812)
);

O2A1O1Ixp33_ASAP7_75t_L g2813 ( 
.A1(n_2222),
.A2(n_2283),
.B(n_2279),
.C(n_2276),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2241),
.A2(n_2242),
.B(n_2232),
.Y(n_2814)
);

AND2x2_ASAP7_75t_SL g2815 ( 
.A(n_1663),
.B(n_1652),
.Y(n_2815)
);

AOI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2082),
.A2(n_1991),
.B1(n_1935),
.B2(n_1977),
.Y(n_2816)
);

AO21x1_ASAP7_75t_L g2817 ( 
.A1(n_2224),
.A2(n_2239),
.B(n_2232),
.Y(n_2817)
);

AND3x2_ASAP7_75t_L g2818 ( 
.A(n_1971),
.B(n_2009),
.C(n_2023),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2239),
.Y(n_2819)
);

NAND3xp33_ASAP7_75t_L g2820 ( 
.A(n_2132),
.B(n_2140),
.C(n_2251),
.Y(n_2820)
);

AOI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2241),
.A2(n_2242),
.B(n_2251),
.Y(n_2821)
);

O2A1O1Ixp33_ASAP7_75t_SL g2822 ( 
.A1(n_2019),
.A2(n_2029),
.B(n_2030),
.C(n_2297),
.Y(n_2822)
);

INVxp67_ASAP7_75t_L g2823 ( 
.A(n_2023),
.Y(n_2823)
);

OAI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2260),
.A2(n_2306),
.B1(n_2297),
.B2(n_2311),
.Y(n_2824)
);

AOI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2082),
.A2(n_1968),
.B1(n_1938),
.B2(n_2295),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_SL g2826 ( 
.A(n_2018),
.B(n_1923),
.Y(n_2826)
);

O2A1O1Ixp33_ASAP7_75t_SL g2827 ( 
.A1(n_2030),
.A2(n_2266),
.B(n_2295),
.C(n_2273),
.Y(n_2827)
);

BUFx8_ASAP7_75t_SL g2828 ( 
.A(n_1652),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2242),
.A2(n_2266),
.B(n_2260),
.Y(n_2829)
);

AOI21x1_ASAP7_75t_L g2830 ( 
.A1(n_2273),
.A2(n_2276),
.B(n_2274),
.Y(n_2830)
);

BUFx2_ASAP7_75t_L g2831 ( 
.A(n_1729),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2024),
.B(n_1781),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2274),
.A2(n_2279),
.B(n_2304),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2304),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_1966),
.B(n_1967),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_1886),
.B(n_1914),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_1837),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2112),
.A2(n_2174),
.B(n_2135),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_1966),
.B(n_1967),
.Y(n_2839)
);

INVx4_ASAP7_75t_L g2840 ( 
.A(n_2257),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2112),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_1783),
.A2(n_1955),
.B(n_1936),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_1886),
.B(n_2257),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_1966),
.B(n_1967),
.Y(n_2844)
);

AO22x1_ASAP7_75t_L g2845 ( 
.A1(n_2140),
.A2(n_1663),
.B1(n_2312),
.B2(n_2290),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_1794),
.B(n_1797),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_1984),
.A2(n_1895),
.B1(n_1947),
.B2(n_1955),
.Y(n_2847)
);

O2A1O1Ixp33_ASAP7_75t_L g2848 ( 
.A1(n_1984),
.A2(n_1872),
.B(n_1960),
.C(n_1947),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_SL g2849 ( 
.A(n_2257),
.B(n_1663),
.Y(n_2849)
);

AOI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2133),
.A2(n_2186),
.B(n_2184),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_1827),
.B(n_1829),
.Y(n_2851)
);

INVx5_ASAP7_75t_L g2852 ( 
.A(n_1663),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_1652),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_1827),
.B(n_1829),
.Y(n_2854)
);

NAND2xp33_ASAP7_75t_L g2855 ( 
.A(n_1652),
.B(n_2055),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_1859),
.B(n_1652),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_1827),
.B(n_1829),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2135),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_1984),
.A2(n_1840),
.B1(n_1960),
.B2(n_1937),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_1799),
.A2(n_1872),
.B1(n_1936),
.B2(n_1856),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_1803),
.A2(n_1835),
.B1(n_1856),
.B2(n_1895),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2154),
.Y(n_2862)
);

AND2x4_ASAP7_75t_L g2863 ( 
.A(n_2080),
.B(n_2114),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_1781),
.B(n_1825),
.Y(n_2864)
);

OR2x6_ASAP7_75t_L g2865 ( 
.A(n_1652),
.B(n_2055),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_1844),
.B(n_1852),
.Y(n_2866)
);

BUFx3_ASAP7_75t_L g2867 ( 
.A(n_1781),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_1844),
.B(n_1852),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_1859),
.B(n_2338),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_1844),
.B(n_1852),
.Y(n_2870)
);

A2O1A1Ixp33_ASAP7_75t_L g2871 ( 
.A1(n_2080),
.A2(n_2290),
.B(n_2312),
.C(n_2286),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2164),
.Y(n_2872)
);

BUFx4f_ASAP7_75t_L g2873 ( 
.A(n_2055),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2164),
.Y(n_2874)
);

AOI21x1_ASAP7_75t_L g2875 ( 
.A1(n_1803),
.A2(n_1835),
.B(n_1893),
.Y(n_2875)
);

BUFx2_ASAP7_75t_L g2876 ( 
.A(n_1795),
.Y(n_2876)
);

AOI22xp33_ASAP7_75t_L g2877 ( 
.A1(n_1820),
.A2(n_1873),
.B1(n_1824),
.B2(n_1883),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_1868),
.B(n_1869),
.Y(n_2878)
);

NOR3xp33_ASAP7_75t_L g2879 ( 
.A(n_2114),
.B(n_2218),
.C(n_2312),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2166),
.Y(n_2880)
);

OAI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_1820),
.A2(n_1873),
.B(n_1824),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_R g2882 ( 
.A(n_2055),
.B(n_2091),
.Y(n_2882)
);

O2A1O1Ixp33_ASAP7_75t_SL g2883 ( 
.A1(n_1881),
.A2(n_1899),
.B(n_1898),
.C(n_1894),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_1868),
.B(n_1869),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_1868),
.B(n_1869),
.Y(n_2885)
);

AOI21x1_ASAP7_75t_L g2886 ( 
.A1(n_1838),
.A2(n_1853),
.B(n_1893),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2168),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_1965),
.B(n_1978),
.Y(n_2888)
);

OAI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_1825),
.A2(n_1883),
.B1(n_1838),
.B2(n_1853),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_1825),
.B(n_1965),
.Y(n_2890)
);

AOI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_1864),
.A2(n_1978),
.B1(n_1859),
.B2(n_1952),
.Y(n_2891)
);

A2O1A1Ixp33_ASAP7_75t_L g2892 ( 
.A1(n_2114),
.A2(n_2199),
.B(n_2218),
.C(n_2290),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_1885),
.B(n_1953),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_SL g2894 ( 
.A(n_1859),
.B(n_2338),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_1885),
.B(n_1934),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_1885),
.B(n_1934),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_1881),
.Y(n_2897)
);

OAI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_1864),
.A2(n_1953),
.B(n_1952),
.Y(n_2898)
);

INVx1_ASAP7_75t_SL g2899 ( 
.A(n_1971),
.Y(n_2899)
);

NAND2x1p5_ASAP7_75t_L g2900 ( 
.A(n_2127),
.B(n_2312),
.Y(n_2900)
);

A2O1A1Ixp33_ASAP7_75t_L g2901 ( 
.A1(n_2127),
.A2(n_2286),
.B(n_2199),
.C(n_2218),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_R g2902 ( 
.A(n_2055),
.B(n_2338),
.Y(n_2902)
);

AOI22x1_ASAP7_75t_L g2903 ( 
.A1(n_1888),
.A2(n_1934),
.B1(n_1953),
.B2(n_1952),
.Y(n_2903)
);

INVx3_ASAP7_75t_L g2904 ( 
.A(n_1881),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2227),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2228),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_1888),
.B(n_1922),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_1881),
.Y(n_2908)
);

OR2x6_ASAP7_75t_SL g2909 ( 
.A(n_1806),
.B(n_2198),
.Y(n_2909)
);

O2A1O1Ixp33_ASAP7_75t_L g2910 ( 
.A1(n_2127),
.A2(n_2199),
.B(n_2218),
.C(n_2286),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2338),
.B(n_2055),
.Y(n_2911)
);

INVx5_ASAP7_75t_L g2912 ( 
.A(n_1894),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2235),
.A2(n_2262),
.B1(n_2284),
.B2(n_2292),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_2091),
.Y(n_2914)
);

AOI21x1_ASAP7_75t_L g2915 ( 
.A1(n_2235),
.A2(n_2292),
.B(n_2284),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2284),
.B(n_2291),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2291),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2037),
.B(n_2028),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_1988),
.B(n_2034),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2037),
.B(n_2034),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2338),
.B(n_2309),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_1988),
.B(n_2034),
.Y(n_2922)
);

O2A1O1Ixp33_ASAP7_75t_L g2923 ( 
.A1(n_2127),
.A2(n_2290),
.B(n_2286),
.C(n_2199),
.Y(n_2923)
);

HB1xp67_ASAP7_75t_L g2924 ( 
.A(n_1957),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_SL g2925 ( 
.A1(n_2091),
.A2(n_2309),
.B1(n_2293),
.B2(n_2219),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_1911),
.Y(n_2926)
);

O2A1O1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_1970),
.A2(n_2012),
.B(n_1899),
.C(n_1898),
.Y(n_2927)
);

O2A1O1Ixp33_ASAP7_75t_L g2928 ( 
.A1(n_1970),
.A2(n_2012),
.B(n_1899),
.C(n_2034),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_2008),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2037),
.B(n_2004),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2091),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_1911),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_1988),
.B(n_2004),
.Y(n_2933)
);

AOI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_1970),
.A2(n_2012),
.B(n_1902),
.Y(n_2934)
);

O2A1O1Ixp33_ASAP7_75t_L g2935 ( 
.A1(n_1988),
.A2(n_2004),
.B(n_1957),
.C(n_2032),
.Y(n_2935)
);

INVx2_ASAP7_75t_SL g2936 ( 
.A(n_2008),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_1902),
.A2(n_1911),
.B(n_1931),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2004),
.B(n_1957),
.Y(n_2938)
);

CKINVDCx20_ASAP7_75t_R g2939 ( 
.A(n_2091),
.Y(n_2939)
);

OR2x2_ASAP7_75t_L g2940 ( 
.A(n_1902),
.B(n_1911),
.Y(n_2940)
);

OAI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_1902),
.A2(n_2032),
.B(n_2003),
.Y(n_2941)
);

OR2x6_ASAP7_75t_SL g2942 ( 
.A(n_2091),
.B(n_2116),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_1911),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2103),
.A2(n_2155),
.B1(n_2293),
.B2(n_2219),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_1931),
.B(n_1943),
.Y(n_2945)
);

O2A1O1Ixp33_ASAP7_75t_L g2946 ( 
.A1(n_2008),
.A2(n_2155),
.B(n_2293),
.C(n_2219),
.Y(n_2946)
);

CKINVDCx20_ASAP7_75t_R g2947 ( 
.A(n_2103),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_1931),
.A2(n_1943),
.B(n_2021),
.Y(n_2948)
);

AOI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_1931),
.A2(n_1943),
.B(n_2021),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_1931),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_1943),
.A2(n_2021),
.B(n_2194),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_1943),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2103),
.A2(n_2194),
.B1(n_2293),
.B2(n_2219),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_L g2954 ( 
.A(n_2008),
.B(n_2194),
.Y(n_2954)
);

AOI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2103),
.A2(n_2194),
.B1(n_2293),
.B2(n_2116),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_1943),
.A2(n_2021),
.B(n_2116),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2116),
.B(n_2309),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2021),
.A2(n_2309),
.B(n_2155),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2116),
.B(n_2155),
.Y(n_2959)
);

AOI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2021),
.A2(n_2116),
.B(n_2155),
.Y(n_2960)
);

NOR3xp33_ASAP7_75t_L g2961 ( 
.A(n_2155),
.B(n_2194),
.C(n_2204),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2194),
.B(n_2204),
.Y(n_2962)
);

AOI221xp5_ASAP7_75t_L g2963 ( 
.A1(n_2293),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.C(n_1433),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2204),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2204),
.B(n_2219),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2204),
.Y(n_2966)
);

NAND2x1_ASAP7_75t_L g2967 ( 
.A(n_2204),
.B(n_2219),
.Y(n_2967)
);

OAI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_1633),
.A2(n_1476),
.B(n_1505),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_1702),
.B(n_1433),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_1702),
.B(n_1433),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_1702),
.B(n_1433),
.Y(n_2971)
);

AOI21xp5_ASAP7_75t_L g2972 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_1631),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_1727),
.B(n_1679),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2341),
.A2(n_1433),
.B1(n_1458),
.B2(n_1457),
.Y(n_2975)
);

NOR2xp67_ASAP7_75t_L g2976 ( 
.A(n_1678),
.B(n_621),
.Y(n_2976)
);

INVxp67_ASAP7_75t_L g2977 ( 
.A(n_1644),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_1727),
.B(n_1679),
.Y(n_2978)
);

OAI22xp5_ASAP7_75t_L g2979 ( 
.A1(n_2334),
.A2(n_1433),
.B1(n_1458),
.B2(n_1457),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2980)
);

AOI21x1_ASAP7_75t_L g2981 ( 
.A1(n_1661),
.A2(n_1763),
.B(n_1800),
.Y(n_2981)
);

OAI21x1_ASAP7_75t_L g2982 ( 
.A1(n_1800),
.A2(n_1969),
.B(n_2026),
.Y(n_2982)
);

AOI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2983)
);

AOI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2984)
);

AO21x1_ASAP7_75t_L g2985 ( 
.A1(n_1633),
.A2(n_2177),
.B(n_2142),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_1702),
.B(n_1433),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_1702),
.B(n_1433),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_1702),
.B(n_1433),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2285),
.B(n_1572),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_2052),
.Y(n_2992)
);

BUFx3_ASAP7_75t_L g2993 ( 
.A(n_2013),
.Y(n_2993)
);

AOI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2994)
);

INVx4_ASAP7_75t_L g2995 ( 
.A(n_1811),
.Y(n_2995)
);

CKINVDCx10_ASAP7_75t_R g2996 ( 
.A(n_2124),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2334),
.A2(n_1433),
.B1(n_1458),
.B2(n_1457),
.Y(n_2997)
);

AOI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_2998)
);

INVxp67_ASAP7_75t_L g2999 ( 
.A(n_1644),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2195),
.B(n_1433),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2195),
.B(n_1433),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_1702),
.B(n_1433),
.Y(n_3002)
);

AOI21xp5_ASAP7_75t_L g3003 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_3003)
);

AOI21x1_ASAP7_75t_L g3004 ( 
.A1(n_1661),
.A2(n_1763),
.B(n_1800),
.Y(n_3004)
);

NOR2x1_ASAP7_75t_R g3005 ( 
.A(n_1759),
.B(n_463),
.Y(n_3005)
);

AO22x1_ASAP7_75t_L g3006 ( 
.A1(n_2171),
.A2(n_792),
.B1(n_1457),
.B2(n_1433),
.Y(n_3006)
);

O2A1O1Ixp33_ASAP7_75t_L g3007 ( 
.A1(n_2104),
.A2(n_1505),
.B(n_1557),
.C(n_1525),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_3008)
);

NOR3xp33_ASAP7_75t_L g3009 ( 
.A(n_2259),
.B(n_1525),
.C(n_1505),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_1628),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_1633),
.A2(n_1476),
.B(n_1505),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_1766),
.B(n_1629),
.Y(n_3012)
);

NOR3xp33_ASAP7_75t_L g3013 ( 
.A(n_2259),
.B(n_1525),
.C(n_1505),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_1702),
.B(n_1433),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_1702),
.B(n_1433),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_1702),
.B(n_1433),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_1631),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_1727),
.B(n_1679),
.Y(n_3018)
);

A2O1A1Ixp33_ASAP7_75t_L g3019 ( 
.A1(n_2142),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3019)
);

AOI21xp5_ASAP7_75t_L g3020 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_3020)
);

A2O1A1Ixp33_ASAP7_75t_L g3021 ( 
.A1(n_2142),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3021)
);

OR2x2_ASAP7_75t_L g3022 ( 
.A(n_1766),
.B(n_1629),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2195),
.B(n_1433),
.Y(n_3023)
);

BUFx8_ASAP7_75t_SL g3024 ( 
.A(n_1759),
.Y(n_3024)
);

OAI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2334),
.A2(n_1433),
.B1(n_1458),
.B2(n_1457),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_1702),
.B(n_1433),
.Y(n_3026)
);

INVx1_ASAP7_75t_SL g3027 ( 
.A(n_1680),
.Y(n_3027)
);

BUFx6f_ASAP7_75t_L g3028 ( 
.A(n_2123),
.Y(n_3028)
);

OR2x2_ASAP7_75t_L g3029 ( 
.A(n_1766),
.B(n_1629),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2195),
.B(n_1433),
.Y(n_3030)
);

BUFx12f_ASAP7_75t_L g3031 ( 
.A(n_1759),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_1800),
.A2(n_1145),
.B(n_1140),
.Y(n_3032)
);

AOI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2171),
.A2(n_1433),
.B1(n_1458),
.B2(n_1457),
.Y(n_3033)
);

NAND2x1p5_ASAP7_75t_L g3034 ( 
.A(n_1944),
.B(n_1811),
.Y(n_3034)
);

OR2x6_ASAP7_75t_L g3035 ( 
.A(n_1969),
.B(n_1823),
.Y(n_3035)
);

INVx3_ASAP7_75t_L g3036 ( 
.A(n_2726),
.Y(n_3036)
);

NAND2x1_ASAP7_75t_L g3037 ( 
.A(n_2520),
.B(n_2995),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2707),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2707),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3040)
);

BUFx12f_ASAP7_75t_L g3041 ( 
.A(n_2432),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2984),
.A2(n_2991),
.B(n_2987),
.Y(n_3043)
);

AOI221x1_ASAP7_75t_L g3044 ( 
.A1(n_3009),
.A2(n_3013),
.B1(n_2392),
.B2(n_3011),
.C(n_2968),
.Y(n_3044)
);

INVx1_ASAP7_75t_SL g3045 ( 
.A(n_2722),
.Y(n_3045)
);

AO31x2_ASAP7_75t_L g3046 ( 
.A1(n_2463),
.A2(n_2817),
.A3(n_2387),
.B(n_2574),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2348),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2994),
.A2(n_3003),
.B(n_2998),
.Y(n_3048)
);

INVx4_ASAP7_75t_L g3049 ( 
.A(n_2567),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3051)
);

INVx5_ASAP7_75t_L g3052 ( 
.A(n_3035),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2729),
.Y(n_3053)
);

AOI21xp33_ASAP7_75t_L g3054 ( 
.A1(n_3007),
.A2(n_3011),
.B(n_2968),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_2344),
.B(n_2403),
.Y(n_3055)
);

AOI21x1_ASAP7_75t_L g3056 ( 
.A1(n_2981),
.A2(n_3004),
.B(n_2421),
.Y(n_3056)
);

OAI21x1_ASAP7_75t_SL g3057 ( 
.A1(n_2491),
.A2(n_2365),
.B(n_2395),
.Y(n_3057)
);

OR2x6_ASAP7_75t_L g3058 ( 
.A(n_2417),
.B(n_3035),
.Y(n_3058)
);

BUFx4_ASAP7_75t_R g3059 ( 
.A(n_3024),
.Y(n_3059)
);

OAI21x1_ASAP7_75t_L g3060 ( 
.A1(n_2903),
.A2(n_2535),
.B(n_2523),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2729),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2736),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_3008),
.A2(n_3032),
.B(n_3020),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2608),
.Y(n_3064)
);

BUFx8_ASAP7_75t_L g3065 ( 
.A(n_2541),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2445),
.B(n_2356),
.Y(n_3066)
);

OAI21x1_ASAP7_75t_L g3067 ( 
.A1(n_2558),
.A2(n_2568),
.B(n_2564),
.Y(n_3067)
);

NAND2x1p5_ASAP7_75t_L g3068 ( 
.A(n_2451),
.B(n_2386),
.Y(n_3068)
);

OAI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2343),
.A2(n_2372),
.B(n_3019),
.Y(n_3069)
);

INVx3_ASAP7_75t_L g3070 ( 
.A(n_2608),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2353),
.B(n_2357),
.Y(n_3071)
);

OAI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2343),
.A2(n_3021),
.B(n_2354),
.Y(n_3072)
);

AOI21xp5_ASAP7_75t_L g3073 ( 
.A1(n_2360),
.A2(n_2440),
.B(n_2425),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2348),
.Y(n_3074)
);

A2O1A1Ixp33_ASAP7_75t_L g3075 ( 
.A1(n_2368),
.A2(n_2351),
.B(n_2346),
.C(n_2354),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2353),
.B(n_2357),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2942),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2377),
.A2(n_2418),
.B(n_2450),
.Y(n_3078)
);

AO31x2_ASAP7_75t_L g3079 ( 
.A1(n_2817),
.A2(n_2574),
.A3(n_2985),
.B(n_2358),
.Y(n_3079)
);

INVxp67_ASAP7_75t_SL g3080 ( 
.A(n_2345),
.Y(n_3080)
);

AOI221xp5_ASAP7_75t_L g3081 ( 
.A1(n_2368),
.A2(n_2975),
.B1(n_2979),
.B2(n_3025),
.C(n_2997),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2479),
.B(n_2625),
.Y(n_3082)
);

OAI21x1_ASAP7_75t_L g3083 ( 
.A1(n_2875),
.A2(n_2886),
.B(n_2553),
.Y(n_3083)
);

A2O1A1Ixp33_ASAP7_75t_L g3084 ( 
.A1(n_3000),
.A2(n_3001),
.B(n_3030),
.C(n_3023),
.Y(n_3084)
);

OAI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_3033),
.A2(n_2969),
.B1(n_2971),
.B2(n_2970),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2736),
.Y(n_3086)
);

A2O1A1Ixp33_ASAP7_75t_L g3087 ( 
.A1(n_3033),
.A2(n_2398),
.B(n_2422),
.C(n_2401),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2479),
.B(n_2625),
.Y(n_3088)
);

A2O1A1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_2422),
.A2(n_2397),
.B(n_2416),
.C(n_2411),
.Y(n_3089)
);

AO31x2_ASAP7_75t_L g3090 ( 
.A1(n_2358),
.A2(n_2985),
.A3(n_2464),
.B(n_2517),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2974),
.B(n_2978),
.Y(n_3091)
);

AO31x2_ASAP7_75t_L g3092 ( 
.A1(n_2517),
.A2(n_2454),
.A3(n_2539),
.B(n_2548),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_2531),
.A2(n_2570),
.B(n_2838),
.Y(n_3093)
);

OAI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2531),
.A2(n_2570),
.B(n_2850),
.Y(n_3094)
);

INVx3_ASAP7_75t_L g3095 ( 
.A(n_2600),
.Y(n_3095)
);

NOR2x1_ASAP7_75t_SL g3096 ( 
.A(n_2417),
.B(n_3035),
.Y(n_3096)
);

O2A1O1Ixp5_ASAP7_75t_L g3097 ( 
.A1(n_3006),
.A2(n_2373),
.B(n_2990),
.C(n_2406),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2583),
.B(n_2618),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2419),
.B(n_2544),
.Y(n_3099)
);

AOI21x1_ASAP7_75t_L g3100 ( 
.A1(n_2421),
.A2(n_2389),
.B(n_2394),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2584),
.A2(n_2373),
.B(n_2631),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2544),
.B(n_2376),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2830),
.Y(n_3103)
);

NOR2x1_ASAP7_75t_SL g3104 ( 
.A(n_2417),
.B(n_3035),
.Y(n_3104)
);

OAI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2518),
.A2(n_2386),
.B(n_3025),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2600),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2376),
.B(n_2383),
.Y(n_3107)
);

AOI21x1_ASAP7_75t_L g3108 ( 
.A1(n_2394),
.A2(n_2527),
.B(n_2459),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_SL g3109 ( 
.A(n_2963),
.B(n_2979),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2571),
.A2(n_2581),
.B(n_2575),
.Y(n_3110)
);

AOI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2465),
.A2(n_2451),
.B(n_2508),
.Y(n_3111)
);

OAI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2997),
.A2(n_2406),
.B(n_2347),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2383),
.B(n_2452),
.Y(n_3113)
);

OAI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_2414),
.A2(n_2452),
.B(n_2976),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2509),
.A2(n_2489),
.B(n_2460),
.Y(n_3115)
);

INVxp67_ASAP7_75t_L g3116 ( 
.A(n_2617),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2460),
.A2(n_2557),
.B(n_2510),
.Y(n_3117)
);

OAI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2986),
.A2(n_2989),
.B1(n_3002),
.B2(n_2988),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_SL g3119 ( 
.A1(n_2946),
.A2(n_2756),
.B(n_2754),
.Y(n_3119)
);

INVxp67_ASAP7_75t_SL g3120 ( 
.A(n_2640),
.Y(n_3120)
);

OAI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2976),
.A2(n_2428),
.B(n_2530),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2557),
.A2(n_3006),
.B(n_2602),
.Y(n_3122)
);

O2A1O1Ixp5_ASAP7_75t_L g3123 ( 
.A1(n_2519),
.A2(n_2540),
.B(n_2526),
.C(n_2539),
.Y(n_3123)
);

A2O1A1Ixp33_ASAP7_75t_L g3124 ( 
.A1(n_2435),
.A2(n_2530),
.B(n_2514),
.C(n_2441),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2499),
.A2(n_2500),
.B(n_2417),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2974),
.B(n_2978),
.Y(n_3126)
);

INVx3_ASAP7_75t_L g3127 ( 
.A(n_2520),
.Y(n_3127)
);

NAND3xp33_ASAP7_75t_L g3128 ( 
.A(n_2423),
.B(n_2433),
.C(n_2367),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2442),
.B(n_2443),
.Y(n_3129)
);

OAI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_3014),
.A2(n_3016),
.B1(n_3015),
.B2(n_3026),
.Y(n_3130)
);

OAI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2537),
.A2(n_2390),
.B(n_2355),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2830),
.Y(n_3132)
);

AOI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_3035),
.A2(n_2498),
.B(n_2492),
.Y(n_3133)
);

BUFx4f_ASAP7_75t_L g3134 ( 
.A(n_2567),
.Y(n_3134)
);

OA21x2_ASAP7_75t_L g3135 ( 
.A1(n_2536),
.A2(n_2802),
.B(n_2580),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2639),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_3018),
.B(n_2458),
.Y(n_3137)
);

OAI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2413),
.A2(n_2471),
.B(n_2410),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2635),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2456),
.B(n_2478),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2522),
.B(n_2349),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2635),
.Y(n_3142)
);

AO31x2_ASAP7_75t_L g3143 ( 
.A1(n_2616),
.A2(n_2889),
.A3(n_2613),
.B(n_2913),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2639),
.Y(n_3144)
);

BUFx2_ASAP7_75t_L g3145 ( 
.A(n_2696),
.Y(n_3145)
);

AOI21x1_ASAP7_75t_L g3146 ( 
.A1(n_2527),
.A2(n_2597),
.B(n_2675),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2495),
.B(n_2620),
.Y(n_3147)
);

AOI21x1_ASAP7_75t_L g3148 ( 
.A1(n_2599),
.A2(n_2693),
.B(n_2695),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_3018),
.B(n_2458),
.Y(n_3149)
);

A2O1A1Ixp33_ASAP7_75t_L g3150 ( 
.A1(n_2514),
.A2(n_2441),
.B(n_2404),
.C(n_2410),
.Y(n_3150)
);

BUFx8_ASAP7_75t_L g3151 ( 
.A(n_2541),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2350),
.B(n_2352),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2620),
.B(n_2511),
.Y(n_3153)
);

AOI21x1_ASAP7_75t_L g3154 ( 
.A1(n_2585),
.A2(n_2845),
.B(n_2697),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_2536),
.A2(n_2827),
.B(n_2848),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2515),
.B(n_2455),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2560),
.B(n_2493),
.Y(n_3157)
);

OAI21x1_ASAP7_75t_L g3158 ( 
.A1(n_2627),
.A2(n_2629),
.B(n_3034),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2455),
.B(n_2483),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2483),
.B(n_2477),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2776),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2681),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2462),
.A2(n_2505),
.B(n_2497),
.Y(n_3163)
);

AO31x2_ASAP7_75t_L g3164 ( 
.A1(n_2889),
.A2(n_2913),
.A3(n_2660),
.B(n_2519),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2477),
.B(n_2404),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2560),
.B(n_2493),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2361),
.B(n_3012),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2653),
.Y(n_3168)
);

CKINVDCx5p33_ASAP7_75t_R g3169 ( 
.A(n_2653),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2703),
.A2(n_2705),
.B(n_2739),
.Y(n_3170)
);

OR2x2_ASAP7_75t_L g3171 ( 
.A(n_2361),
.B(n_3012),
.Y(n_3171)
);

O2A1O1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_2522),
.A2(n_2633),
.B(n_2481),
.C(n_2490),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_3022),
.B(n_3029),
.Y(n_3173)
);

A2O1A1Ixp33_ASAP7_75t_L g3174 ( 
.A1(n_2470),
.A2(n_2494),
.B(n_2525),
.C(n_2580),
.Y(n_3174)
);

O2A1O1Ixp5_ASAP7_75t_L g3175 ( 
.A1(n_2554),
.A2(n_2552),
.B(n_2696),
.C(n_2662),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3022),
.B(n_3029),
.Y(n_3176)
);

OAI21x1_ASAP7_75t_L g3177 ( 
.A1(n_2682),
.A2(n_2898),
.B(n_2689),
.Y(n_3177)
);

OR2x6_ASAP7_75t_L g3178 ( 
.A(n_2656),
.B(n_2663),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2789),
.Y(n_3179)
);

OAI21x1_ASAP7_75t_SL g3180 ( 
.A1(n_2641),
.A2(n_2590),
.B(n_2589),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2638),
.B(n_2506),
.Y(n_3181)
);

AOI31xp33_ASAP7_75t_SL g3182 ( 
.A1(n_2482),
.A2(n_2566),
.A3(n_2810),
.B(n_2446),
.Y(n_3182)
);

OAI22xp5_ASAP7_75t_L g3183 ( 
.A1(n_2429),
.A2(n_2369),
.B1(n_2374),
.B2(n_2363),
.Y(n_3183)
);

BUFx4_ASAP7_75t_SL g3184 ( 
.A(n_2773),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2506),
.B(n_2601),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2789),
.Y(n_3186)
);

NAND2x1p5_ASAP7_75t_L g3187 ( 
.A(n_2520),
.B(n_2995),
.Y(n_3187)
);

O2A1O1Ixp5_ASAP7_75t_L g3188 ( 
.A1(n_2751),
.A2(n_2582),
.B(n_2802),
.C(n_2621),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2601),
.B(n_2375),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2855),
.A2(n_2674),
.B(n_2426),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2674),
.A2(n_2426),
.B(n_2567),
.Y(n_3191)
);

BUFx2_ASAP7_75t_L g3192 ( 
.A(n_2503),
.Y(n_3192)
);

OAI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2775),
.A2(n_2476),
.B(n_2446),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2378),
.B(n_2379),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2380),
.B(n_2385),
.Y(n_3195)
);

INVx4_ASAP7_75t_L g3196 ( 
.A(n_2652),
.Y(n_3196)
);

OAI21x1_ASAP7_75t_L g3197 ( 
.A1(n_2713),
.A2(n_2723),
.B(n_2716),
.Y(n_3197)
);

BUFx3_ASAP7_75t_L g3198 ( 
.A(n_2942),
.Y(n_3198)
);

OAI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_2429),
.A2(n_2391),
.B1(n_2399),
.B2(n_2393),
.Y(n_3199)
);

OAI21x1_ASAP7_75t_L g3200 ( 
.A1(n_2733),
.A2(n_2833),
.B(n_2738),
.Y(n_3200)
);

AO31x2_ASAP7_75t_L g3201 ( 
.A1(n_2503),
.A2(n_2598),
.A3(n_2724),
.B(n_2587),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2582),
.B(n_2549),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2728),
.B(n_2734),
.Y(n_3203)
);

BUFx3_ASAP7_75t_L g3204 ( 
.A(n_2667),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2415),
.Y(n_3205)
);

AOI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_2778),
.A2(n_2822),
.B(n_2765),
.Y(n_3206)
);

OAI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_2405),
.A2(n_2412),
.B1(n_2447),
.B2(n_2431),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2448),
.B(n_2449),
.Y(n_3208)
);

OAI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_2467),
.A2(n_2472),
.B1(n_2473),
.B2(n_2469),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2765),
.A2(n_2829),
.B(n_2883),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2439),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2475),
.B(n_2486),
.Y(n_3212)
);

NOR2xp33_ASAP7_75t_L g3213 ( 
.A(n_2496),
.B(n_2342),
.Y(n_3213)
);

NAND2xp33_ASAP7_75t_SL g3214 ( 
.A(n_2882),
.B(n_2902),
.Y(n_3214)
);

OAI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2446),
.A2(n_2710),
.B(n_2549),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2520),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2439),
.Y(n_3217)
);

NAND3xp33_ASAP7_75t_L g3218 ( 
.A(n_2642),
.B(n_2658),
.C(n_2566),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_2596),
.A2(n_2610),
.B(n_2609),
.Y(n_3219)
);

AOI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_2468),
.A2(n_2642),
.B1(n_2550),
.B2(n_2496),
.Y(n_3220)
);

NAND3xp33_ASAP7_75t_SL g3221 ( 
.A(n_2717),
.B(n_2603),
.C(n_2759),
.Y(n_3221)
);

A2O1A1Ixp33_ASAP7_75t_L g3222 ( 
.A1(n_2686),
.A2(n_2710),
.B(n_2766),
.C(n_2825),
.Y(n_3222)
);

A2O1A1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_2686),
.A2(n_2825),
.B(n_2732),
.C(n_2735),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_2871),
.A2(n_2901),
.B(n_2892),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2487),
.B(n_2630),
.Y(n_3225)
);

OAI21x1_ASAP7_75t_L g3226 ( 
.A1(n_2637),
.A2(n_2763),
.B(n_2738),
.Y(n_3226)
);

OAI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_2814),
.A2(n_2821),
.B(n_2590),
.Y(n_3227)
);

AND2x4_ASAP7_75t_L g3228 ( 
.A(n_2344),
.B(n_2403),
.Y(n_3228)
);

AOI21x1_ASAP7_75t_L g3229 ( 
.A1(n_2845),
.A2(n_2949),
.B(n_2948),
.Y(n_3229)
);

OR2x6_ASAP7_75t_L g3230 ( 
.A(n_2724),
.B(n_2579),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2521),
.B(n_2702),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_2837),
.A2(n_2923),
.B(n_2910),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2702),
.B(n_2720),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2856),
.A2(n_2894),
.B(n_2869),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_2415),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_2995),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_2728),
.B(n_2734),
.Y(n_3237)
);

BUFx2_ASAP7_75t_L g3238 ( 
.A(n_2661),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2720),
.B(n_2741),
.Y(n_3239)
);

AOI221x1_ASAP7_75t_L g3240 ( 
.A1(n_2687),
.A2(n_2651),
.B1(n_2750),
.B2(n_2694),
.C(n_2961),
.Y(n_3240)
);

AND2x2_ASAP7_75t_SL g3241 ( 
.A(n_2800),
.B(n_2815),
.Y(n_3241)
);

NAND2x1_ASAP7_75t_L g3242 ( 
.A(n_2995),
.B(n_2652),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2741),
.B(n_2744),
.Y(n_3243)
);

OR2x6_ASAP7_75t_L g3244 ( 
.A(n_2579),
.B(n_2344),
.Y(n_3244)
);

OAI21x1_ASAP7_75t_L g3245 ( 
.A1(n_2837),
.A2(n_2881),
.B(n_2842),
.Y(n_3245)
);

OAI21x1_ASAP7_75t_SL g3246 ( 
.A1(n_2927),
.A2(n_2813),
.B(n_2928),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2790),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_2760),
.A2(n_2786),
.B(n_2774),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2744),
.B(n_2555),
.Y(n_3249)
);

CKINVDCx5p33_ASAP7_75t_R g3250 ( 
.A(n_2654),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2790),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2555),
.B(n_2661),
.Y(n_3252)
);

OR2x6_ASAP7_75t_L g3253 ( 
.A(n_2579),
.B(n_2344),
.Y(n_3253)
);

OAI21x1_ASAP7_75t_L g3254 ( 
.A1(n_2837),
.A2(n_2881),
.B(n_2842),
.Y(n_3254)
);

OAI21x1_ASAP7_75t_L g3255 ( 
.A1(n_2753),
.A2(n_2937),
.B(n_2900),
.Y(n_3255)
);

AND3x2_ASAP7_75t_L g3256 ( 
.A(n_2752),
.B(n_2876),
.C(n_2742),
.Y(n_3256)
);

OAI21x1_ASAP7_75t_L g3257 ( 
.A1(n_2753),
.A2(n_2900),
.B(n_2801),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2645),
.B(n_2668),
.Y(n_3258)
);

OAI21x1_ASAP7_75t_L g3259 ( 
.A1(n_2801),
.A2(n_2900),
.B(n_2897),
.Y(n_3259)
);

NOR2xp67_ASAP7_75t_L g3260 ( 
.A(n_2755),
.B(n_2777),
.Y(n_3260)
);

NAND3xp33_ASAP7_75t_L g3261 ( 
.A(n_2634),
.B(n_2659),
.C(n_2619),
.Y(n_3261)
);

OAI21x1_ASAP7_75t_L g3262 ( 
.A1(n_2801),
.A2(n_2904),
.B(n_2897),
.Y(n_3262)
);

OAI21x1_ASAP7_75t_L g3263 ( 
.A1(n_2897),
.A2(n_2908),
.B(n_2904),
.Y(n_3263)
);

OAI21x1_ASAP7_75t_L g3264 ( 
.A1(n_2897),
.A2(n_2908),
.B(n_2904),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_2496),
.A2(n_2808),
.B(n_2788),
.Y(n_3265)
);

OAI21x1_ASAP7_75t_L g3266 ( 
.A1(n_2904),
.A2(n_2908),
.B(n_2951),
.Y(n_3266)
);

INVxp67_ASAP7_75t_L g3267 ( 
.A(n_2364),
.Y(n_3267)
);

AOI21x1_ASAP7_75t_L g3268 ( 
.A1(n_2761),
.A2(n_2770),
.B(n_2762),
.Y(n_3268)
);

OAI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_2782),
.A2(n_2891),
.B(n_2809),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_2958),
.A2(n_2960),
.B(n_2755),
.Y(n_3270)
);

BUFx3_ASAP7_75t_L g3271 ( 
.A(n_2667),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_2956),
.A2(n_2852),
.B(n_2698),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_2712),
.B(n_2730),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_2852),
.A2(n_2704),
.B(n_2683),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2852),
.A2(n_2725),
.B(n_2709),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_2852),
.A2(n_2849),
.B(n_2806),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_2852),
.A2(n_2797),
.B(n_2803),
.Y(n_3277)
);

INVx1_ASAP7_75t_SL g3278 ( 
.A(n_2722),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2819),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2439),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_2444),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2819),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2645),
.B(n_2668),
.Y(n_3283)
);

INVxp67_ASAP7_75t_L g3284 ( 
.A(n_2644),
.Y(n_3284)
);

AO31x2_ASAP7_75t_L g3285 ( 
.A1(n_2757),
.A2(n_2771),
.A3(n_2824),
.B(n_2812),
.Y(n_3285)
);

AOI221xp5_ASAP7_75t_L g3286 ( 
.A1(n_2592),
.A2(n_2561),
.B1(n_2562),
.B2(n_2538),
.C(n_2532),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2706),
.B(n_2916),
.Y(n_3287)
);

HB1xp67_ASAP7_75t_L g3288 ( 
.A(n_2591),
.Y(n_3288)
);

OAI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2468),
.A2(n_2586),
.B1(n_2573),
.B2(n_2577),
.Y(n_3289)
);

NOR2xp67_ASAP7_75t_L g3290 ( 
.A(n_2777),
.B(n_2792),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2444),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2834),
.Y(n_3292)
);

BUFx2_ASAP7_75t_L g3293 ( 
.A(n_2371),
.Y(n_3293)
);

AND2x4_ASAP7_75t_L g3294 ( 
.A(n_2403),
.B(n_2794),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2796),
.A2(n_2559),
.B(n_2524),
.Y(n_3295)
);

A2O1A1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_2811),
.A2(n_2769),
.B(n_2820),
.C(n_2941),
.Y(n_3296)
);

OAI21x1_ASAP7_75t_SL g3297 ( 
.A1(n_2935),
.A2(n_2941),
.B(n_2859),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2706),
.B(n_2916),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2444),
.B(n_2973),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2973),
.B(n_3017),
.Y(n_3300)
);

AO21x2_ASAP7_75t_L g3301 ( 
.A1(n_2891),
.A2(n_2859),
.B(n_2847),
.Y(n_3301)
);

INVx3_ASAP7_75t_L g3302 ( 
.A(n_2359),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_2480),
.B(n_2488),
.Y(n_3303)
);

INVx8_ASAP7_75t_L g3304 ( 
.A(n_2667),
.Y(n_3304)
);

AOI21xp33_ASAP7_75t_L g3305 ( 
.A1(n_2468),
.A2(n_2594),
.B(n_2793),
.Y(n_3305)
);

A2O1A1Ixp33_ASAP7_75t_L g3306 ( 
.A1(n_2811),
.A2(n_2820),
.B(n_2791),
.C(n_2700),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2973),
.B(n_3017),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_2359),
.Y(n_3308)
);

AOI21x1_ASAP7_75t_L g3309 ( 
.A1(n_2651),
.A2(n_2750),
.B(n_2694),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2847),
.A2(n_2861),
.B(n_2860),
.Y(n_3310)
);

BUFx12f_ASAP7_75t_L g3311 ( 
.A(n_2432),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2524),
.A2(n_2873),
.B(n_2559),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_2524),
.A2(n_2873),
.B(n_2559),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_2873),
.A2(n_2805),
.B(n_2665),
.Y(n_3314)
);

AO21x2_ASAP7_75t_L g3315 ( 
.A1(n_2860),
.A2(n_2861),
.B(n_2780),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3017),
.B(n_2746),
.Y(n_3316)
);

AOI21x1_ASAP7_75t_L g3317 ( 
.A1(n_2911),
.A2(n_2957),
.B(n_2921),
.Y(n_3317)
);

AOI21xp33_ASAP7_75t_L g3318 ( 
.A1(n_2749),
.A2(n_3027),
.B(n_2569),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2381),
.B(n_2384),
.Y(n_3319)
);

INVx4_ASAP7_75t_L g3320 ( 
.A(n_2652),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_2652),
.A2(n_2840),
.B(n_2665),
.Y(n_3321)
);

HB1xp67_ASAP7_75t_L g3322 ( 
.A(n_2591),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2737),
.Y(n_3323)
);

OAI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_2823),
.A2(n_2877),
.B(n_2578),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_2665),
.A2(n_2840),
.B(n_2962),
.Y(n_3325)
);

BUFx10_ASAP7_75t_L g3326 ( 
.A(n_2541),
.Y(n_3326)
);

OAI21x1_ASAP7_75t_L g3327 ( 
.A1(n_2436),
.A2(n_2614),
.B(n_2547),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2665),
.A2(n_2840),
.B(n_2918),
.Y(n_3328)
);

HB1xp67_ASAP7_75t_L g3329 ( 
.A(n_2636),
.Y(n_3329)
);

AOI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_2840),
.A2(n_2678),
.B(n_2605),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_2678),
.A2(n_2605),
.B(n_2542),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_2542),
.A2(n_2815),
.B(n_2800),
.Y(n_3332)
);

BUFx6f_ASAP7_75t_L g3333 ( 
.A(n_2800),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_2815),
.A2(n_2843),
.B(n_2912),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_2712),
.B(n_2569),
.Y(n_3335)
);

OAI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_2572),
.A2(n_2909),
.B1(n_3027),
.B2(n_2556),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3010),
.B(n_2835),
.Y(n_3337)
);

A2O1A1Ixp33_ASAP7_75t_L g3338 ( 
.A1(n_2876),
.A2(n_2890),
.B(n_2669),
.C(n_2671),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3010),
.B(n_2835),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_2480),
.B(n_2488),
.Y(n_3340)
);

CKINVDCx20_ASAP7_75t_R g3341 ( 
.A(n_2507),
.Y(n_3341)
);

NAND2x1p5_ASAP7_75t_L g3342 ( 
.A(n_2721),
.B(n_2912),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_L g3343 ( 
.A(n_2342),
.B(n_2623),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2839),
.B(n_2844),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2839),
.B(n_2844),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_2768),
.B(n_2785),
.Y(n_3346)
);

OAI21x1_ASAP7_75t_L g3347 ( 
.A1(n_2846),
.A2(n_2857),
.B(n_2851),
.Y(n_3347)
);

INVx1_ASAP7_75t_SL g3348 ( 
.A(n_2899),
.Y(n_3348)
);

A2O1A1Ixp33_ASAP7_75t_L g3349 ( 
.A1(n_2831),
.A2(n_2721),
.B(n_2864),
.C(n_2832),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2768),
.B(n_2785),
.Y(n_3350)
);

O2A1O1Ixp5_ASAP7_75t_L g3351 ( 
.A1(n_2622),
.A2(n_2657),
.B(n_2666),
.C(n_2836),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2868),
.A2(n_2878),
.B(n_2870),
.Y(n_3352)
);

OAI21x1_ASAP7_75t_L g3353 ( 
.A1(n_2884),
.A2(n_2893),
.B(n_2885),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_2758),
.B(n_2945),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_2895),
.A2(n_2907),
.B(n_2896),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2388),
.Y(n_3356)
);

AO31x2_ASAP7_75t_L g3357 ( 
.A1(n_2474),
.A2(n_2533),
.A3(n_2543),
.B(n_2484),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_2400),
.B(n_2402),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_SL g3359 ( 
.A1(n_2382),
.A2(n_2453),
.B(n_2437),
.Y(n_3359)
);

AO21x1_ASAP7_75t_L g3360 ( 
.A1(n_2783),
.A2(n_2784),
.B(n_2779),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_2474),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2400),
.Y(n_3362)
);

AOI21x1_ASAP7_75t_L g3363 ( 
.A1(n_2781),
.A2(n_2807),
.B(n_2798),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2420),
.B(n_2424),
.Y(n_3364)
);

CKINVDCx5p33_ASAP7_75t_R g3365 ( 
.A(n_2654),
.Y(n_3365)
);

AND2x6_ASAP7_75t_L g3366 ( 
.A(n_2382),
.B(n_2437),
.Y(n_3366)
);

NAND2x1p5_ASAP7_75t_L g3367 ( 
.A(n_2912),
.B(n_2944),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_2420),
.B(n_2424),
.Y(n_3368)
);

OAI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_2934),
.A2(n_2879),
.B(n_2798),
.Y(n_3369)
);

AOI21x1_ASAP7_75t_L g3370 ( 
.A1(n_2781),
.A2(n_2807),
.B(n_2799),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2474),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_2758),
.B(n_2507),
.Y(n_3372)
);

NAND2x1p5_ASAP7_75t_L g3373 ( 
.A(n_2912),
.B(n_2944),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2438),
.B(n_2457),
.Y(n_3374)
);

OAI21xp33_ASAP7_75t_L g3375 ( 
.A1(n_2606),
.A2(n_2643),
.B(n_2408),
.Y(n_3375)
);

AO31x2_ASAP7_75t_L g3376 ( 
.A1(n_2533),
.A2(n_2563),
.A3(n_2680),
.B(n_2747),
.Y(n_3376)
);

INVxp67_ASAP7_75t_L g3377 ( 
.A(n_2626),
.Y(n_3377)
);

INVx2_ASAP7_75t_SL g3378 ( 
.A(n_2415),
.Y(n_3378)
);

INVx4_ASAP7_75t_L g3379 ( 
.A(n_2382),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_2758),
.B(n_2407),
.Y(n_3380)
);

OAI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_2690),
.A2(n_2692),
.B(n_2920),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_2912),
.A2(n_2865),
.B(n_2758),
.Y(n_3382)
);

OAI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_2930),
.A2(n_2745),
.B(n_2743),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_2912),
.A2(n_2865),
.B(n_2953),
.Y(n_3384)
);

OAI222xp33_ASAP7_75t_L g3385 ( 
.A1(n_2748),
.A2(n_2759),
.B1(n_2512),
.B2(n_2999),
.C1(n_2565),
.C2(n_2977),
.Y(n_3385)
);

NOR2x1_ASAP7_75t_L g3386 ( 
.A(n_2461),
.B(n_2551),
.Y(n_3386)
);

A2O1A1Ixp33_ASAP7_75t_L g3387 ( 
.A1(n_2831),
.A2(n_2953),
.B(n_2955),
.C(n_2816),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_2909),
.A2(n_2939),
.B1(n_2947),
.B2(n_2529),
.Y(n_3388)
);

AOI21x1_ASAP7_75t_L g3389 ( 
.A1(n_2863),
.A2(n_2943),
.B(n_2926),
.Y(n_3389)
);

NOR2xp67_ASAP7_75t_L g3390 ( 
.A(n_2955),
.B(n_2964),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_2593),
.B(n_2636),
.Y(n_3391)
);

A2O1A1Ixp33_ASAP7_75t_L g3392 ( 
.A1(n_2816),
.A2(n_2826),
.B(n_2461),
.C(n_2804),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_2945),
.B(n_2888),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_SL g3394 ( 
.A(n_2670),
.B(n_2672),
.Y(n_3394)
);

INVx3_ASAP7_75t_L g3395 ( 
.A(n_2632),
.Y(n_3395)
);

OAI22xp5_ASAP7_75t_L g3396 ( 
.A1(n_2914),
.A2(n_2366),
.B1(n_2993),
.B2(n_2925),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2865),
.A2(n_2731),
.B(n_2673),
.Y(n_3397)
);

INVx3_ASAP7_75t_L g3398 ( 
.A(n_2650),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2502),
.B(n_2504),
.Y(n_3399)
);

INVx4_ASAP7_75t_L g3400 ( 
.A(n_2382),
.Y(n_3400)
);

OAI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_2933),
.A2(n_2919),
.B(n_2922),
.Y(n_3401)
);

AO31x2_ASAP7_75t_L g3402 ( 
.A1(n_2650),
.A2(n_2767),
.A3(n_2685),
.B(n_2714),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_SL g3403 ( 
.A1(n_2382),
.A2(n_2528),
.B(n_3028),
.Y(n_3403)
);

AOI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_2396),
.A2(n_3031),
.B1(n_2604),
.B2(n_2534),
.Y(n_3404)
);

OAI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_2938),
.A2(n_2866),
.B(n_2854),
.Y(n_3405)
);

O2A1O1Ixp5_ASAP7_75t_L g3406 ( 
.A1(n_2964),
.A2(n_2967),
.B(n_2932),
.C(n_2952),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2504),
.B(n_2516),
.Y(n_3407)
);

OAI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_2854),
.A2(n_2866),
.B(n_2880),
.Y(n_3408)
);

NOR3xp33_ASAP7_75t_L g3409 ( 
.A(n_3005),
.B(n_2546),
.C(n_2764),
.Y(n_3409)
);

OAI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_2914),
.A2(n_2366),
.B1(n_2993),
.B2(n_2784),
.Y(n_3410)
);

NOR2x1_ASAP7_75t_L g3411 ( 
.A(n_2551),
.B(n_2865),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_2676),
.B(n_2677),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_2865),
.A2(n_2740),
.B(n_2679),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_2888),
.B(n_2932),
.Y(n_3414)
);

OAI22xp5_ASAP7_75t_L g3415 ( 
.A1(n_2366),
.A2(n_2993),
.B1(n_2779),
.B2(n_2795),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_2684),
.A2(n_2727),
.B(n_2688),
.Y(n_3416)
);

INVx2_ASAP7_75t_SL g3417 ( 
.A(n_2551),
.Y(n_3417)
);

HB1xp67_ASAP7_75t_L g3418 ( 
.A(n_2899),
.Y(n_3418)
);

AOI21xp33_ASAP7_75t_L g3419 ( 
.A1(n_2371),
.A2(n_2434),
.B(n_2612),
.Y(n_3419)
);

AO31x2_ASAP7_75t_L g3420 ( 
.A1(n_2767),
.A2(n_2787),
.A3(n_2917),
.B(n_2874),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_2787),
.Y(n_3421)
);

AO21x2_ASAP7_75t_L g3422 ( 
.A1(n_2545),
.A2(n_2607),
.B(n_2648),
.Y(n_3422)
);

BUFx2_ASAP7_75t_L g3423 ( 
.A(n_2434),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_2699),
.B(n_2701),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_2950),
.B(n_2952),
.Y(n_3425)
);

NAND2x1p5_ASAP7_75t_L g3426 ( 
.A(n_2967),
.B(n_2437),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_2711),
.A2(n_2719),
.B(n_2466),
.Y(n_3427)
);

NAND2x1p5_ASAP7_75t_L g3428 ( 
.A(n_2437),
.B(n_2453),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_2576),
.B(n_2612),
.Y(n_3429)
);

AOI21xp33_ASAP7_75t_L g3430 ( 
.A1(n_2615),
.A2(n_2715),
.B(n_2648),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_2437),
.A2(n_2513),
.B(n_2595),
.Y(n_3431)
);

NOR2x1_ASAP7_75t_L g3432 ( 
.A(n_2940),
.B(n_2858),
.Y(n_3432)
);

NOR2x1_ASAP7_75t_SL g3433 ( 
.A(n_2453),
.B(n_2513),
.Y(n_3433)
);

INVx2_ASAP7_75t_SL g3434 ( 
.A(n_2818),
.Y(n_3434)
);

INVx8_ASAP7_75t_L g3435 ( 
.A(n_2667),
.Y(n_3435)
);

AO31x2_ASAP7_75t_L g3436 ( 
.A1(n_2862),
.A2(n_2872),
.A3(n_2628),
.B(n_2715),
.Y(n_3436)
);

A2O1A1Ixp33_ASAP7_75t_L g3437 ( 
.A1(n_2959),
.A2(n_2954),
.B(n_2867),
.C(n_2624),
.Y(n_3437)
);

NAND2x1_ASAP7_75t_L g3438 ( 
.A(n_2667),
.B(n_2950),
.Y(n_3438)
);

NOR3xp33_ASAP7_75t_L g3439 ( 
.A(n_3005),
.B(n_2546),
.C(n_2664),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2841),
.B(n_2887),
.Y(n_3440)
);

OAI21x1_ASAP7_75t_L g3441 ( 
.A1(n_2841),
.A2(n_2906),
.B(n_2905),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_2453),
.A2(n_2528),
.B(n_2595),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2905),
.B(n_2924),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2940),
.B(n_2867),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_2453),
.A2(n_2501),
.B(n_2624),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_2867),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2965),
.B(n_2929),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_2965),
.B(n_2929),
.Y(n_3448)
);

OAI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_2936),
.A2(n_2611),
.B(n_2992),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_2646),
.B(n_2655),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_2646),
.B(n_2655),
.Y(n_3451)
);

OAI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_2992),
.A2(n_2795),
.B(n_2501),
.Y(n_3452)
);

NAND3xp33_ASAP7_75t_L g3453 ( 
.A(n_2432),
.B(n_2624),
.C(n_2595),
.Y(n_3453)
);

OA21x2_ASAP7_75t_L g3454 ( 
.A1(n_2646),
.A2(n_2772),
.B(n_2718),
.Y(n_3454)
);

AO21x1_ASAP7_75t_L g3455 ( 
.A1(n_2828),
.A2(n_2646),
.B(n_2853),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_2646),
.B(n_2931),
.Y(n_3456)
);

CKINVDCx5p33_ASAP7_75t_R g3457 ( 
.A(n_2691),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_2655),
.B(n_2931),
.Y(n_3458)
);

AOI21x1_ASAP7_75t_L g3459 ( 
.A1(n_2655),
.A2(n_2931),
.B(n_2772),
.Y(n_3459)
);

AOI21x1_ASAP7_75t_SL g3460 ( 
.A1(n_2649),
.A2(n_2432),
.B(n_2708),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_2466),
.A2(n_2624),
.B(n_2595),
.Y(n_3461)
);

A2O1A1Ixp33_ASAP7_75t_L g3462 ( 
.A1(n_2466),
.A2(n_2624),
.B(n_2595),
.C(n_2501),
.Y(n_3462)
);

OAI21xp5_ASAP7_75t_L g3463 ( 
.A1(n_2466),
.A2(n_3028),
.B(n_2528),
.Y(n_3463)
);

HB1xp67_ASAP7_75t_L g3464 ( 
.A(n_2718),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_2501),
.A2(n_3028),
.B(n_2528),
.Y(n_3465)
);

OAI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2501),
.A2(n_3028),
.B(n_2528),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_2718),
.B(n_2931),
.Y(n_3467)
);

A2O1A1Ixp33_ASAP7_75t_L g3468 ( 
.A1(n_2513),
.A2(n_3028),
.B(n_2772),
.C(n_2966),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_2718),
.B(n_2966),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2513),
.A2(n_2853),
.B(n_2772),
.Y(n_3470)
);

A2O1A1Ixp33_ASAP7_75t_L g3471 ( 
.A1(n_2513),
.A2(n_2966),
.B(n_2853),
.C(n_2996),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_2853),
.B(n_2966),
.Y(n_3472)
);

OAI21x1_ASAP7_75t_L g3473 ( 
.A1(n_2853),
.A2(n_2708),
.B(n_2691),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_2649),
.B(n_2396),
.Y(n_3474)
);

OR2x2_ASAP7_75t_L g3475 ( 
.A(n_2534),
.B(n_2588),
.Y(n_3475)
);

AND2x4_ASAP7_75t_L g3476 ( 
.A(n_2588),
.B(n_2604),
.Y(n_3476)
);

AO31x2_ASAP7_75t_L g3477 ( 
.A1(n_2430),
.A2(n_2463),
.A3(n_2817),
.B(n_2387),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3031),
.B(n_2430),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_2996),
.B(n_2409),
.Y(n_3479)
);

A2O1A1Ixp33_ASAP7_75t_L g3480 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3481)
);

NOR2xp33_ASAP7_75t_L g3482 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_2344),
.B(n_2403),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3486)
);

OAI21x1_ASAP7_75t_L g3487 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3488)
);

OAI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3490)
);

OAI21x1_ASAP7_75t_L g3491 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3491)
);

OAI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3492)
);

NOR2xp33_ASAP7_75t_L g3493 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3493)
);

AOI21x1_ASAP7_75t_L g3494 ( 
.A1(n_2981),
.A2(n_1661),
.B(n_1763),
.Y(n_3494)
);

A2O1A1Ixp33_ASAP7_75t_L g3495 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3033),
.B(n_1572),
.Y(n_3496)
);

AOI21xp33_ASAP7_75t_L g3497 ( 
.A1(n_3007),
.A2(n_792),
.B(n_2142),
.Y(n_3497)
);

OAI21x1_ASAP7_75t_L g3498 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3499)
);

BUFx2_ASAP7_75t_L g3500 ( 
.A(n_2647),
.Y(n_3500)
);

AO21x1_ASAP7_75t_L g3501 ( 
.A1(n_2968),
.A2(n_792),
.B(n_3011),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3502)
);

OAI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3033),
.A2(n_1457),
.B1(n_1458),
.B2(n_1433),
.Y(n_3503)
);

NAND2x1p5_ASAP7_75t_L g3504 ( 
.A(n_2451),
.B(n_2386),
.Y(n_3504)
);

OAI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3033),
.A2(n_1457),
.B1(n_1458),
.B2(n_1433),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3507)
);

OAI21x1_ASAP7_75t_L g3508 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3509)
);

OAI21x1_ASAP7_75t_SL g3510 ( 
.A1(n_2491),
.A2(n_2365),
.B(n_2395),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3512)
);

A2O1A1Ixp33_ASAP7_75t_L g3513 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3513)
);

A2O1A1Ixp33_ASAP7_75t_L g3514 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3514)
);

AO31x2_ASAP7_75t_L g3515 ( 
.A1(n_2463),
.A2(n_2817),
.A3(n_2387),
.B(n_2574),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_3033),
.B(n_1572),
.Y(n_3516)
);

INVx2_ASAP7_75t_SL g3517 ( 
.A(n_2415),
.Y(n_3517)
);

BUFx8_ASAP7_75t_L g3518 ( 
.A(n_2541),
.Y(n_3518)
);

INVx3_ASAP7_75t_L g3519 ( 
.A(n_2726),
.Y(n_3519)
);

AOI21xp5_ASAP7_75t_L g3520 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3523)
);

A2O1A1Ixp33_ASAP7_75t_L g3524 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3524)
);

OAI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3525)
);

HB1xp67_ASAP7_75t_L g3526 ( 
.A(n_2364),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3527)
);

OR2x2_ASAP7_75t_L g3528 ( 
.A(n_2361),
.B(n_3012),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_2707),
.Y(n_3529)
);

INVx2_ASAP7_75t_SL g3530 ( 
.A(n_2415),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3531)
);

AND3x4_ASAP7_75t_L g3532 ( 
.A(n_3009),
.B(n_2171),
.C(n_2136),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3534)
);

A2O1A1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3535)
);

AOI21x1_ASAP7_75t_L g3536 ( 
.A1(n_2981),
.A2(n_1661),
.B(n_1763),
.Y(n_3536)
);

NAND2x1p5_ASAP7_75t_L g3537 ( 
.A(n_2451),
.B(n_2386),
.Y(n_3537)
);

HB1xp67_ASAP7_75t_L g3538 ( 
.A(n_2364),
.Y(n_3538)
);

OAI21x1_ASAP7_75t_L g3539 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3540)
);

OAI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3033),
.A2(n_1457),
.B1(n_1458),
.B2(n_1433),
.Y(n_3541)
);

BUFx3_ASAP7_75t_L g3542 ( 
.A(n_2942),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_2707),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3544)
);

O2A1O1Ixp5_ASAP7_75t_L g3545 ( 
.A1(n_3006),
.A2(n_792),
.B(n_1457),
.C(n_1433),
.Y(n_3545)
);

INVx3_ASAP7_75t_L g3546 ( 
.A(n_2726),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3033),
.B(n_1572),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3549)
);

NOR2xp33_ASAP7_75t_L g3550 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3551)
);

A2O1A1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3554)
);

INVx4_ASAP7_75t_L g3555 ( 
.A(n_2567),
.Y(n_3555)
);

OAI21x1_ASAP7_75t_L g3556 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3033),
.B(n_1572),
.Y(n_3557)
);

OAI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3558)
);

OAI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3559)
);

AOI21xp33_ASAP7_75t_L g3560 ( 
.A1(n_3007),
.A2(n_792),
.B(n_2142),
.Y(n_3560)
);

A2O1A1Ixp33_ASAP7_75t_L g3561 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_2364),
.Y(n_3563)
);

INVx6_ASAP7_75t_L g3564 ( 
.A(n_2652),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_SL g3565 ( 
.A1(n_2584),
.A2(n_1146),
.B(n_2946),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2707),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3568)
);

OR2x2_ASAP7_75t_L g3569 ( 
.A(n_2361),
.B(n_3012),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_2707),
.Y(n_3570)
);

CKINVDCx20_ASAP7_75t_R g3571 ( 
.A(n_2507),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3572)
);

A2O1A1Ixp33_ASAP7_75t_L g3573 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3573)
);

OAI21xp33_ASAP7_75t_SL g3574 ( 
.A1(n_2446),
.A2(n_773),
.B(n_1669),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3577)
);

OAI21x1_ASAP7_75t_L g3578 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3579)
);

NOR4xp25_ASAP7_75t_L g3580 ( 
.A(n_3007),
.B(n_1505),
.C(n_1557),
.D(n_1525),
.Y(n_3580)
);

AOI221xp5_ASAP7_75t_L g3581 ( 
.A1(n_3009),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.C(n_1433),
.Y(n_3581)
);

BUFx12f_ASAP7_75t_L g3582 ( 
.A(n_2432),
.Y(n_3582)
);

AOI222xp33_ASAP7_75t_L g3583 ( 
.A1(n_2429),
.A2(n_2368),
.B1(n_2209),
.B2(n_2422),
.C1(n_1458),
.C2(n_1457),
.Y(n_3583)
);

BUFx3_ASAP7_75t_L g3584 ( 
.A(n_2942),
.Y(n_3584)
);

BUFx8_ASAP7_75t_SL g3585 ( 
.A(n_3024),
.Y(n_3585)
);

AOI21x1_ASAP7_75t_SL g3586 ( 
.A1(n_2969),
.A2(n_1445),
.B(n_1443),
.Y(n_3586)
);

OAI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3587)
);

CKINVDCx5p33_ASAP7_75t_R g3588 ( 
.A(n_2653),
.Y(n_3588)
);

A2O1A1Ixp33_ASAP7_75t_L g3589 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3589)
);

AO31x2_ASAP7_75t_L g3590 ( 
.A1(n_2463),
.A2(n_2817),
.A3(n_2387),
.B(n_2574),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3591)
);

AOI211x1_ASAP7_75t_L g3592 ( 
.A1(n_2368),
.A2(n_3006),
.B(n_1525),
.C(n_1557),
.Y(n_3592)
);

BUFx12f_ASAP7_75t_L g3593 ( 
.A(n_2432),
.Y(n_3593)
);

INVx4_ASAP7_75t_L g3594 ( 
.A(n_2567),
.Y(n_3594)
);

BUFx4_ASAP7_75t_SL g3595 ( 
.A(n_2773),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3596)
);

INVx5_ASAP7_75t_L g3597 ( 
.A(n_3035),
.Y(n_3597)
);

NAND2x1p5_ASAP7_75t_L g3598 ( 
.A(n_2451),
.B(n_2386),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_2915),
.Y(n_3599)
);

AOI21x1_ASAP7_75t_L g3600 ( 
.A1(n_2981),
.A2(n_1661),
.B(n_1763),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3603)
);

NAND2xp33_ASAP7_75t_L g3604 ( 
.A(n_3009),
.B(n_366),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3606)
);

AND2x4_ASAP7_75t_L g3607 ( 
.A(n_2344),
.B(n_2403),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_2707),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_SL g3609 ( 
.A1(n_2584),
.A2(n_1146),
.B(n_2946),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3611)
);

HB1xp67_ASAP7_75t_L g3612 ( 
.A(n_2364),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_2707),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3615)
);

INVx4_ASAP7_75t_L g3616 ( 
.A(n_2567),
.Y(n_3616)
);

CKINVDCx5p33_ASAP7_75t_R g3617 ( 
.A(n_2653),
.Y(n_3617)
);

INVxp67_ASAP7_75t_L g3618 ( 
.A(n_2617),
.Y(n_3618)
);

INVx3_ASAP7_75t_SL g3619 ( 
.A(n_2795),
.Y(n_3619)
);

HB1xp67_ASAP7_75t_L g3620 ( 
.A(n_2364),
.Y(n_3620)
);

AOI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3007),
.A2(n_792),
.B(n_2142),
.Y(n_3621)
);

AND2x2_ASAP7_75t_SL g3622 ( 
.A(n_2435),
.B(n_2392),
.Y(n_3622)
);

OAI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_3033),
.A2(n_1457),
.B1(n_1458),
.B2(n_1433),
.Y(n_3623)
);

AOI22xp5_ASAP7_75t_L g3624 ( 
.A1(n_2368),
.A2(n_1433),
.B1(n_1458),
.B2(n_1457),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_SL g3625 ( 
.A1(n_2491),
.A2(n_2365),
.B(n_2395),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3626)
);

INVxp67_ASAP7_75t_SL g3627 ( 
.A(n_2345),
.Y(n_3627)
);

OAI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3628)
);

BUFx12f_ASAP7_75t_L g3629 ( 
.A(n_2432),
.Y(n_3629)
);

INVx5_ASAP7_75t_L g3630 ( 
.A(n_3035),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_2707),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_L g3632 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_2707),
.Y(n_3633)
);

OR2x2_ASAP7_75t_L g3634 ( 
.A(n_2361),
.B(n_3012),
.Y(n_3634)
);

INVxp67_ASAP7_75t_L g3635 ( 
.A(n_2617),
.Y(n_3635)
);

INVx4_ASAP7_75t_L g3636 ( 
.A(n_2567),
.Y(n_3636)
);

A2O1A1Ixp33_ASAP7_75t_L g3637 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3637)
);

AOI221xp5_ASAP7_75t_L g3638 ( 
.A1(n_3009),
.A2(n_1458),
.B1(n_1478),
.B2(n_1457),
.C(n_1433),
.Y(n_3638)
);

OAI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3639)
);

A2O1A1Ixp33_ASAP7_75t_L g3640 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3642)
);

AOI221x1_ASAP7_75t_L g3643 ( 
.A1(n_3009),
.A2(n_3013),
.B1(n_2171),
.B2(n_2104),
.C(n_2392),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3645)
);

BUFx2_ASAP7_75t_L g3646 ( 
.A(n_2647),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_L g3647 ( 
.A(n_2368),
.B(n_2349),
.Y(n_3647)
);

OAI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3648)
);

OAI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3007),
.A2(n_1476),
.B(n_792),
.Y(n_3649)
);

AND2x4_ASAP7_75t_L g3650 ( 
.A(n_2344),
.B(n_2403),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3651)
);

AO31x2_ASAP7_75t_L g3652 ( 
.A1(n_2463),
.A2(n_2817),
.A3(n_2387),
.B(n_2574),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3653)
);

INVx4_ASAP7_75t_L g3654 ( 
.A(n_2567),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3655)
);

AOI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_2972),
.A2(n_2983),
.B(n_2980),
.Y(n_3656)
);

OAI21x1_ASAP7_75t_L g3657 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3657)
);

NOR2xp67_ASAP7_75t_SL g3658 ( 
.A(n_2691),
.B(n_1505),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_2915),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_2915),
.Y(n_3660)
);

O2A1O1Ixp5_ASAP7_75t_L g3661 ( 
.A1(n_3006),
.A2(n_792),
.B(n_1457),
.C(n_1433),
.Y(n_3661)
);

AOI221x1_ASAP7_75t_L g3662 ( 
.A1(n_3009),
.A2(n_3013),
.B1(n_2171),
.B2(n_2104),
.C(n_2392),
.Y(n_3662)
);

BUFx6f_ASAP7_75t_L g3663 ( 
.A(n_2726),
.Y(n_3663)
);

AND2x2_ASAP7_75t_L g3664 ( 
.A(n_2409),
.B(n_2427),
.Y(n_3664)
);

A2O1A1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_2368),
.A2(n_1433),
.B(n_1458),
.C(n_1457),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_2915),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_2707),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_2982),
.A2(n_1800),
.B(n_2362),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_2485),
.B(n_2370),
.Y(n_3669)
);

INVx1_ASAP7_75t_SL g3670 ( 
.A(n_3045),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3230),
.B(n_3244),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3179),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3663),
.Y(n_3673)
);

BUFx2_ASAP7_75t_L g3674 ( 
.A(n_3244),
.Y(n_3674)
);

CKINVDCx16_ASAP7_75t_R g3675 ( 
.A(n_3041),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3230),
.B(n_3244),
.Y(n_3676)
);

INVx4_ASAP7_75t_L g3677 ( 
.A(n_3134),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3179),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3052),
.B(n_3597),
.Y(n_3679)
);

INVx4_ASAP7_75t_L g3680 ( 
.A(n_3134),
.Y(n_3680)
);

INVx5_ASAP7_75t_L g3681 ( 
.A(n_3058),
.Y(n_3681)
);

BUFx12f_ASAP7_75t_L g3682 ( 
.A(n_3250),
.Y(n_3682)
);

INVx2_ASAP7_75t_SL g3683 ( 
.A(n_3047),
.Y(n_3683)
);

INVx2_ASAP7_75t_SL g3684 ( 
.A(n_3047),
.Y(n_3684)
);

HB1xp67_ASAP7_75t_L g3685 ( 
.A(n_3432),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3186),
.Y(n_3686)
);

BUFx4f_ASAP7_75t_L g3687 ( 
.A(n_3366),
.Y(n_3687)
);

HB1xp67_ASAP7_75t_L g3688 ( 
.A(n_3432),
.Y(n_3688)
);

NAND2x1p5_ASAP7_75t_L g3689 ( 
.A(n_3052),
.B(n_3597),
.Y(n_3689)
);

BUFx3_ASAP7_75t_L g3690 ( 
.A(n_3065),
.Y(n_3690)
);

HB1xp67_ASAP7_75t_L g3691 ( 
.A(n_3162),
.Y(n_3691)
);

INVxp67_ASAP7_75t_SL g3692 ( 
.A(n_3050),
.Y(n_3692)
);

BUFx3_ASAP7_75t_L g3693 ( 
.A(n_3065),
.Y(n_3693)
);

BUFx8_ASAP7_75t_L g3694 ( 
.A(n_3041),
.Y(n_3694)
);

INVx3_ASAP7_75t_L g3695 ( 
.A(n_3047),
.Y(n_3695)
);

INVx5_ASAP7_75t_L g3696 ( 
.A(n_3058),
.Y(n_3696)
);

INVx6_ASAP7_75t_SL g3697 ( 
.A(n_3244),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3186),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_3585),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3247),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_L g3701 ( 
.A(n_3141),
.B(n_3084),
.Y(n_3701)
);

BUFx3_ASAP7_75t_L g3702 ( 
.A(n_3065),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3247),
.Y(n_3703)
);

INVx1_ASAP7_75t_SL g3704 ( 
.A(n_3045),
.Y(n_3704)
);

OR2x2_ASAP7_75t_L g3705 ( 
.A(n_3201),
.B(n_3162),
.Y(n_3705)
);

INVx1_ASAP7_75t_SL g3706 ( 
.A(n_3278),
.Y(n_3706)
);

BUFx2_ASAP7_75t_R g3707 ( 
.A(n_3457),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3251),
.Y(n_3708)
);

INVx3_ASAP7_75t_L g3709 ( 
.A(n_3074),
.Y(n_3709)
);

INVx3_ASAP7_75t_L g3710 ( 
.A(n_3074),
.Y(n_3710)
);

INVx6_ASAP7_75t_L g3711 ( 
.A(n_3065),
.Y(n_3711)
);

BUFx2_ASAP7_75t_R g3712 ( 
.A(n_3619),
.Y(n_3712)
);

INVx5_ASAP7_75t_SL g3713 ( 
.A(n_3058),
.Y(n_3713)
);

INVx1_ASAP7_75t_SL g3714 ( 
.A(n_3278),
.Y(n_3714)
);

BUFx12f_ASAP7_75t_L g3715 ( 
.A(n_3365),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3251),
.Y(n_3716)
);

BUFx3_ASAP7_75t_L g3717 ( 
.A(n_3151),
.Y(n_3717)
);

BUFx4f_ASAP7_75t_SL g3718 ( 
.A(n_3041),
.Y(n_3718)
);

BUFx3_ASAP7_75t_L g3719 ( 
.A(n_3151),
.Y(n_3719)
);

AND2x6_ASAP7_75t_L g3720 ( 
.A(n_3204),
.B(n_3271),
.Y(n_3720)
);

BUFx12f_ASAP7_75t_L g3721 ( 
.A(n_3168),
.Y(n_3721)
);

BUFx3_ASAP7_75t_L g3722 ( 
.A(n_3151),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3147),
.B(n_3153),
.Y(n_3723)
);

BUFx12f_ASAP7_75t_L g3724 ( 
.A(n_3169),
.Y(n_3724)
);

BUFx2_ASAP7_75t_SL g3725 ( 
.A(n_3455),
.Y(n_3725)
);

BUFx2_ASAP7_75t_L g3726 ( 
.A(n_3253),
.Y(n_3726)
);

CKINVDCx20_ASAP7_75t_R g3727 ( 
.A(n_3341),
.Y(n_3727)
);

BUFx2_ASAP7_75t_L g3728 ( 
.A(n_3253),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3147),
.B(n_3153),
.Y(n_3729)
);

INVx6_ASAP7_75t_L g3730 ( 
.A(n_3151),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3279),
.Y(n_3731)
);

BUFx12f_ASAP7_75t_L g3732 ( 
.A(n_3588),
.Y(n_3732)
);

INVx3_ASAP7_75t_SL g3733 ( 
.A(n_3622),
.Y(n_3733)
);

NAND2x1p5_ASAP7_75t_L g3734 ( 
.A(n_3052),
.B(n_3597),
.Y(n_3734)
);

BUFx2_ASAP7_75t_SL g3735 ( 
.A(n_3455),
.Y(n_3735)
);

BUFx3_ASAP7_75t_L g3736 ( 
.A(n_3518),
.Y(n_3736)
);

BUFx2_ASAP7_75t_R g3737 ( 
.A(n_3619),
.Y(n_3737)
);

BUFx6f_ASAP7_75t_SL g3738 ( 
.A(n_3326),
.Y(n_3738)
);

INVx5_ASAP7_75t_L g3739 ( 
.A(n_3058),
.Y(n_3739)
);

INVx4_ASAP7_75t_L g3740 ( 
.A(n_3134),
.Y(n_3740)
);

NAND2x1p5_ASAP7_75t_L g3741 ( 
.A(n_3052),
.B(n_3597),
.Y(n_3741)
);

BUFx3_ASAP7_75t_L g3742 ( 
.A(n_3518),
.Y(n_3742)
);

INVx3_ASAP7_75t_SL g3743 ( 
.A(n_3622),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3279),
.Y(n_3744)
);

AOI22xp33_ASAP7_75t_L g3745 ( 
.A1(n_3532),
.A2(n_3638),
.B1(n_3581),
.B2(n_3583),
.Y(n_3745)
);

BUFx3_ASAP7_75t_L g3746 ( 
.A(n_3518),
.Y(n_3746)
);

CKINVDCx5p33_ASAP7_75t_R g3747 ( 
.A(n_3059),
.Y(n_3747)
);

BUFx3_ASAP7_75t_L g3748 ( 
.A(n_3518),
.Y(n_3748)
);

INVx3_ASAP7_75t_L g3749 ( 
.A(n_3074),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3282),
.Y(n_3750)
);

INVxp67_ASAP7_75t_SL g3751 ( 
.A(n_3050),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3099),
.B(n_3125),
.Y(n_3752)
);

INVx4_ASAP7_75t_L g3753 ( 
.A(n_3134),
.Y(n_3753)
);

INVx6_ASAP7_75t_L g3754 ( 
.A(n_3326),
.Y(n_3754)
);

BUFx3_ASAP7_75t_L g3755 ( 
.A(n_3326),
.Y(n_3755)
);

INVx4_ASAP7_75t_L g3756 ( 
.A(n_3049),
.Y(n_3756)
);

CKINVDCx20_ASAP7_75t_R g3757 ( 
.A(n_3571),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3099),
.B(n_3113),
.Y(n_3758)
);

CKINVDCx20_ASAP7_75t_R g3759 ( 
.A(n_3617),
.Y(n_3759)
);

BUFx3_ASAP7_75t_L g3760 ( 
.A(n_3326),
.Y(n_3760)
);

BUFx8_ASAP7_75t_SL g3761 ( 
.A(n_3311),
.Y(n_3761)
);

CKINVDCx5p33_ASAP7_75t_R g3762 ( 
.A(n_3184),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3292),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3113),
.B(n_3120),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3323),
.Y(n_3765)
);

BUFx2_ASAP7_75t_SL g3766 ( 
.A(n_3434),
.Y(n_3766)
);

INVx5_ASAP7_75t_L g3767 ( 
.A(n_3058),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3323),
.Y(n_3768)
);

INVx3_ASAP7_75t_SL g3769 ( 
.A(n_3622),
.Y(n_3769)
);

INVx4_ASAP7_75t_L g3770 ( 
.A(n_3049),
.Y(n_3770)
);

BUFx12f_ASAP7_75t_L g3771 ( 
.A(n_3311),
.Y(n_3771)
);

INVx1_ASAP7_75t_SL g3772 ( 
.A(n_3348),
.Y(n_3772)
);

NAND2x1p5_ASAP7_75t_L g3773 ( 
.A(n_3052),
.B(n_3597),
.Y(n_3773)
);

BUFx12f_ASAP7_75t_L g3774 ( 
.A(n_3311),
.Y(n_3774)
);

BUFx3_ASAP7_75t_L g3775 ( 
.A(n_3454),
.Y(n_3775)
);

INVx3_ASAP7_75t_SL g3776 ( 
.A(n_3476),
.Y(n_3776)
);

CKINVDCx20_ASAP7_75t_R g3777 ( 
.A(n_3619),
.Y(n_3777)
);

NOR2xp33_ASAP7_75t_L g3778 ( 
.A(n_3532),
.B(n_3183),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3038),
.Y(n_3779)
);

BUFx2_ASAP7_75t_SL g3780 ( 
.A(n_3434),
.Y(n_3780)
);

BUFx2_ASAP7_75t_L g3781 ( 
.A(n_3253),
.Y(n_3781)
);

CKINVDCx20_ASAP7_75t_R g3782 ( 
.A(n_3404),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3181),
.B(n_3160),
.Y(n_3783)
);

INVx3_ASAP7_75t_L g3784 ( 
.A(n_3074),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3230),
.B(n_3253),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3230),
.B(n_3201),
.Y(n_3786)
);

INVx4_ASAP7_75t_L g3787 ( 
.A(n_3049),
.Y(n_3787)
);

INVx6_ASAP7_75t_L g3788 ( 
.A(n_3304),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3599),
.Y(n_3789)
);

INVx3_ASAP7_75t_SL g3790 ( 
.A(n_3476),
.Y(n_3790)
);

NAND2x1p5_ASAP7_75t_L g3791 ( 
.A(n_3052),
.B(n_3597),
.Y(n_3791)
);

BUFx12f_ASAP7_75t_L g3792 ( 
.A(n_3582),
.Y(n_3792)
);

INVx3_ASAP7_75t_SL g3793 ( 
.A(n_3476),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3038),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3039),
.Y(n_3795)
);

INVx1_ASAP7_75t_SL g3796 ( 
.A(n_3348),
.Y(n_3796)
);

BUFx2_ASAP7_75t_SL g3797 ( 
.A(n_3290),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3659),
.Y(n_3798)
);

BUFx12f_ASAP7_75t_L g3799 ( 
.A(n_3582),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3532),
.B(n_3183),
.Y(n_3800)
);

INVx5_ASAP7_75t_SL g3801 ( 
.A(n_3301),
.Y(n_3801)
);

INVx8_ASAP7_75t_L g3802 ( 
.A(n_3366),
.Y(n_3802)
);

NAND2x1p5_ASAP7_75t_L g3803 ( 
.A(n_3630),
.B(n_3049),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3659),
.Y(n_3804)
);

INVx2_ASAP7_75t_SL g3805 ( 
.A(n_3095),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3659),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3660),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3181),
.B(n_3160),
.Y(n_3808)
);

INVx4_ASAP7_75t_L g3809 ( 
.A(n_3555),
.Y(n_3809)
);

BUFx2_ASAP7_75t_R g3810 ( 
.A(n_3474),
.Y(n_3810)
);

BUFx4f_ASAP7_75t_SL g3811 ( 
.A(n_3582),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3660),
.Y(n_3812)
);

NOR2xp33_ASAP7_75t_SL g3813 ( 
.A(n_3075),
.B(n_3072),
.Y(n_3813)
);

INVx1_ASAP7_75t_SL g3814 ( 
.A(n_3293),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3660),
.Y(n_3815)
);

INVx1_ASAP7_75t_SL g3816 ( 
.A(n_3293),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3039),
.Y(n_3817)
);

BUFx2_ASAP7_75t_L g3818 ( 
.A(n_3201),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3581),
.A2(n_3638),
.B1(n_3583),
.B2(n_3072),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3489),
.B(n_3492),
.Y(n_3820)
);

BUFx3_ASAP7_75t_L g3821 ( 
.A(n_3454),
.Y(n_3821)
);

INVx4_ASAP7_75t_L g3822 ( 
.A(n_3555),
.Y(n_3822)
);

BUFx3_ASAP7_75t_L g3823 ( 
.A(n_3454),
.Y(n_3823)
);

INVxp67_ASAP7_75t_SL g3824 ( 
.A(n_3486),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3666),
.Y(n_3825)
);

CKINVDCx5p33_ASAP7_75t_R g3826 ( 
.A(n_3595),
.Y(n_3826)
);

INVx2_ASAP7_75t_SL g3827 ( 
.A(n_3106),
.Y(n_3827)
);

CKINVDCx6p67_ASAP7_75t_R g3828 ( 
.A(n_3593),
.Y(n_3828)
);

AND2x4_ASAP7_75t_L g3829 ( 
.A(n_3630),
.B(n_3055),
.Y(n_3829)
);

INVx4_ASAP7_75t_L g3830 ( 
.A(n_3555),
.Y(n_3830)
);

CKINVDCx16_ASAP7_75t_R g3831 ( 
.A(n_3593),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3161),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3053),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3230),
.B(n_3201),
.Y(n_3834)
);

BUFx12f_ASAP7_75t_L g3835 ( 
.A(n_3593),
.Y(n_3835)
);

BUFx3_ASAP7_75t_L g3836 ( 
.A(n_3454),
.Y(n_3836)
);

AND2x4_ASAP7_75t_L g3837 ( 
.A(n_3630),
.B(n_3055),
.Y(n_3837)
);

CKINVDCx16_ASAP7_75t_R g3838 ( 
.A(n_3629),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3053),
.Y(n_3839)
);

INVxp67_ASAP7_75t_SL g3840 ( 
.A(n_3486),
.Y(n_3840)
);

OR2x2_ASAP7_75t_L g3841 ( 
.A(n_3201),
.B(n_3139),
.Y(n_3841)
);

INVx2_ASAP7_75t_SL g3842 ( 
.A(n_3106),
.Y(n_3842)
);

INVx1_ASAP7_75t_SL g3843 ( 
.A(n_3423),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3102),
.B(n_3107),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3062),
.Y(n_3845)
);

BUFx3_ASAP7_75t_L g3846 ( 
.A(n_3473),
.Y(n_3846)
);

CKINVDCx16_ASAP7_75t_R g3847 ( 
.A(n_3629),
.Y(n_3847)
);

BUFx3_ASAP7_75t_L g3848 ( 
.A(n_3473),
.Y(n_3848)
);

BUFx3_ASAP7_75t_L g3849 ( 
.A(n_3367),
.Y(n_3849)
);

BUFx3_ASAP7_75t_L g3850 ( 
.A(n_3367),
.Y(n_3850)
);

INVx3_ASAP7_75t_L g3851 ( 
.A(n_3106),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3062),
.Y(n_3852)
);

INVx1_ASAP7_75t_SL g3853 ( 
.A(n_3423),
.Y(n_3853)
);

BUFx4f_ASAP7_75t_SL g3854 ( 
.A(n_3629),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3103),
.Y(n_3855)
);

BUFx2_ASAP7_75t_SL g3856 ( 
.A(n_3290),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3103),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3161),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3161),
.Y(n_3859)
);

INVx1_ASAP7_75t_SL g3860 ( 
.A(n_3418),
.Y(n_3860)
);

BUFx3_ASAP7_75t_L g3861 ( 
.A(n_3367),
.Y(n_3861)
);

INVx2_ASAP7_75t_SL g3862 ( 
.A(n_3106),
.Y(n_3862)
);

BUFx3_ASAP7_75t_L g3863 ( 
.A(n_3373),
.Y(n_3863)
);

BUFx8_ASAP7_75t_L g3864 ( 
.A(n_3366),
.Y(n_3864)
);

BUFx4_ASAP7_75t_SL g3865 ( 
.A(n_3453),
.Y(n_3865)
);

BUFx3_ASAP7_75t_L g3866 ( 
.A(n_3373),
.Y(n_3866)
);

BUFx4_ASAP7_75t_SL g3867 ( 
.A(n_3453),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3132),
.Y(n_3868)
);

NAND2x1p5_ASAP7_75t_L g3869 ( 
.A(n_3630),
.B(n_3555),
.Y(n_3869)
);

BUFx3_ASAP7_75t_L g3870 ( 
.A(n_3373),
.Y(n_3870)
);

BUFx2_ASAP7_75t_SL g3871 ( 
.A(n_3077),
.Y(n_3871)
);

CKINVDCx5p33_ASAP7_75t_R g3872 ( 
.A(n_3404),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3135),
.B(n_3425),
.Y(n_3873)
);

CKINVDCx11_ASAP7_75t_R g3874 ( 
.A(n_3476),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_L g3875 ( 
.A1(n_3128),
.A2(n_3503),
.B1(n_3541),
.B2(n_3505),
.Y(n_3875)
);

BUFx2_ASAP7_75t_L g3876 ( 
.A(n_3411),
.Y(n_3876)
);

NAND2x1p5_ASAP7_75t_L g3877 ( 
.A(n_3630),
.B(n_3594),
.Y(n_3877)
);

BUFx8_ASAP7_75t_L g3878 ( 
.A(n_3366),
.Y(n_3878)
);

INVx5_ASAP7_75t_SL g3879 ( 
.A(n_3301),
.Y(n_3879)
);

BUFx2_ASAP7_75t_SL g3880 ( 
.A(n_3077),
.Y(n_3880)
);

INVx2_ASAP7_75t_SL g3881 ( 
.A(n_3630),
.Y(n_3881)
);

BUFx12f_ASAP7_75t_L g3882 ( 
.A(n_3475),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3061),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3132),
.Y(n_3884)
);

INVx2_ASAP7_75t_SL g3885 ( 
.A(n_3257),
.Y(n_3885)
);

OR2x6_ASAP7_75t_L g3886 ( 
.A(n_3073),
.B(n_3178),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3529),
.Y(n_3887)
);

INVx6_ASAP7_75t_L g3888 ( 
.A(n_3435),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3529),
.Y(n_3889)
);

BUFx12f_ASAP7_75t_L g3890 ( 
.A(n_3475),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3061),
.Y(n_3891)
);

BUFx3_ASAP7_75t_L g3892 ( 
.A(n_3438),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3543),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3543),
.Y(n_3894)
);

INVx1_ASAP7_75t_SL g3895 ( 
.A(n_3526),
.Y(n_3895)
);

INVx6_ASAP7_75t_SL g3896 ( 
.A(n_3178),
.Y(n_3896)
);

CKINVDCx16_ASAP7_75t_R g3897 ( 
.A(n_3214),
.Y(n_3897)
);

BUFx3_ASAP7_75t_L g3898 ( 
.A(n_3257),
.Y(n_3898)
);

BUFx2_ASAP7_75t_SL g3899 ( 
.A(n_3077),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3102),
.B(n_3107),
.Y(n_3900)
);

INVx8_ASAP7_75t_L g3901 ( 
.A(n_3366),
.Y(n_3901)
);

BUFx3_ASAP7_75t_L g3902 ( 
.A(n_3435),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3086),
.Y(n_3903)
);

AOI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3503),
.A2(n_3505),
.B1(n_3623),
.B2(n_3541),
.Y(n_3904)
);

NAND2x1p5_ASAP7_75t_L g3905 ( 
.A(n_3594),
.B(n_3616),
.Y(n_3905)
);

CKINVDCx16_ASAP7_75t_R g3906 ( 
.A(n_3198),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3566),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3566),
.Y(n_3908)
);

BUFx3_ASAP7_75t_L g3909 ( 
.A(n_3435),
.Y(n_3909)
);

INVx4_ASAP7_75t_L g3910 ( 
.A(n_3594),
.Y(n_3910)
);

NAND2x1p5_ASAP7_75t_L g3911 ( 
.A(n_3594),
.B(n_3616),
.Y(n_3911)
);

INVx6_ASAP7_75t_L g3912 ( 
.A(n_3435),
.Y(n_3912)
);

BUFx3_ASAP7_75t_L g3913 ( 
.A(n_3068),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_L g3914 ( 
.A1(n_3128),
.A2(n_3623),
.B1(n_3109),
.B2(n_3218),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3570),
.Y(n_3915)
);

INVxp67_ASAP7_75t_SL g3916 ( 
.A(n_3490),
.Y(n_3916)
);

BUFx2_ASAP7_75t_SL g3917 ( 
.A(n_3198),
.Y(n_3917)
);

INVx4_ASAP7_75t_L g3918 ( 
.A(n_3616),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3570),
.Y(n_3919)
);

INVx3_ASAP7_75t_SL g3920 ( 
.A(n_3564),
.Y(n_3920)
);

AND2x4_ASAP7_75t_L g3921 ( 
.A(n_3055),
.B(n_3228),
.Y(n_3921)
);

INVx1_ASAP7_75t_SL g3922 ( 
.A(n_3538),
.Y(n_3922)
);

INVx1_ASAP7_75t_SL g3923 ( 
.A(n_3563),
.Y(n_3923)
);

BUFx3_ASAP7_75t_L g3924 ( 
.A(n_3068),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3608),
.Y(n_3925)
);

AOI22xp5_ASAP7_75t_L g3926 ( 
.A1(n_3218),
.A2(n_3624),
.B1(n_3081),
.B2(n_3199),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3608),
.Y(n_3927)
);

BUFx12f_ASAP7_75t_L g3928 ( 
.A(n_3478),
.Y(n_3928)
);

INVx5_ASAP7_75t_L g3929 ( 
.A(n_3178),
.Y(n_3929)
);

HB1xp67_ASAP7_75t_SL g3930 ( 
.A(n_3198),
.Y(n_3930)
);

INVx4_ASAP7_75t_L g3931 ( 
.A(n_3616),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3081),
.A2(n_3069),
.B1(n_3492),
.B2(n_3489),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3613),
.Y(n_3933)
);

CKINVDCx20_ASAP7_75t_R g3934 ( 
.A(n_3478),
.Y(n_3934)
);

INVx3_ASAP7_75t_L g3935 ( 
.A(n_3064),
.Y(n_3935)
);

BUFx12f_ASAP7_75t_L g3936 ( 
.A(n_3379),
.Y(n_3936)
);

BUFx10_ASAP7_75t_L g3937 ( 
.A(n_3213),
.Y(n_3937)
);

INVx3_ASAP7_75t_SL g3938 ( 
.A(n_3564),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3156),
.B(n_3219),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3613),
.Y(n_3940)
);

INVx3_ASAP7_75t_L g3941 ( 
.A(n_3070),
.Y(n_3941)
);

CKINVDCx6p67_ASAP7_75t_R g3942 ( 
.A(n_3474),
.Y(n_3942)
);

INVx1_ASAP7_75t_SL g3943 ( 
.A(n_3612),
.Y(n_3943)
);

CKINVDCx20_ASAP7_75t_R g3944 ( 
.A(n_3116),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3631),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3156),
.B(n_3082),
.Y(n_3946)
);

INVx4_ASAP7_75t_L g3947 ( 
.A(n_3636),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3082),
.B(n_3088),
.Y(n_3948)
);

INVx3_ASAP7_75t_L g3949 ( 
.A(n_3070),
.Y(n_3949)
);

INVxp67_ASAP7_75t_SL g3950 ( 
.A(n_3490),
.Y(n_3950)
);

INVx1_ASAP7_75t_SL g3951 ( 
.A(n_3620),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3631),
.Y(n_3952)
);

BUFx3_ASAP7_75t_L g3953 ( 
.A(n_3068),
.Y(n_3953)
);

CKINVDCx6p67_ASAP7_75t_R g3954 ( 
.A(n_3542),
.Y(n_3954)
);

INVx1_ASAP7_75t_SL g3955 ( 
.A(n_3288),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3088),
.B(n_3159),
.Y(n_3956)
);

BUFx2_ASAP7_75t_L g3957 ( 
.A(n_3411),
.Y(n_3957)
);

BUFx12f_ASAP7_75t_L g3958 ( 
.A(n_3379),
.Y(n_3958)
);

INVxp67_ASAP7_75t_SL g3959 ( 
.A(n_3502),
.Y(n_3959)
);

BUFx2_ASAP7_75t_SL g3960 ( 
.A(n_3542),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_3315),
.Y(n_3961)
);

BUFx3_ASAP7_75t_L g3962 ( 
.A(n_3504),
.Y(n_3962)
);

BUFx2_ASAP7_75t_SL g3963 ( 
.A(n_3542),
.Y(n_3963)
);

BUFx4f_ASAP7_75t_L g3964 ( 
.A(n_3241),
.Y(n_3964)
);

BUFx12f_ASAP7_75t_L g3965 ( 
.A(n_3379),
.Y(n_3965)
);

INVx3_ASAP7_75t_SL g3966 ( 
.A(n_3564),
.Y(n_3966)
);

AO22x2_ASAP7_75t_L g3967 ( 
.A1(n_3044),
.A2(n_3199),
.B1(n_3202),
.B2(n_3643),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3633),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3633),
.Y(n_3969)
);

NAND2x1p5_ASAP7_75t_L g3970 ( 
.A(n_3636),
.B(n_3654),
.Y(n_3970)
);

BUFx2_ASAP7_75t_SL g3971 ( 
.A(n_3584),
.Y(n_3971)
);

NOR2xp33_ASAP7_75t_L g3972 ( 
.A(n_3497),
.B(n_3560),
.Y(n_3972)
);

INVx3_ASAP7_75t_L g3973 ( 
.A(n_3070),
.Y(n_3973)
);

BUFx6f_ASAP7_75t_L g3974 ( 
.A(n_3178),
.Y(n_3974)
);

BUFx6f_ASAP7_75t_L g3975 ( 
.A(n_3178),
.Y(n_3975)
);

INVx1_ASAP7_75t_SL g3976 ( 
.A(n_3322),
.Y(n_3976)
);

INVx3_ASAP7_75t_L g3977 ( 
.A(n_3070),
.Y(n_3977)
);

BUFx3_ASAP7_75t_L g3978 ( 
.A(n_3504),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3667),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3667),
.Y(n_3980)
);

INVxp67_ASAP7_75t_SL g3981 ( 
.A(n_3502),
.Y(n_3981)
);

AND2x4_ASAP7_75t_L g3982 ( 
.A(n_3055),
.B(n_3228),
.Y(n_3982)
);

INVx3_ASAP7_75t_L g3983 ( 
.A(n_3036),
.Y(n_3983)
);

BUFx6f_ASAP7_75t_L g3984 ( 
.A(n_3229),
.Y(n_3984)
);

BUFx12f_ASAP7_75t_L g3985 ( 
.A(n_3379),
.Y(n_3985)
);

BUFx6f_ASAP7_75t_L g3986 ( 
.A(n_3229),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3422),
.Y(n_3987)
);

BUFx3_ASAP7_75t_L g3988 ( 
.A(n_3504),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3159),
.B(n_3165),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3422),
.Y(n_3990)
);

BUFx3_ASAP7_75t_L g3991 ( 
.A(n_3537),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3165),
.B(n_3167),
.Y(n_3992)
);

INVx3_ASAP7_75t_L g3993 ( 
.A(n_3036),
.Y(n_3993)
);

NAND2x1p5_ASAP7_75t_L g3994 ( 
.A(n_3636),
.B(n_3654),
.Y(n_3994)
);

BUFx3_ASAP7_75t_L g3995 ( 
.A(n_3537),
.Y(n_3995)
);

INVx6_ASAP7_75t_SL g3996 ( 
.A(n_3228),
.Y(n_3996)
);

INVxp67_ASAP7_75t_SL g3997 ( 
.A(n_3512),
.Y(n_3997)
);

INVx1_ASAP7_75t_SL g3998 ( 
.A(n_3329),
.Y(n_3998)
);

BUFx3_ASAP7_75t_L g3999 ( 
.A(n_3537),
.Y(n_3999)
);

INVx4_ASAP7_75t_L g4000 ( 
.A(n_3636),
.Y(n_4000)
);

BUFx3_ASAP7_75t_L g4001 ( 
.A(n_3598),
.Y(n_4001)
);

INVx4_ASAP7_75t_L g4002 ( 
.A(n_3654),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3356),
.Y(n_4003)
);

CKINVDCx5p33_ASAP7_75t_R g4004 ( 
.A(n_3618),
.Y(n_4004)
);

BUFx12f_ASAP7_75t_L g4005 ( 
.A(n_3400),
.Y(n_4005)
);

INVxp67_ASAP7_75t_SL g4006 ( 
.A(n_3512),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3356),
.Y(n_4007)
);

BUFx12f_ASAP7_75t_L g4008 ( 
.A(n_3400),
.Y(n_4008)
);

CKINVDCx14_ASAP7_75t_R g4009 ( 
.A(n_3479),
.Y(n_4009)
);

INVx3_ASAP7_75t_SL g4010 ( 
.A(n_3564),
.Y(n_4010)
);

BUFx2_ASAP7_75t_L g4011 ( 
.A(n_3192),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3362),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_3635),
.Y(n_4013)
);

INVx3_ASAP7_75t_L g4014 ( 
.A(n_3036),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3362),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3167),
.B(n_3173),
.Y(n_4016)
);

INVx3_ASAP7_75t_L g4017 ( 
.A(n_3036),
.Y(n_4017)
);

INVx1_ASAP7_75t_SL g4018 ( 
.A(n_3425),
.Y(n_4018)
);

OR2x2_ASAP7_75t_L g4019 ( 
.A(n_3139),
.B(n_3142),
.Y(n_4019)
);

NOR2xp33_ASAP7_75t_L g4020 ( 
.A(n_3497),
.B(n_3560),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3135),
.B(n_3228),
.Y(n_4021)
);

INVx1_ASAP7_75t_SL g4022 ( 
.A(n_3444),
.Y(n_4022)
);

AND2x4_ASAP7_75t_L g4023 ( 
.A(n_3483),
.B(n_3607),
.Y(n_4023)
);

BUFx2_ASAP7_75t_SL g4024 ( 
.A(n_3584),
.Y(n_4024)
);

BUFx12f_ASAP7_75t_L g4025 ( 
.A(n_3400),
.Y(n_4025)
);

INVx1_ASAP7_75t_SL g4026 ( 
.A(n_3444),
.Y(n_4026)
);

OR2x2_ASAP7_75t_L g4027 ( 
.A(n_3139),
.B(n_3142),
.Y(n_4027)
);

NAND2x1p5_ASAP7_75t_L g4028 ( 
.A(n_3654),
.B(n_3197),
.Y(n_4028)
);

NAND2x1p5_ASAP7_75t_L g4029 ( 
.A(n_3197),
.B(n_3154),
.Y(n_4029)
);

BUFx2_ASAP7_75t_SL g4030 ( 
.A(n_3584),
.Y(n_4030)
);

INVx1_ASAP7_75t_SL g4031 ( 
.A(n_3447),
.Y(n_4031)
);

INVxp67_ASAP7_75t_SL g4032 ( 
.A(n_3521),
.Y(n_4032)
);

INVx1_ASAP7_75t_SL g4033 ( 
.A(n_3447),
.Y(n_4033)
);

NAND2x1p5_ASAP7_75t_L g4034 ( 
.A(n_3154),
.B(n_3117),
.Y(n_4034)
);

INVx2_ASAP7_75t_SL g4035 ( 
.A(n_3255),
.Y(n_4035)
);

INVx1_ASAP7_75t_SL g4036 ( 
.A(n_3448),
.Y(n_4036)
);

BUFx3_ASAP7_75t_L g4037 ( 
.A(n_3342),
.Y(n_4037)
);

INVx2_ASAP7_75t_SL g4038 ( 
.A(n_3255),
.Y(n_4038)
);

BUFx2_ASAP7_75t_L g4039 ( 
.A(n_3192),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3135),
.B(n_3483),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3135),
.B(n_3483),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3483),
.B(n_3607),
.Y(n_4042)
);

INVx2_ASAP7_75t_SL g4043 ( 
.A(n_3607),
.Y(n_4043)
);

INVx1_ASAP7_75t_SL g4044 ( 
.A(n_3448),
.Y(n_4044)
);

INVx1_ASAP7_75t_SL g4045 ( 
.A(n_3391),
.Y(n_4045)
);

NAND2x1p5_ASAP7_75t_L g4046 ( 
.A(n_3108),
.B(n_3115),
.Y(n_4046)
);

AND2x4_ASAP7_75t_L g4047 ( 
.A(n_3607),
.B(n_3650),
.Y(n_4047)
);

INVx3_ASAP7_75t_L g4048 ( 
.A(n_3519),
.Y(n_4048)
);

INVx4_ASAP7_75t_L g4049 ( 
.A(n_3196),
.Y(n_4049)
);

BUFx4f_ASAP7_75t_L g4050 ( 
.A(n_3241),
.Y(n_4050)
);

OR2x2_ASAP7_75t_L g4051 ( 
.A(n_3142),
.B(n_3046),
.Y(n_4051)
);

CKINVDCx20_ASAP7_75t_R g4052 ( 
.A(n_3335),
.Y(n_4052)
);

NAND2x1p5_ASAP7_75t_L g4053 ( 
.A(n_3108),
.B(n_3037),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_3436),
.Y(n_4054)
);

BUFx2_ASAP7_75t_SL g4055 ( 
.A(n_3390),
.Y(n_4055)
);

BUFx3_ASAP7_75t_L g4056 ( 
.A(n_3342),
.Y(n_4056)
);

BUFx4_ASAP7_75t_SL g4057 ( 
.A(n_3261),
.Y(n_4057)
);

INVx1_ASAP7_75t_SL g4058 ( 
.A(n_3171),
.Y(n_4058)
);

CKINVDCx20_ASAP7_75t_R g4059 ( 
.A(n_3449),
.Y(n_4059)
);

INVx5_ASAP7_75t_L g4060 ( 
.A(n_3546),
.Y(n_4060)
);

BUFx12f_ASAP7_75t_L g4061 ( 
.A(n_3400),
.Y(n_4061)
);

BUFx2_ASAP7_75t_SL g4062 ( 
.A(n_3390),
.Y(n_4062)
);

INVx4_ASAP7_75t_L g4063 ( 
.A(n_3196),
.Y(n_4063)
);

INVx5_ASAP7_75t_L g4064 ( 
.A(n_3500),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3069),
.A2(n_3525),
.B1(n_3558),
.B2(n_3534),
.Y(n_4065)
);

INVx5_ASAP7_75t_SL g4066 ( 
.A(n_3301),
.Y(n_4066)
);

CKINVDCx20_ASAP7_75t_R g4067 ( 
.A(n_3449),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_3046),
.B(n_3515),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3342),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3226),
.Y(n_4070)
);

INVx3_ASAP7_75t_L g4071 ( 
.A(n_3389),
.Y(n_4071)
);

BUFx4_ASAP7_75t_SL g4072 ( 
.A(n_3261),
.Y(n_4072)
);

INVx5_ASAP7_75t_L g4073 ( 
.A(n_3500),
.Y(n_4073)
);

INVx3_ASAP7_75t_L g4074 ( 
.A(n_3389),
.Y(n_4074)
);

INVx1_ASAP7_75t_SL g4075 ( 
.A(n_3171),
.Y(n_4075)
);

INVx1_ASAP7_75t_SL g4076 ( 
.A(n_3528),
.Y(n_4076)
);

BUFx4f_ASAP7_75t_L g4077 ( 
.A(n_3241),
.Y(n_4077)
);

INVx3_ASAP7_75t_SL g4078 ( 
.A(n_3273),
.Y(n_4078)
);

NAND2x1p5_ASAP7_75t_L g4079 ( 
.A(n_3037),
.B(n_3210),
.Y(n_4079)
);

BUFx12f_ASAP7_75t_L g4080 ( 
.A(n_3428),
.Y(n_4080)
);

INVx3_ASAP7_75t_SL g4081 ( 
.A(n_3196),
.Y(n_4081)
);

CKINVDCx5p33_ASAP7_75t_R g4082 ( 
.A(n_3284),
.Y(n_4082)
);

BUFx3_ASAP7_75t_L g4083 ( 
.A(n_3259),
.Y(n_4083)
);

CKINVDCx20_ASAP7_75t_R g4084 ( 
.A(n_3354),
.Y(n_4084)
);

CKINVDCx8_ASAP7_75t_R g4085 ( 
.A(n_3333),
.Y(n_4085)
);

NAND2x1p5_ASAP7_75t_L g4086 ( 
.A(n_3210),
.B(n_3100),
.Y(n_4086)
);

BUFx12f_ASAP7_75t_L g4087 ( 
.A(n_3428),
.Y(n_4087)
);

CKINVDCx20_ASAP7_75t_R g4088 ( 
.A(n_3354),
.Y(n_4088)
);

CKINVDCx5p33_ASAP7_75t_R g4089 ( 
.A(n_3375),
.Y(n_4089)
);

INVxp67_ASAP7_75t_SL g4090 ( 
.A(n_3521),
.Y(n_4090)
);

OR2x6_ASAP7_75t_L g4091 ( 
.A(n_3111),
.B(n_3110),
.Y(n_4091)
);

NAND2x1p5_ASAP7_75t_L g4092 ( 
.A(n_3100),
.B(n_3170),
.Y(n_4092)
);

NAND2x1_ASAP7_75t_L g4093 ( 
.A(n_3119),
.B(n_3565),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3176),
.B(n_3189),
.Y(n_4094)
);

BUFx4_ASAP7_75t_SL g4095 ( 
.A(n_3446),
.Y(n_4095)
);

AND2x4_ASAP7_75t_L g4096 ( 
.A(n_3096),
.B(n_3104),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3189),
.B(n_3569),
.Y(n_4097)
);

CKINVDCx20_ASAP7_75t_R g4098 ( 
.A(n_3452),
.Y(n_4098)
);

NAND2x1p5_ASAP7_75t_L g4099 ( 
.A(n_3170),
.B(n_3646),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_3046),
.B(n_3515),
.Y(n_4100)
);

NAND2x1p5_ASAP7_75t_L g4101 ( 
.A(n_3646),
.B(n_3093),
.Y(n_4101)
);

NAND2x1p5_ASAP7_75t_L g4102 ( 
.A(n_3093),
.B(n_3094),
.Y(n_4102)
);

BUFx3_ASAP7_75t_L g4103 ( 
.A(n_3426),
.Y(n_4103)
);

BUFx3_ASAP7_75t_L g4104 ( 
.A(n_3426),
.Y(n_4104)
);

INVx1_ASAP7_75t_SL g4105 ( 
.A(n_3569),
.Y(n_4105)
);

BUFx3_ASAP7_75t_L g4106 ( 
.A(n_3426),
.Y(n_4106)
);

BUFx8_ASAP7_75t_L g4107 ( 
.A(n_3145),
.Y(n_4107)
);

INVx5_ASAP7_75t_L g4108 ( 
.A(n_3196),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_3525),
.B(n_3534),
.Y(n_4109)
);

INVx1_ASAP7_75t_SL g4110 ( 
.A(n_3634),
.Y(n_4110)
);

INVx4_ASAP7_75t_L g4111 ( 
.A(n_3320),
.Y(n_4111)
);

BUFx2_ASAP7_75t_SL g4112 ( 
.A(n_3260),
.Y(n_4112)
);

BUFx12f_ASAP7_75t_L g4113 ( 
.A(n_3428),
.Y(n_4113)
);

INVx1_ASAP7_75t_SL g4114 ( 
.A(n_3634),
.Y(n_4114)
);

INVx5_ASAP7_75t_L g4115 ( 
.A(n_3320),
.Y(n_4115)
);

INVx5_ASAP7_75t_L g4116 ( 
.A(n_3320),
.Y(n_4116)
);

AOI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3624),
.A2(n_3482),
.B1(n_3506),
.B2(n_3493),
.Y(n_4117)
);

INVxp67_ASAP7_75t_SL g4118 ( 
.A(n_3522),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_3096),
.B(n_3104),
.Y(n_4119)
);

BUFx2_ASAP7_75t_SL g4120 ( 
.A(n_3260),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_3375),
.Y(n_4121)
);

INVxp67_ASAP7_75t_L g4122 ( 
.A(n_3522),
.Y(n_4122)
);

BUFx2_ASAP7_75t_SL g4123 ( 
.A(n_3205),
.Y(n_4123)
);

BUFx10_ASAP7_75t_L g4124 ( 
.A(n_3256),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3098),
.B(n_3080),
.Y(n_4125)
);

INVx5_ASAP7_75t_L g4126 ( 
.A(n_3320),
.Y(n_4126)
);

BUFx12f_ASAP7_75t_L g4127 ( 
.A(n_3479),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3319),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_SL g4129 ( 
.A1(n_3131),
.A2(n_3112),
.B1(n_3215),
.B2(n_3574),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_3046),
.B(n_3515),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3319),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_3098),
.B(n_3627),
.Y(n_4132)
);

AND2x4_ASAP7_75t_L g4133 ( 
.A(n_3294),
.B(n_3204),
.Y(n_4133)
);

CKINVDCx11_ASAP7_75t_R g4134 ( 
.A(n_3388),
.Y(n_4134)
);

INVx6_ASAP7_75t_SL g4135 ( 
.A(n_3294),
.Y(n_4135)
);

BUFx4_ASAP7_75t_SL g4136 ( 
.A(n_3446),
.Y(n_4136)
);

BUFx2_ASAP7_75t_L g4137 ( 
.A(n_3205),
.Y(n_4137)
);

BUFx12f_ASAP7_75t_L g4138 ( 
.A(n_3235),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3185),
.B(n_3231),
.Y(n_4139)
);

AND2x2_ASAP7_75t_L g4140 ( 
.A(n_3515),
.B(n_3590),
.Y(n_4140)
);

CKINVDCx20_ASAP7_75t_R g4141 ( 
.A(n_3452),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_3235),
.Y(n_4142)
);

CKINVDCx5p33_ASAP7_75t_R g4143 ( 
.A(n_3343),
.Y(n_4143)
);

CKINVDCx16_ASAP7_75t_R g4144 ( 
.A(n_3388),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3185),
.B(n_3231),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_3590),
.B(n_3652),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3207),
.B(n_3209),
.Y(n_4147)
);

CKINVDCx6p67_ASAP7_75t_R g4148 ( 
.A(n_3271),
.Y(n_4148)
);

INVx1_ASAP7_75t_SL g4149 ( 
.A(n_3464),
.Y(n_4149)
);

NAND2x1p5_ASAP7_75t_L g4150 ( 
.A(n_3155),
.B(n_3242),
.Y(n_4150)
);

NAND2x1p5_ASAP7_75t_L g4151 ( 
.A(n_3242),
.B(n_3248),
.Y(n_4151)
);

BUFx2_ASAP7_75t_SL g4152 ( 
.A(n_3378),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3207),
.B(n_3209),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3054),
.B(n_3085),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3054),
.B(n_3085),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3523),
.B(n_3527),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_3267),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3441),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_SL g4159 ( 
.A(n_3558),
.B(n_3559),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3441),
.Y(n_4160)
);

NAND2x1p5_ASAP7_75t_L g4161 ( 
.A(n_3248),
.B(n_3232),
.Y(n_4161)
);

CKINVDCx20_ASAP7_75t_R g4162 ( 
.A(n_3157),
.Y(n_4162)
);

CKINVDCx5p33_ASAP7_75t_R g4163 ( 
.A(n_3152),
.Y(n_4163)
);

BUFx2_ASAP7_75t_SL g4164 ( 
.A(n_3417),
.Y(n_4164)
);

INVxp33_ASAP7_75t_L g4165 ( 
.A(n_3409),
.Y(n_4165)
);

BUFx3_ASAP7_75t_L g4166 ( 
.A(n_3517),
.Y(n_4166)
);

INVx2_ASAP7_75t_SL g4167 ( 
.A(n_3517),
.Y(n_4167)
);

INVx2_ASAP7_75t_SL g4168 ( 
.A(n_3530),
.Y(n_4168)
);

NAND2x1p5_ASAP7_75t_L g4169 ( 
.A(n_3232),
.B(n_3200),
.Y(n_4169)
);

INVx2_ASAP7_75t_SL g4170 ( 
.A(n_3530),
.Y(n_4170)
);

CKINVDCx6p67_ASAP7_75t_R g4171 ( 
.A(n_3523),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_3527),
.B(n_3531),
.Y(n_4172)
);

INVx3_ASAP7_75t_L g4173 ( 
.A(n_3266),
.Y(n_4173)
);

BUFx2_ASAP7_75t_R g4174 ( 
.A(n_3372),
.Y(n_4174)
);

BUFx2_ASAP7_75t_L g4175 ( 
.A(n_3227),
.Y(n_4175)
);

CKINVDCx14_ASAP7_75t_R g4176 ( 
.A(n_3203),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_3590),
.B(n_3652),
.Y(n_4177)
);

BUFx4_ASAP7_75t_SL g4178 ( 
.A(n_3460),
.Y(n_4178)
);

BUFx2_ASAP7_75t_L g4179 ( 
.A(n_3227),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3590),
.B(n_3652),
.Y(n_4180)
);

AOI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_3550),
.A2(n_3632),
.B1(n_3647),
.B2(n_3562),
.Y(n_4181)
);

BUFx2_ASAP7_75t_L g4182 ( 
.A(n_3369),
.Y(n_4182)
);

BUFx6f_ASAP7_75t_L g4183 ( 
.A(n_3083),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3531),
.B(n_3544),
.Y(n_4184)
);

CKINVDCx5p33_ASAP7_75t_R g4185 ( 
.A(n_3377),
.Y(n_4185)
);

INVxp67_ASAP7_75t_SL g4186 ( 
.A(n_3544),
.Y(n_4186)
);

INVxp33_ASAP7_75t_SL g4187 ( 
.A(n_3658),
.Y(n_4187)
);

BUFx4f_ASAP7_75t_SL g4188 ( 
.A(n_3380),
.Y(n_4188)
);

AND2x4_ASAP7_75t_L g4189 ( 
.A(n_3158),
.B(n_3127),
.Y(n_4189)
);

OR2x6_ASAP7_75t_L g4190 ( 
.A(n_3119),
.B(n_3384),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_3360),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3360),
.Y(n_4192)
);

CKINVDCx20_ASAP7_75t_R g4193 ( 
.A(n_3157),
.Y(n_4193)
);

OR2x6_ASAP7_75t_L g4194 ( 
.A(n_3078),
.B(n_3122),
.Y(n_4194)
);

BUFx2_ASAP7_75t_L g4195 ( 
.A(n_3369),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3590),
.B(n_3652),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_4122),
.B(n_3066),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_3832),
.Y(n_4198)
);

BUFx2_ASAP7_75t_R g4199 ( 
.A(n_3761),
.Y(n_4199)
);

AO31x2_ASAP7_75t_L g4200 ( 
.A1(n_3987),
.A2(n_3501),
.A3(n_3043),
.B(n_3048),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_3691),
.Y(n_4201)
);

A2O1A1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_4093),
.A2(n_3778),
.B(n_3800),
.C(n_3813),
.Y(n_4202)
);

OAI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_4065),
.A2(n_3044),
.B(n_3559),
.Y(n_4203)
);

AOI21x1_ASAP7_75t_L g4204 ( 
.A1(n_3820),
.A2(n_3662),
.B(n_3643),
.Y(n_4204)
);

AO21x2_ASAP7_75t_L g4205 ( 
.A1(n_3987),
.A2(n_3579),
.B(n_3577),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_3813),
.A2(n_3131),
.B1(n_3605),
.B2(n_3587),
.Y(n_4206)
);

OAI21xp5_ASAP7_75t_L g4207 ( 
.A1(n_4065),
.A2(n_3605),
.B(n_3587),
.Y(n_4207)
);

AO21x2_ASAP7_75t_L g4208 ( 
.A1(n_3990),
.A2(n_3579),
.B(n_3577),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_4163),
.B(n_3385),
.Y(n_4209)
);

A2O1A1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_4093),
.A2(n_3800),
.B(n_3778),
.C(n_3701),
.Y(n_4210)
);

AOI221xp5_ASAP7_75t_L g4211 ( 
.A1(n_3745),
.A2(n_3580),
.B1(n_3621),
.B2(n_3592),
.C(n_3628),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_3832),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3691),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_3832),
.Y(n_4214)
);

OAI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_3926),
.A2(n_4117),
.B1(n_4181),
.B2(n_3904),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4122),
.B(n_3066),
.Y(n_4216)
);

NOR2xp33_ASAP7_75t_L g4217 ( 
.A(n_4187),
.B(n_3118),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3672),
.Y(n_4218)
);

AOI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_3745),
.A2(n_3628),
.B1(n_3648),
.B2(n_3639),
.Y(n_4219)
);

BUFx2_ASAP7_75t_L g4220 ( 
.A(n_3697),
.Y(n_4220)
);

OAI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_3926),
.A2(n_3648),
.B(n_3639),
.Y(n_4221)
);

OR2x2_ASAP7_75t_L g4222 ( 
.A(n_4058),
.B(n_3652),
.Y(n_4222)
);

INVx5_ASAP7_75t_L g4223 ( 
.A(n_4190),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_3873),
.B(n_4021),
.Y(n_4224)
);

BUFx2_ASAP7_75t_L g4225 ( 
.A(n_3697),
.Y(n_4225)
);

BUFx3_ASAP7_75t_L g4226 ( 
.A(n_3694),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_3873),
.B(n_3145),
.Y(n_4227)
);

AND2x2_ASAP7_75t_L g4228 ( 
.A(n_3873),
.B(n_3136),
.Y(n_4228)
);

AOI22xp5_ASAP7_75t_L g4229 ( 
.A1(n_3819),
.A2(n_3604),
.B1(n_3574),
.B2(n_3516),
.Y(n_4229)
);

OAI21x1_ASAP7_75t_L g4230 ( 
.A1(n_4029),
.A2(n_3603),
.B(n_3063),
.Y(n_4230)
);

INVx4_ASAP7_75t_L g4231 ( 
.A(n_3711),
.Y(n_4231)
);

A2O1A1Ixp33_ASAP7_75t_L g4232 ( 
.A1(n_3701),
.A2(n_3123),
.B(n_3101),
.C(n_3172),
.Y(n_4232)
);

CKINVDCx5p33_ASAP7_75t_R g4233 ( 
.A(n_3762),
.Y(n_4233)
);

OAI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4109),
.A2(n_3649),
.B(n_3580),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_3672),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3678),
.Y(n_4236)
);

OAI21x1_ASAP7_75t_L g4237 ( 
.A1(n_4029),
.A2(n_3603),
.B(n_3481),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3678),
.Y(n_4238)
);

OAI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_4159),
.A2(n_3649),
.B(n_3662),
.Y(n_4239)
);

BUFx6f_ASAP7_75t_L g4240 ( 
.A(n_3689),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3939),
.B(n_3548),
.Y(n_4241)
);

OAI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4117),
.A2(n_3220),
.B1(n_3215),
.B2(n_3112),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_4091),
.A2(n_3484),
.B(n_3040),
.Y(n_4243)
);

AOI31xp67_ASAP7_75t_L g4244 ( 
.A1(n_4181),
.A2(n_3496),
.A3(n_3557),
.B(n_3547),
.Y(n_4244)
);

OAI21x1_ASAP7_75t_L g4245 ( 
.A1(n_4169),
.A2(n_3499),
.B(n_3485),
.Y(n_4245)
);

OR2x6_ASAP7_75t_L g4246 ( 
.A(n_3689),
.B(n_3509),
.Y(n_4246)
);

INVx3_ASAP7_75t_L g4247 ( 
.A(n_3775),
.Y(n_4247)
);

AND2x4_ASAP7_75t_L g4248 ( 
.A(n_3681),
.B(n_3477),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_3858),
.Y(n_4249)
);

OAI21x1_ASAP7_75t_L g4250 ( 
.A1(n_4169),
.A2(n_3520),
.B(n_3511),
.Y(n_4250)
);

OAI21x1_ASAP7_75t_L g4251 ( 
.A1(n_4169),
.A2(n_3540),
.B(n_3533),
.Y(n_4251)
);

BUFx2_ASAP7_75t_L g4252 ( 
.A(n_3697),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3686),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_3858),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3686),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3939),
.B(n_3548),
.Y(n_4256)
);

OAI22xp5_ASAP7_75t_L g4257 ( 
.A1(n_3819),
.A2(n_3124),
.B1(n_3592),
.B2(n_3087),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_3858),
.Y(n_4258)
);

AOI22xp33_ASAP7_75t_L g4259 ( 
.A1(n_3932),
.A2(n_4020),
.B1(n_3972),
.B2(n_3914),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3698),
.Y(n_4260)
);

OAI21x1_ASAP7_75t_L g4261 ( 
.A1(n_4169),
.A2(n_3606),
.B(n_3568),
.Y(n_4261)
);

OAI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_3932),
.A2(n_3220),
.B1(n_3150),
.B2(n_3480),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_3859),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_3859),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4156),
.B(n_3549),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_3859),
.Y(n_4266)
);

OAI21x1_ASAP7_75t_L g4267 ( 
.A1(n_4092),
.A2(n_3641),
.B(n_3626),
.Y(n_4267)
);

NAND2x1p5_ASAP7_75t_L g4268 ( 
.A(n_3681),
.B(n_3696),
.Y(n_4268)
);

NAND2x1_ASAP7_75t_L g4269 ( 
.A(n_4190),
.B(n_3057),
.Y(n_4269)
);

INVx3_ASAP7_75t_L g4270 ( 
.A(n_3775),
.Y(n_4270)
);

INVx1_ASAP7_75t_SL g4271 ( 
.A(n_3814),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4021),
.B(n_3144),
.Y(n_4272)
);

AOI21xp5_ASAP7_75t_L g4273 ( 
.A1(n_4091),
.A2(n_3656),
.B(n_3644),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4021),
.B(n_3144),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_3883),
.Y(n_4275)
);

O2A1O1Ixp33_ASAP7_75t_SL g4276 ( 
.A1(n_3934),
.A2(n_3392),
.B(n_3513),
.C(n_3495),
.Y(n_4276)
);

INVx1_ASAP7_75t_SL g4277 ( 
.A(n_3814),
.Y(n_4277)
);

OAI22xp5_ASAP7_75t_L g4278 ( 
.A1(n_3914),
.A2(n_3514),
.B1(n_3535),
.B2(n_3524),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4156),
.B(n_4172),
.Y(n_4279)
);

BUFx6f_ASAP7_75t_L g4280 ( 
.A(n_3689),
.Y(n_4280)
);

AOI22xp33_ASAP7_75t_L g4281 ( 
.A1(n_3972),
.A2(n_3621),
.B1(n_3138),
.B2(n_3501),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_R g4282 ( 
.A(n_3699),
.B(n_3221),
.Y(n_4282)
);

INVx2_ASAP7_75t_SL g4283 ( 
.A(n_4060),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3698),
.Y(n_4284)
);

NOR2xp67_ASAP7_75t_SL g4285 ( 
.A(n_3771),
.B(n_3565),
.Y(n_4285)
);

OAI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4020),
.A2(n_3661),
.B(n_3545),
.Y(n_4286)
);

BUFx2_ASAP7_75t_SL g4287 ( 
.A(n_3777),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_3883),
.Y(n_4288)
);

INVx2_ASAP7_75t_SL g4289 ( 
.A(n_4060),
.Y(n_4289)
);

NOR2xp33_ASAP7_75t_L g4290 ( 
.A(n_4143),
.B(n_3118),
.Y(n_4290)
);

AOI21x1_ASAP7_75t_L g4291 ( 
.A1(n_3967),
.A2(n_3268),
.B(n_3658),
.Y(n_4291)
);

NAND2xp33_ASAP7_75t_L g4292 ( 
.A(n_3967),
.B(n_3552),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4172),
.B(n_3549),
.Y(n_4293)
);

AO21x2_ASAP7_75t_L g4294 ( 
.A1(n_4191),
.A2(n_3056),
.B(n_3146),
.Y(n_4294)
);

NAND2x1_ASAP7_75t_L g4295 ( 
.A(n_4190),
.B(n_3720),
.Y(n_4295)
);

OAI22xp5_ASAP7_75t_L g4296 ( 
.A1(n_3967),
.A2(n_3561),
.B1(n_3576),
.B2(n_3573),
.Y(n_4296)
);

INVx2_ASAP7_75t_SL g4297 ( 
.A(n_4060),
.Y(n_4297)
);

OAI21x1_ASAP7_75t_L g4298 ( 
.A1(n_4092),
.A2(n_3067),
.B(n_3060),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4053),
.A2(n_3067),
.B(n_3060),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3700),
.Y(n_4300)
);

AO21x2_ASAP7_75t_L g4301 ( 
.A1(n_4191),
.A2(n_3056),
.B(n_3146),
.Y(n_4301)
);

OAI21x1_ASAP7_75t_L g4302 ( 
.A1(n_4053),
.A2(n_3491),
.B(n_3487),
.Y(n_4302)
);

INVx3_ASAP7_75t_L g4303 ( 
.A(n_3775),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4040),
.B(n_3285),
.Y(n_4304)
);

HB1xp67_ASAP7_75t_L g4305 ( 
.A(n_3705),
.Y(n_4305)
);

AOI22xp33_ASAP7_75t_L g4306 ( 
.A1(n_3967),
.A2(n_4129),
.B1(n_3875),
.B2(n_3138),
.Y(n_4306)
);

BUFx3_ASAP7_75t_L g4307 ( 
.A(n_3694),
.Y(n_4307)
);

INVx3_ASAP7_75t_L g4308 ( 
.A(n_3821),
.Y(n_4308)
);

OAI21x1_ASAP7_75t_L g4309 ( 
.A1(n_4053),
.A2(n_3491),
.B(n_3487),
.Y(n_4309)
);

BUFx3_ASAP7_75t_L g4310 ( 
.A(n_3694),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4040),
.B(n_3285),
.Y(n_4311)
);

OAI21x1_ASAP7_75t_L g4312 ( 
.A1(n_4053),
.A2(n_3508),
.B(n_3498),
.Y(n_4312)
);

INVx3_ASAP7_75t_L g4313 ( 
.A(n_3821),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_3700),
.Y(n_4314)
);

INVxp67_ASAP7_75t_L g4315 ( 
.A(n_3685),
.Y(n_4315)
);

AOI21xp5_ASAP7_75t_L g4316 ( 
.A1(n_4091),
.A2(n_3553),
.B(n_3551),
.Y(n_4316)
);

BUFx6f_ASAP7_75t_L g4317 ( 
.A(n_3689),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3703),
.Y(n_4318)
);

AOI22xp33_ASAP7_75t_L g4319 ( 
.A1(n_3967),
.A2(n_3114),
.B1(n_3121),
.B2(n_3105),
.Y(n_4319)
);

OAI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4129),
.A2(n_3097),
.B(n_3174),
.Y(n_4320)
);

BUFx3_ASAP7_75t_L g4321 ( 
.A(n_3694),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_3697),
.Y(n_4322)
);

NAND3xp33_ASAP7_75t_SL g4323 ( 
.A(n_3875),
.B(n_3193),
.C(n_3589),
.Y(n_4323)
);

CKINVDCx11_ASAP7_75t_R g4324 ( 
.A(n_3727),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_3703),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_3708),
.Y(n_4326)
);

BUFx2_ASAP7_75t_L g4327 ( 
.A(n_3697),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4184),
.B(n_3551),
.Y(n_4328)
);

OAI22xp5_ASAP7_75t_L g4329 ( 
.A1(n_3904),
.A2(n_3637),
.B1(n_3665),
.B2(n_3640),
.Y(n_4329)
);

O2A1O1Ixp33_ASAP7_75t_SL g4330 ( 
.A1(n_4057),
.A2(n_3129),
.B(n_3140),
.C(n_3338),
.Y(n_4330)
);

HB1xp67_ASAP7_75t_L g4331 ( 
.A(n_3705),
.Y(n_4331)
);

AOI222xp33_ASAP7_75t_L g4332 ( 
.A1(n_4154),
.A2(n_3114),
.B1(n_3105),
.B2(n_3121),
.C1(n_3130),
.C2(n_3193),
.Y(n_4332)
);

AOI21xp5_ASAP7_75t_L g4333 ( 
.A1(n_4091),
.A2(n_3554),
.B(n_3553),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_3708),
.Y(n_4334)
);

AOI21xp5_ASAP7_75t_R g4335 ( 
.A1(n_4057),
.A2(n_3130),
.B(n_3336),
.Y(n_4335)
);

OAI21x1_ASAP7_75t_L g4336 ( 
.A1(n_4086),
.A2(n_3556),
.B(n_3539),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4040),
.B(n_3285),
.Y(n_4337)
);

BUFx3_ASAP7_75t_L g4338 ( 
.A(n_3694),
.Y(n_4338)
);

AOI21xp33_ASAP7_75t_L g4339 ( 
.A1(n_4154),
.A2(n_3567),
.B(n_3554),
.Y(n_4339)
);

BUFx6f_ASAP7_75t_L g4340 ( 
.A(n_3734),
.Y(n_4340)
);

INVx8_ASAP7_75t_L g4341 ( 
.A(n_3771),
.Y(n_4341)
);

AND2x4_ASAP7_75t_L g4342 ( 
.A(n_3681),
.B(n_3477),
.Y(n_4342)
);

INVx1_ASAP7_75t_SL g4343 ( 
.A(n_3816),
.Y(n_4343)
);

BUFx6f_ASAP7_75t_L g4344 ( 
.A(n_3734),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4041),
.B(n_3786),
.Y(n_4345)
);

AOI22xp33_ASAP7_75t_SL g4346 ( 
.A1(n_4144),
.A2(n_4121),
.B1(n_4089),
.B2(n_4050),
.Y(n_4346)
);

OAI221xp5_ASAP7_75t_L g4347 ( 
.A1(n_4155),
.A2(n_3182),
.B1(n_3089),
.B2(n_3222),
.C(n_3175),
.Y(n_4347)
);

OAI22xp5_ASAP7_75t_L g4348 ( 
.A1(n_3964),
.A2(n_3140),
.B1(n_3129),
.B2(n_3609),
.Y(n_4348)
);

OAI21x1_ASAP7_75t_L g4349 ( 
.A1(n_4086),
.A2(n_3578),
.B(n_3572),
.Y(n_4349)
);

HB1xp67_ASAP7_75t_L g4350 ( 
.A(n_3705),
.Y(n_4350)
);

OAI21x1_ASAP7_75t_L g4351 ( 
.A1(n_4086),
.A2(n_4034),
.B(n_4071),
.Y(n_4351)
);

NAND2xp33_ASAP7_75t_L g4352 ( 
.A(n_3733),
.B(n_3439),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_4086),
.A2(n_3578),
.B(n_3572),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3716),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3716),
.Y(n_4355)
);

OR2x6_ASAP7_75t_L g4356 ( 
.A(n_3734),
.B(n_3133),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4041),
.B(n_3285),
.Y(n_4357)
);

AND2x4_ASAP7_75t_L g4358 ( 
.A(n_3681),
.B(n_3477),
.Y(n_4358)
);

AO21x1_ASAP7_75t_L g4359 ( 
.A1(n_4155),
.A2(n_3265),
.B(n_3206),
.Y(n_4359)
);

O2A1O1Ixp5_ASAP7_75t_L g4360 ( 
.A1(n_4147),
.A2(n_3188),
.B(n_3191),
.C(n_3190),
.Y(n_4360)
);

OAI21x1_ASAP7_75t_L g4361 ( 
.A1(n_4034),
.A2(n_4074),
.B(n_4071),
.Y(n_4361)
);

INVxp33_ASAP7_75t_L g4362 ( 
.A(n_3874),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_3891),
.Y(n_4363)
);

INVx4_ASAP7_75t_SL g4364 ( 
.A(n_3720),
.Y(n_4364)
);

AOI21x1_ASAP7_75t_L g4365 ( 
.A1(n_4147),
.A2(n_3268),
.B(n_3494),
.Y(n_4365)
);

NAND2x1p5_ASAP7_75t_L g4366 ( 
.A(n_3681),
.B(n_3386),
.Y(n_4366)
);

NAND2x1p5_ASAP7_75t_L g4367 ( 
.A(n_3681),
.B(n_3386),
.Y(n_4367)
);

INVx3_ASAP7_75t_L g4368 ( 
.A(n_3821),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3731),
.Y(n_4369)
);

AND2x4_ASAP7_75t_L g4370 ( 
.A(n_3696),
.B(n_3477),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_3731),
.Y(n_4371)
);

INVx4_ASAP7_75t_SL g4372 ( 
.A(n_3720),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_3891),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_4041),
.B(n_3285),
.Y(n_4374)
);

OAI21xp5_ASAP7_75t_L g4375 ( 
.A1(n_4153),
.A2(n_3609),
.B(n_3575),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_3733),
.A2(n_3336),
.B1(n_3510),
.B2(n_3057),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_3903),
.Y(n_4377)
);

INVx1_ASAP7_75t_SL g4378 ( 
.A(n_3816),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_3786),
.B(n_3477),
.Y(n_4379)
);

OAI21x1_ASAP7_75t_L g4380 ( 
.A1(n_4102),
.A2(n_4173),
.B(n_3657),
.Y(n_4380)
);

O2A1O1Ixp33_ASAP7_75t_L g4381 ( 
.A1(n_4153),
.A2(n_3182),
.B(n_3223),
.C(n_3510),
.Y(n_4381)
);

INVxp67_ASAP7_75t_L g4382 ( 
.A(n_3685),
.Y(n_4382)
);

AOI22xp5_ASAP7_75t_L g4383 ( 
.A1(n_4144),
.A2(n_3289),
.B1(n_3286),
.B2(n_3396),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_3744),
.Y(n_4384)
);

AOI221xp5_ASAP7_75t_L g4385 ( 
.A1(n_3752),
.A2(n_3289),
.B1(n_3305),
.B2(n_3310),
.C(n_3567),
.Y(n_4385)
);

AND2x4_ASAP7_75t_L g4386 ( 
.A(n_3696),
.B(n_3477),
.Y(n_4386)
);

OAI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_4182),
.A2(n_3601),
.B(n_3575),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3744),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_3750),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_3903),
.Y(n_4390)
);

INVx3_ASAP7_75t_L g4391 ( 
.A(n_3823),
.Y(n_4391)
);

BUFx12f_ASAP7_75t_L g4392 ( 
.A(n_3771),
.Y(n_4392)
);

INVx2_ASAP7_75t_SL g4393 ( 
.A(n_4060),
.Y(n_4393)
);

HB1xp67_ASAP7_75t_L g4394 ( 
.A(n_4011),
.Y(n_4394)
);

NAND2x1p5_ASAP7_75t_L g4395 ( 
.A(n_3696),
.B(n_3200),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_4091),
.A2(n_3602),
.B(n_3601),
.Y(n_4396)
);

INVx2_ASAP7_75t_SL g4397 ( 
.A(n_4060),
.Y(n_4397)
);

NOR4xp25_ASAP7_75t_L g4398 ( 
.A(n_4072),
.B(n_3305),
.C(n_3310),
.D(n_3602),
.Y(n_4398)
);

BUFx3_ASAP7_75t_L g4399 ( 
.A(n_3774),
.Y(n_4399)
);

OAI21x1_ASAP7_75t_L g4400 ( 
.A1(n_4173),
.A2(n_3668),
.B(n_3148),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4184),
.B(n_3610),
.Y(n_4401)
);

INVx5_ASAP7_75t_L g4402 ( 
.A(n_4190),
.Y(n_4402)
);

OAI22xp5_ASAP7_75t_L g4403 ( 
.A1(n_3964),
.A2(n_3194),
.B1(n_3208),
.B2(n_3195),
.Y(n_4403)
);

AOI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4091),
.A2(n_3611),
.B(n_3610),
.Y(n_4404)
);

AOI21xp5_ASAP7_75t_L g4405 ( 
.A1(n_4190),
.A2(n_3615),
.B(n_3611),
.Y(n_4405)
);

INVx2_ASAP7_75t_SL g4406 ( 
.A(n_4060),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_3723),
.B(n_3615),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_3723),
.B(n_3642),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_L g4409 ( 
.A(n_4165),
.B(n_3412),
.Y(n_4409)
);

OA21x2_ASAP7_75t_L g4410 ( 
.A1(n_4068),
.A2(n_3269),
.B(n_3270),
.Y(n_4410)
);

OR2x6_ASAP7_75t_L g4411 ( 
.A(n_3734),
.B(n_3382),
.Y(n_4411)
);

INVx4_ASAP7_75t_SL g4412 ( 
.A(n_3720),
.Y(n_4412)
);

INVx3_ASAP7_75t_L g4413 ( 
.A(n_3823),
.Y(n_4413)
);

INVx1_ASAP7_75t_SL g4414 ( 
.A(n_3843),
.Y(n_4414)
);

CKINVDCx6p67_ASAP7_75t_R g4415 ( 
.A(n_3774),
.Y(n_4415)
);

INVx3_ASAP7_75t_L g4416 ( 
.A(n_3823),
.Y(n_4416)
);

NOR2xp33_ASAP7_75t_L g4417 ( 
.A(n_4004),
.B(n_3394),
.Y(n_4417)
);

OAI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_4182),
.A2(n_3645),
.B(n_3642),
.Y(n_4418)
);

OAI21x1_ASAP7_75t_SL g4419 ( 
.A1(n_3677),
.A2(n_3297),
.B(n_3246),
.Y(n_4419)
);

CKINVDCx5p33_ASAP7_75t_R g4420 ( 
.A(n_3826),
.Y(n_4420)
);

INVx3_ASAP7_75t_L g4421 ( 
.A(n_3836),
.Y(n_4421)
);

BUFx12f_ASAP7_75t_L g4422 ( 
.A(n_3774),
.Y(n_4422)
);

OAI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_4195),
.A2(n_3651),
.B(n_3645),
.Y(n_4423)
);

OAI21x1_ASAP7_75t_L g4424 ( 
.A1(n_4046),
.A2(n_3177),
.B(n_3494),
.Y(n_4424)
);

AO32x2_ASAP7_75t_L g4425 ( 
.A1(n_4043),
.A2(n_3415),
.A3(n_3410),
.B1(n_3396),
.B2(n_3079),
.Y(n_4425)
);

OR2x6_ASAP7_75t_L g4426 ( 
.A(n_3741),
.B(n_3277),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_L g4427 ( 
.A1(n_3733),
.A2(n_3625),
.B1(n_3238),
.B2(n_3415),
.Y(n_4427)
);

O2A1O1Ixp33_ASAP7_75t_SL g4428 ( 
.A1(n_4072),
.A2(n_3471),
.B(n_3296),
.C(n_3306),
.Y(n_4428)
);

AND2x4_ASAP7_75t_L g4429 ( 
.A(n_3696),
.B(n_3739),
.Y(n_4429)
);

INVx8_ASAP7_75t_L g4430 ( 
.A(n_3792),
.Y(n_4430)
);

OAI21xp5_ASAP7_75t_L g4431 ( 
.A1(n_4195),
.A2(n_3653),
.B(n_3651),
.Y(n_4431)
);

AOI22xp5_ASAP7_75t_L g4432 ( 
.A1(n_4059),
.A2(n_3286),
.B1(n_3410),
.B2(n_3238),
.Y(n_4432)
);

OA21x2_ASAP7_75t_L g4433 ( 
.A1(n_4068),
.A2(n_4140),
.B(n_4100),
.Y(n_4433)
);

OAI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_3752),
.A2(n_3655),
.B(n_3653),
.Y(n_4434)
);

INVx3_ASAP7_75t_SL g4435 ( 
.A(n_4171),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_3729),
.B(n_3655),
.Y(n_4436)
);

AOI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4067),
.A2(n_3424),
.B1(n_3387),
.B2(n_3301),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_3763),
.Y(n_4438)
);

AOI21x1_ASAP7_75t_L g4439 ( 
.A1(n_4192),
.A2(n_3600),
.B(n_3536),
.Y(n_4439)
);

AOI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_4190),
.A2(n_3669),
.B(n_3625),
.Y(n_4440)
);

AO21x2_ASAP7_75t_L g4441 ( 
.A1(n_4192),
.A2(n_4100),
.B(n_4068),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_3786),
.B(n_3092),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_L g4443 ( 
.A1(n_3743),
.A2(n_3333),
.B1(n_3297),
.B2(n_3381),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_3729),
.B(n_3669),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3765),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_3765),
.Y(n_4446)
);

OA21x2_ASAP7_75t_L g4447 ( 
.A1(n_4140),
.A2(n_3269),
.B(n_3240),
.Y(n_4447)
);

OAI21xp5_ASAP7_75t_L g4448 ( 
.A1(n_4175),
.A2(n_3351),
.B(n_3240),
.Y(n_4448)
);

OR2x2_ASAP7_75t_L g4449 ( 
.A(n_4058),
.B(n_3079),
.Y(n_4449)
);

INVxp33_ASAP7_75t_L g4450 ( 
.A(n_4134),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_3758),
.B(n_3692),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_3834),
.B(n_3092),
.Y(n_4452)
);

OAI21x1_ASAP7_75t_L g4453 ( 
.A1(n_4161),
.A2(n_4099),
.B(n_4101),
.Y(n_4453)
);

INVx1_ASAP7_75t_SL g4454 ( 
.A(n_3843),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_3834),
.B(n_3092),
.Y(n_4455)
);

NOR2x1_ASAP7_75t_L g4456 ( 
.A(n_3725),
.B(n_3331),
.Y(n_4456)
);

OAI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_4175),
.A2(n_3163),
.B(n_3224),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_3768),
.Y(n_4458)
);

INVx3_ASAP7_75t_L g4459 ( 
.A(n_3836),
.Y(n_4459)
);

NOR2xp33_ASAP7_75t_SL g4460 ( 
.A(n_3712),
.B(n_3462),
.Y(n_4460)
);

INVx2_ASAP7_75t_SL g4461 ( 
.A(n_4060),
.Y(n_4461)
);

AOI22xp33_ASAP7_75t_L g4462 ( 
.A1(n_3743),
.A2(n_3381),
.B1(n_3180),
.B2(n_3397),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_3758),
.B(n_3090),
.Y(n_4463)
);

BUFx6f_ASAP7_75t_L g4464 ( 
.A(n_3741),
.Y(n_4464)
);

OAI21x1_ASAP7_75t_L g4465 ( 
.A1(n_4101),
.A2(n_3276),
.B(n_3254),
.Y(n_4465)
);

OAI21x1_ASAP7_75t_SL g4466 ( 
.A1(n_3677),
.A2(n_3246),
.B(n_3180),
.Y(n_4466)
);

AND2x4_ASAP7_75t_L g4467 ( 
.A(n_3739),
.B(n_3414),
.Y(n_4467)
);

OAI21x1_ASAP7_75t_L g4468 ( 
.A1(n_4101),
.A2(n_3254),
.B(n_3245),
.Y(n_4468)
);

CKINVDCx11_ASAP7_75t_R g4469 ( 
.A(n_3757),
.Y(n_4469)
);

OAI21x1_ASAP7_75t_L g4470 ( 
.A1(n_4101),
.A2(n_4079),
.B(n_4150),
.Y(n_4470)
);

BUFx3_ASAP7_75t_L g4471 ( 
.A(n_3792),
.Y(n_4471)
);

INVx4_ASAP7_75t_SL g4472 ( 
.A(n_3720),
.Y(n_4472)
);

BUFx10_ASAP7_75t_L g4473 ( 
.A(n_3738),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_4079),
.A2(n_3245),
.B(n_3272),
.Y(n_4474)
);

BUFx2_ASAP7_75t_SL g4475 ( 
.A(n_4064),
.Y(n_4475)
);

CKINVDCx20_ASAP7_75t_R g4476 ( 
.A(n_3759),
.Y(n_4476)
);

AOI22xp33_ASAP7_75t_L g4477 ( 
.A1(n_3743),
.A2(n_3413),
.B1(n_3383),
.B2(n_3427),
.Y(n_4477)
);

AND2x4_ASAP7_75t_L g4478 ( 
.A(n_3739),
.B(n_3327),
.Y(n_4478)
);

OAI21xp5_ASAP7_75t_L g4479 ( 
.A1(n_4179),
.A2(n_3163),
.B(n_3349),
.Y(n_4479)
);

NAND2x1p5_ASAP7_75t_L g4480 ( 
.A(n_3739),
.B(n_3127),
.Y(n_4480)
);

BUFx3_ASAP7_75t_L g4481 ( 
.A(n_3792),
.Y(n_4481)
);

INVx2_ASAP7_75t_SL g4482 ( 
.A(n_3836),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_3692),
.B(n_3090),
.Y(n_4483)
);

OAI21xp5_ASAP7_75t_L g4484 ( 
.A1(n_4179),
.A2(n_3314),
.B(n_3234),
.Y(n_4484)
);

OAI21xp5_ASAP7_75t_L g4485 ( 
.A1(n_4194),
.A2(n_3275),
.B(n_3274),
.Y(n_4485)
);

OAI21xp5_ASAP7_75t_L g4486 ( 
.A1(n_4194),
.A2(n_3295),
.B(n_3328),
.Y(n_4486)
);

AOI21xp5_ASAP7_75t_L g4487 ( 
.A1(n_4194),
.A2(n_3468),
.B(n_3321),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_3779),
.Y(n_4488)
);

INVx1_ASAP7_75t_SL g4489 ( 
.A(n_3853),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_3779),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_3794),
.Y(n_4491)
);

AND2x4_ASAP7_75t_L g4492 ( 
.A(n_3739),
.B(n_3767),
.Y(n_4492)
);

AND2x4_ASAP7_75t_L g4493 ( 
.A(n_3739),
.B(n_3327),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4194),
.A2(n_3325),
.B(n_3330),
.Y(n_4494)
);

INVx1_ASAP7_75t_SL g4495 ( 
.A(n_3853),
.Y(n_4495)
);

A2O1A1Ixp33_ASAP7_75t_L g4496 ( 
.A1(n_3964),
.A2(n_3332),
.B(n_3334),
.C(n_3312),
.Y(n_4496)
);

OAI21x1_ASAP7_75t_SL g4497 ( 
.A1(n_3677),
.A2(n_3309),
.B(n_3316),
.Y(n_4497)
);

BUFx2_ASAP7_75t_L g4498 ( 
.A(n_3996),
.Y(n_4498)
);

INVx5_ASAP7_75t_SL g4499 ( 
.A(n_4171),
.Y(n_4499)
);

OR2x6_ASAP7_75t_L g4500 ( 
.A(n_3741),
.B(n_3187),
.Y(n_4500)
);

OAI21xp5_ASAP7_75t_L g4501 ( 
.A1(n_4194),
.A2(n_3324),
.B(n_3309),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_3794),
.Y(n_4502)
);

INVx2_ASAP7_75t_SL g4503 ( 
.A(n_4064),
.Y(n_4503)
);

AOI22xp33_ASAP7_75t_L g4504 ( 
.A1(n_3769),
.A2(n_4050),
.B1(n_4077),
.B2(n_3964),
.Y(n_4504)
);

AOI22xp33_ASAP7_75t_L g4505 ( 
.A1(n_3769),
.A2(n_3383),
.B1(n_3416),
.B2(n_3324),
.Y(n_4505)
);

OAI21x1_ASAP7_75t_SL g4506 ( 
.A1(n_3677),
.A2(n_3316),
.B(n_3433),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_3751),
.B(n_3090),
.Y(n_4507)
);

O2A1O1Ixp33_ASAP7_75t_L g4508 ( 
.A1(n_3769),
.A2(n_3194),
.B(n_3195),
.C(n_3208),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_3795),
.Y(n_4509)
);

OAI21x1_ASAP7_75t_L g4510 ( 
.A1(n_4028),
.A2(n_3262),
.B(n_3406),
.Y(n_4510)
);

O2A1O1Ixp33_ASAP7_75t_SL g4511 ( 
.A1(n_3782),
.A2(n_3437),
.B(n_3212),
.C(n_3225),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_3751),
.B(n_3090),
.Y(n_4512)
);

OAI21x1_ASAP7_75t_L g4513 ( 
.A1(n_4028),
.A2(n_3264),
.B(n_3263),
.Y(n_4513)
);

O2A1O1Ixp33_ASAP7_75t_SL g4514 ( 
.A1(n_3712),
.A2(n_3212),
.B(n_3225),
.C(n_3313),
.Y(n_4514)
);

AOI22xp33_ASAP7_75t_L g4515 ( 
.A1(n_4050),
.A2(n_3318),
.B1(n_3166),
.B2(n_3664),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_R g4516 ( 
.A(n_4009),
.B(n_3747),
.Y(n_4516)
);

AOI21xp5_ASAP7_75t_L g4517 ( 
.A1(n_4194),
.A2(n_3470),
.B(n_3403),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_3795),
.Y(n_4518)
);

BUFx2_ASAP7_75t_L g4519 ( 
.A(n_3996),
.Y(n_4519)
);

HB1xp67_ASAP7_75t_L g4520 ( 
.A(n_3841),
.Y(n_4520)
);

BUFx3_ASAP7_75t_L g4521 ( 
.A(n_3799),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_3824),
.B(n_3090),
.Y(n_4522)
);

OAI22xp5_ASAP7_75t_L g4523 ( 
.A1(n_4050),
.A2(n_3243),
.B1(n_3252),
.B2(n_3249),
.Y(n_4523)
);

AO22x1_ASAP7_75t_L g4524 ( 
.A1(n_3776),
.A2(n_3466),
.B1(n_3463),
.B2(n_3401),
.Y(n_4524)
);

NAND2x1p5_ASAP7_75t_L g4525 ( 
.A(n_3767),
.B(n_3127),
.Y(n_4525)
);

O2A1O1Ixp33_ASAP7_75t_L g4526 ( 
.A1(n_3989),
.A2(n_3808),
.B(n_3783),
.C(n_3956),
.Y(n_4526)
);

O2A1O1Ixp33_ASAP7_75t_L g4527 ( 
.A1(n_3989),
.A2(n_3318),
.B(n_3401),
.C(n_3419),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_3834),
.B(n_3092),
.Y(n_4528)
);

AOI21xp5_ASAP7_75t_L g4529 ( 
.A1(n_3886),
.A2(n_3403),
.B(n_3359),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3817),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_3824),
.B(n_3090),
.Y(n_4531)
);

AO21x2_ASAP7_75t_L g4532 ( 
.A1(n_4146),
.A2(n_3430),
.B(n_3419),
.Y(n_4532)
);

AND2x4_ASAP7_75t_L g4533 ( 
.A(n_3767),
.B(n_3393),
.Y(n_4533)
);

OR2x2_ASAP7_75t_L g4534 ( 
.A(n_4075),
.B(n_3079),
.Y(n_4534)
);

AOI22xp33_ASAP7_75t_L g4535 ( 
.A1(n_4077),
.A2(n_4120),
.B1(n_4112),
.B2(n_3740),
.Y(n_4535)
);

BUFx2_ASAP7_75t_L g4536 ( 
.A(n_3996),
.Y(n_4536)
);

AND2x4_ASAP7_75t_L g4537 ( 
.A(n_3767),
.B(n_3393),
.Y(n_4537)
);

OR2x2_ASAP7_75t_L g4538 ( 
.A(n_4075),
.B(n_3079),
.Y(n_4538)
);

NAND3xp33_ASAP7_75t_SL g4539 ( 
.A(n_4082),
.B(n_3944),
.C(n_4013),
.Y(n_4539)
);

AOI21xp5_ASAP7_75t_L g4540 ( 
.A1(n_3886),
.A2(n_3359),
.B(n_3433),
.Y(n_4540)
);

AND2x4_ASAP7_75t_L g4541 ( 
.A(n_3767),
.B(n_3092),
.Y(n_4541)
);

BUFx6f_ASAP7_75t_L g4542 ( 
.A(n_3741),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_3840),
.B(n_3079),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_3817),
.Y(n_4544)
);

OAI21x1_ASAP7_75t_SL g4545 ( 
.A1(n_3680),
.A2(n_3370),
.B(n_3317),
.Y(n_4545)
);

AOI22xp33_ASAP7_75t_L g4546 ( 
.A1(n_4077),
.A2(n_3166),
.B1(n_3051),
.B2(n_3664),
.Y(n_4546)
);

AND2x2_ASAP7_75t_SL g4547 ( 
.A(n_4077),
.B(n_3164),
.Y(n_4547)
);

INVx1_ASAP7_75t_SL g4548 ( 
.A(n_3670),
.Y(n_4548)
);

AOI22xp33_ASAP7_75t_L g4549 ( 
.A1(n_4112),
.A2(n_3042),
.B1(n_3051),
.B2(n_3596),
.Y(n_4549)
);

AOI22xp33_ASAP7_75t_L g4550 ( 
.A1(n_4120),
.A2(n_3042),
.B1(n_3596),
.B2(n_3591),
.Y(n_4550)
);

BUFx6f_ASAP7_75t_L g4551 ( 
.A(n_3773),
.Y(n_4551)
);

A2O1A1Ixp33_ASAP7_75t_L g4552 ( 
.A1(n_3725),
.A2(n_3431),
.B(n_3461),
.C(n_3442),
.Y(n_4552)
);

OAI21x1_ASAP7_75t_L g4553 ( 
.A1(n_3851),
.A2(n_3791),
.B(n_3773),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_3680),
.A2(n_3591),
.B1(n_3507),
.B2(n_3488),
.Y(n_4554)
);

INVx1_ASAP7_75t_SL g4555 ( 
.A(n_3670),
.Y(n_4555)
);

AND2x6_ASAP7_75t_L g4556 ( 
.A(n_3713),
.B(n_3216),
.Y(n_4556)
);

INVx2_ASAP7_75t_SL g4557 ( 
.A(n_4064),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_3671),
.B(n_3164),
.Y(n_4558)
);

BUFx6f_ASAP7_75t_L g4559 ( 
.A(n_3791),
.Y(n_4559)
);

BUFx6f_ASAP7_75t_L g4560 ( 
.A(n_3791),
.Y(n_4560)
);

OAI22xp5_ASAP7_75t_L g4561 ( 
.A1(n_4176),
.A2(n_3243),
.B1(n_3239),
.B2(n_3249),
.Y(n_4561)
);

OAI21x1_ASAP7_75t_L g4562 ( 
.A1(n_4051),
.A2(n_4151),
.B(n_4158),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_3833),
.Y(n_4563)
);

INVx1_ASAP7_75t_SL g4564 ( 
.A(n_3704),
.Y(n_4564)
);

O2A1O1Ixp33_ASAP7_75t_SL g4565 ( 
.A1(n_3737),
.A2(n_3463),
.B(n_3466),
.C(n_3465),
.Y(n_4565)
);

INVx1_ASAP7_75t_SL g4566 ( 
.A(n_3704),
.Y(n_4566)
);

AO21x2_ASAP7_75t_L g4567 ( 
.A1(n_4177),
.A2(n_3352),
.B(n_3355),
.Y(n_4567)
);

OAI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_3840),
.A2(n_3445),
.B(n_3352),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_3671),
.B(n_3164),
.Y(n_4569)
);

HB1xp67_ASAP7_75t_L g4570 ( 
.A(n_3841),
.Y(n_4570)
);

AND2x4_ASAP7_75t_L g4571 ( 
.A(n_4096),
.B(n_3216),
.Y(n_4571)
);

NAND2x1p5_ASAP7_75t_L g4572 ( 
.A(n_3929),
.B(n_3216),
.Y(n_4572)
);

NAND2x1p5_ASAP7_75t_L g4573 ( 
.A(n_3929),
.B(n_3236),
.Y(n_4573)
);

BUFx12f_ASAP7_75t_L g4574 ( 
.A(n_3799),
.Y(n_4574)
);

OAI222xp33_ASAP7_75t_L g4575 ( 
.A1(n_3783),
.A2(n_3071),
.B1(n_3076),
.B2(n_3091),
.C1(n_3126),
.C2(n_3137),
.Y(n_4575)
);

OAI21x1_ASAP7_75t_L g4576 ( 
.A1(n_4051),
.A2(n_4151),
.B(n_4158),
.Y(n_4576)
);

AOI221xp5_ASAP7_75t_L g4577 ( 
.A1(n_3808),
.A2(n_3405),
.B1(n_3076),
.B2(n_3091),
.C(n_3126),
.Y(n_4577)
);

HB1xp67_ASAP7_75t_L g4578 ( 
.A(n_3841),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_3833),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_3839),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_3839),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_3845),
.Y(n_4582)
);

INVx1_ASAP7_75t_SL g4583 ( 
.A(n_3706),
.Y(n_4583)
);

INVx3_ASAP7_75t_SL g4584 ( 
.A(n_4171),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_3845),
.Y(n_4585)
);

AND2x4_ASAP7_75t_L g4586 ( 
.A(n_4096),
.B(n_3236),
.Y(n_4586)
);

BUFx2_ASAP7_75t_L g4587 ( 
.A(n_3996),
.Y(n_4587)
);

INVx2_ASAP7_75t_SL g4588 ( 
.A(n_4064),
.Y(n_4588)
);

BUFx3_ASAP7_75t_L g4589 ( 
.A(n_3799),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_3852),
.Y(n_4590)
);

INVx3_ASAP7_75t_L g4591 ( 
.A(n_3898),
.Y(n_4591)
);

O2A1O1Ixp33_ASAP7_75t_SL g4592 ( 
.A1(n_3737),
.A2(n_3458),
.B(n_3467),
.C(n_3450),
.Y(n_4592)
);

AOI22xp33_ASAP7_75t_L g4593 ( 
.A1(n_3680),
.A2(n_3507),
.B1(n_3488),
.B2(n_3614),
.Y(n_4593)
);

OAI21x1_ASAP7_75t_L g4594 ( 
.A1(n_4151),
.A2(n_4160),
.B(n_4054),
.Y(n_4594)
);

HB1xp67_ASAP7_75t_L g4595 ( 
.A(n_4011),
.Y(n_4595)
);

OR2x6_ASAP7_75t_L g4596 ( 
.A(n_3803),
.B(n_3405),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_3886),
.A2(n_3408),
.B(n_3429),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_3852),
.Y(n_4598)
);

OAI21x1_ASAP7_75t_L g4599 ( 
.A1(n_4160),
.A2(n_3459),
.B(n_3363),
.Y(n_4599)
);

AOI22xp33_ASAP7_75t_L g4600 ( 
.A1(n_3680),
.A2(n_3614),
.B1(n_3137),
.B2(n_3149),
.Y(n_4600)
);

OR2x6_ASAP7_75t_L g4601 ( 
.A(n_3803),
.B(n_3408),
.Y(n_4601)
);

BUFx6f_ASAP7_75t_L g4602 ( 
.A(n_3673),
.Y(n_4602)
);

NAND2x1p5_ASAP7_75t_L g4603 ( 
.A(n_3929),
.B(n_3302),
.Y(n_4603)
);

BUFx3_ASAP7_75t_L g4604 ( 
.A(n_3835),
.Y(n_4604)
);

OAI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_3916),
.A2(n_3347),
.B(n_3353),
.Y(n_4605)
);

BUFx12f_ASAP7_75t_L g4606 ( 
.A(n_3835),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_3855),
.Y(n_4607)
);

AOI222xp33_ASAP7_75t_L g4608 ( 
.A1(n_3956),
.A2(n_3203),
.B1(n_3237),
.B2(n_3071),
.C1(n_3239),
.C2(n_3233),
.Y(n_4608)
);

AOI22xp33_ASAP7_75t_L g4609 ( 
.A1(n_3740),
.A2(n_3149),
.B1(n_3340),
.B2(n_3303),
.Y(n_4609)
);

AOI21xp5_ASAP7_75t_L g4610 ( 
.A1(n_3886),
.A2(n_3364),
.B(n_3358),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_3671),
.B(n_3164),
.Y(n_4611)
);

AOI22xp33_ASAP7_75t_L g4612 ( 
.A1(n_3740),
.A2(n_3753),
.B1(n_3937),
.B2(n_4078),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_3855),
.Y(n_4613)
);

AOI21xp5_ASAP7_75t_L g4614 ( 
.A1(n_3886),
.A2(n_3368),
.B(n_3358),
.Y(n_4614)
);

HB1xp67_ASAP7_75t_L g4615 ( 
.A(n_4039),
.Y(n_4615)
);

AOI21x1_ASAP7_75t_L g4616 ( 
.A1(n_3688),
.A2(n_3467),
.B(n_3458),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_3857),
.Y(n_4617)
);

AO21x2_ASAP7_75t_L g4618 ( 
.A1(n_4180),
.A2(n_4196),
.B(n_3961),
.Y(n_4618)
);

OAI22xp5_ASAP7_75t_L g4619 ( 
.A1(n_3810),
.A2(n_3237),
.B1(n_3350),
.B2(n_3346),
.Y(n_4619)
);

INVx3_ASAP7_75t_L g4620 ( 
.A(n_3898),
.Y(n_4620)
);

AND2x4_ASAP7_75t_L g4621 ( 
.A(n_4096),
.B(n_4119),
.Y(n_4621)
);

AND2x4_ASAP7_75t_L g4622 ( 
.A(n_4096),
.B(n_3395),
.Y(n_4622)
);

OAI22xp5_ASAP7_75t_L g4623 ( 
.A1(n_3810),
.A2(n_3350),
.B1(n_3346),
.B2(n_3233),
.Y(n_4623)
);

HB1xp67_ASAP7_75t_L g4624 ( 
.A(n_4039),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_3857),
.Y(n_4625)
);

O2A1O1Ixp33_ASAP7_75t_L g4626 ( 
.A1(n_3946),
.A2(n_3586),
.B(n_3443),
.C(n_3469),
.Y(n_4626)
);

OAI21x1_ASAP7_75t_SL g4627 ( 
.A1(n_3740),
.A2(n_3443),
.B(n_3374),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_L g4628 ( 
.A(n_3916),
.B(n_3143),
.Y(n_4628)
);

NOR2xp33_ASAP7_75t_L g4629 ( 
.A(n_3937),
.B(n_3340),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_3868),
.Y(n_4630)
);

OAI21x1_ASAP7_75t_SL g4631 ( 
.A1(n_3753),
.A2(n_3374),
.B(n_3440),
.Y(n_4631)
);

BUFx2_ASAP7_75t_L g4632 ( 
.A(n_3996),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_3676),
.B(n_3143),
.Y(n_4633)
);

HB1xp67_ASAP7_75t_L g4634 ( 
.A(n_3688),
.Y(n_4634)
);

OAI21xp5_ASAP7_75t_L g4635 ( 
.A1(n_3950),
.A2(n_3472),
.B(n_3469),
.Y(n_4635)
);

INVx1_ASAP7_75t_SL g4636 ( 
.A(n_3706),
.Y(n_4636)
);

O2A1O1Ixp33_ASAP7_75t_L g4637 ( 
.A1(n_3946),
.A2(n_3472),
.B(n_3456),
.C(n_3451),
.Y(n_4637)
);

OAI21xp5_ASAP7_75t_L g4638 ( 
.A1(n_3950),
.A2(n_3456),
.B(n_3451),
.Y(n_4638)
);

OAI22xp33_ASAP7_75t_L g4639 ( 
.A1(n_4188),
.A2(n_3298),
.B1(n_3345),
.B2(n_3344),
.Y(n_4639)
);

NAND2x1p5_ASAP7_75t_L g4640 ( 
.A(n_3929),
.B(n_3308),
.Y(n_4640)
);

OR2x6_ASAP7_75t_L g4641 ( 
.A(n_3803),
.B(n_3869),
.Y(n_4641)
);

INVx2_ASAP7_75t_SL g4642 ( 
.A(n_4064),
.Y(n_4642)
);

NOR2x1_ASAP7_75t_R g4643 ( 
.A(n_3928),
.B(n_3835),
.Y(n_4643)
);

A2O1A1Ixp33_ASAP7_75t_L g4644 ( 
.A1(n_3735),
.A2(n_3303),
.B(n_3339),
.C(n_3337),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_3959),
.B(n_3143),
.Y(n_4645)
);

INVx1_ASAP7_75t_SL g4646 ( 
.A(n_3714),
.Y(n_4646)
);

NOR2xp33_ASAP7_75t_L g4647 ( 
.A(n_3937),
.B(n_3344),
.Y(n_4647)
);

BUFx6f_ASAP7_75t_L g4648 ( 
.A(n_3673),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_3676),
.B(n_3143),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_3959),
.B(n_3143),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_3868),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_3884),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_3884),
.Y(n_4653)
);

OAI22xp5_ASAP7_75t_SL g4654 ( 
.A1(n_4052),
.A2(n_3450),
.B1(n_3339),
.B2(n_3337),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_3887),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_3887),
.Y(n_4656)
);

CKINVDCx8_ASAP7_75t_R g4657 ( 
.A(n_3735),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_3937),
.B(n_3345),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_3889),
.Y(n_4659)
);

A2O1A1Ixp33_ASAP7_75t_L g4660 ( 
.A1(n_4055),
.A2(n_3302),
.B(n_3308),
.C(n_3258),
.Y(n_4660)
);

NOR2xp33_ASAP7_75t_L g4661 ( 
.A(n_4185),
.B(n_3287),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_3721),
.Y(n_4662)
);

INVx1_ASAP7_75t_SL g4663 ( 
.A(n_3714),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_3889),
.Y(n_4664)
);

BUFx4_ASAP7_75t_SL g4665 ( 
.A(n_3690),
.Y(n_4665)
);

INVx3_ASAP7_75t_L g4666 ( 
.A(n_3898),
.Y(n_4666)
);

OAI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_3981),
.A2(n_3407),
.B(n_3399),
.Y(n_4667)
);

OAI21x1_ASAP7_75t_L g4668 ( 
.A1(n_4130),
.A2(n_3399),
.B(n_3398),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_3893),
.Y(n_4669)
);

NAND3xp33_ASAP7_75t_L g4670 ( 
.A(n_3981),
.B(n_4006),
.C(n_3997),
.Y(n_4670)
);

BUFx3_ASAP7_75t_L g4671 ( 
.A(n_4037),
.Y(n_4671)
);

NAND2xp33_ASAP7_75t_R g4672 ( 
.A(n_3872),
.B(n_3283),
.Y(n_4672)
);

OAI21xp5_ASAP7_75t_L g4673 ( 
.A1(n_3997),
.A2(n_4032),
.B(n_4006),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_3893),
.Y(n_4674)
);

NAND2x1p5_ASAP7_75t_L g4675 ( 
.A(n_3929),
.B(n_4108),
.Y(n_4675)
);

AOI221xp5_ASAP7_75t_L g4676 ( 
.A1(n_3948),
.A2(n_3258),
.B1(n_3298),
.B2(n_3283),
.C(n_3287),
.Y(n_4676)
);

AOI21x1_ASAP7_75t_L g4677 ( 
.A1(n_3894),
.A2(n_3307),
.B(n_3300),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4032),
.B(n_3211),
.Y(n_4678)
);

AOI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4098),
.A2(n_3308),
.B1(n_3302),
.B2(n_3281),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_3894),
.Y(n_4680)
);

A2O1A1Ixp33_ASAP7_75t_L g4681 ( 
.A1(n_4055),
.A2(n_3308),
.B(n_3302),
.C(n_3300),
.Y(n_4681)
);

CKINVDCx5p33_ASAP7_75t_R g4682 ( 
.A(n_3721),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_3907),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_3886),
.A2(n_3299),
.B(n_3280),
.Y(n_4684)
);

OAI21x1_ASAP7_75t_L g4685 ( 
.A1(n_3869),
.A2(n_3877),
.B(n_3709),
.Y(n_4685)
);

AOI211xp5_ASAP7_75t_L g4686 ( 
.A1(n_4078),
.A2(n_3299),
.B(n_3280),
.C(n_3281),
.Y(n_4686)
);

AND2x2_ASAP7_75t_SL g4687 ( 
.A(n_3785),
.B(n_3679),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_3907),
.Y(n_4688)
);

OAI22xp5_ASAP7_75t_L g4689 ( 
.A1(n_3930),
.A2(n_4085),
.B1(n_4174),
.B2(n_3801),
.Y(n_4689)
);

AOI21xp5_ASAP7_75t_L g4690 ( 
.A1(n_4090),
.A2(n_3217),
.B(n_3281),
.Y(n_4690)
);

OR2x2_ASAP7_75t_L g4691 ( 
.A(n_4076),
.B(n_4105),
.Y(n_4691)
);

CKINVDCx5p33_ASAP7_75t_R g4692 ( 
.A(n_3721),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_3908),
.Y(n_4693)
);

OA21x2_ASAP7_75t_L g4694 ( 
.A1(n_3818),
.A2(n_3217),
.B(n_3291),
.Y(n_4694)
);

OAI21x1_ASAP7_75t_L g4695 ( 
.A1(n_3877),
.A2(n_3709),
.B(n_3695),
.Y(n_4695)
);

BUFx2_ASAP7_75t_R g4696 ( 
.A(n_3690),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_3908),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_3915),
.Y(n_4698)
);

INVx3_ASAP7_75t_L g4699 ( 
.A(n_4070),
.Y(n_4699)
);

BUFx10_ASAP7_75t_L g4700 ( 
.A(n_3738),
.Y(n_4700)
);

A2O1A1Ixp33_ASAP7_75t_L g4701 ( 
.A1(n_4062),
.A2(n_3421),
.B(n_3361),
.C(n_3371),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_3915),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_3919),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_3785),
.B(n_3357),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_3919),
.Y(n_4705)
);

XOR2x2_ASAP7_75t_SL g4706 ( 
.A(n_3905),
.B(n_3357),
.Y(n_4706)
);

AOI21x1_ASAP7_75t_L g4707 ( 
.A1(n_3925),
.A2(n_3933),
.B(n_3927),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_3925),
.Y(n_4708)
);

NAND2x1p5_ASAP7_75t_L g4709 ( 
.A(n_3929),
.B(n_3376),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_3927),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_3933),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4042),
.B(n_3376),
.Y(n_4712)
);

BUFx3_ASAP7_75t_L g4713 ( 
.A(n_4037),
.Y(n_4713)
);

INVx2_ASAP7_75t_SL g4714 ( 
.A(n_4064),
.Y(n_4714)
);

INVx4_ASAP7_75t_L g4715 ( 
.A(n_3711),
.Y(n_4715)
);

OAI22xp33_ASAP7_75t_L g4716 ( 
.A1(n_4188),
.A2(n_3402),
.B1(n_3420),
.B2(n_3897),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_L g4717 ( 
.A(n_4157),
.B(n_3420),
.Y(n_4717)
);

AOI22xp33_ASAP7_75t_L g4718 ( 
.A1(n_3882),
.A2(n_3420),
.B1(n_3890),
.B2(n_4141),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4118),
.B(n_4186),
.Y(n_4719)
);

AOI21x1_ASAP7_75t_L g4720 ( 
.A1(n_3940),
.A2(n_3952),
.B(n_3945),
.Y(n_4720)
);

INVx2_ASAP7_75t_SL g4721 ( 
.A(n_4064),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4042),
.B(n_3674),
.Y(n_4722)
);

OR2x2_ASAP7_75t_L g4723 ( 
.A(n_4076),
.B(n_4105),
.Y(n_4723)
);

BUFx2_ASAP7_75t_L g4724 ( 
.A(n_4135),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_3940),
.Y(n_4725)
);

OAI221xp5_ASAP7_75t_L g4726 ( 
.A1(n_4118),
.A2(n_4186),
.B1(n_4132),
.B2(n_4125),
.C(n_4045),
.Y(n_4726)
);

OAI21x1_ASAP7_75t_L g4727 ( 
.A1(n_3710),
.A2(n_3784),
.B(n_3749),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4042),
.B(n_3674),
.Y(n_4728)
);

OAI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_3897),
.A2(n_3906),
.B1(n_4127),
.B2(n_3942),
.Y(n_4729)
);

O2A1O1Ixp33_ASAP7_75t_L g4730 ( 
.A1(n_4125),
.A2(n_4132),
.B(n_4045),
.C(n_3922),
.Y(n_4730)
);

OAI21x1_ASAP7_75t_L g4731 ( 
.A1(n_3749),
.A2(n_3784),
.B(n_4019),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_3945),
.Y(n_4732)
);

AOI21xp5_ASAP7_75t_L g4733 ( 
.A1(n_3929),
.A2(n_3881),
.B(n_3679),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4022),
.B(n_4026),
.Y(n_4734)
);

CKINVDCx20_ASAP7_75t_R g4735 ( 
.A(n_3718),
.Y(n_4735)
);

OAI21x1_ASAP7_75t_L g4736 ( 
.A1(n_3749),
.A2(n_3784),
.B(n_4027),
.Y(n_4736)
);

OR3x4_ASAP7_75t_SL g4737 ( 
.A(n_3707),
.B(n_3928),
.C(n_4127),
.Y(n_4737)
);

AOI21x1_ASAP7_75t_L g4738 ( 
.A1(n_3952),
.A2(n_3969),
.B(n_3968),
.Y(n_4738)
);

NAND2x1p5_ASAP7_75t_L g4739 ( 
.A(n_4108),
.B(n_4115),
.Y(n_4739)
);

OAI21x1_ASAP7_75t_L g4740 ( 
.A1(n_3784),
.A2(n_4027),
.B(n_3798),
.Y(n_4740)
);

INVx2_ASAP7_75t_SL g4741 ( 
.A(n_4073),
.Y(n_4741)
);

OAI21x1_ASAP7_75t_L g4742 ( 
.A1(n_4027),
.A2(n_3798),
.B(n_3789),
.Y(n_4742)
);

OAI21xp5_ASAP7_75t_L g4743 ( 
.A1(n_3764),
.A2(n_4145),
.B(n_4139),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4022),
.B(n_4026),
.Y(n_4744)
);

OA21x2_ASAP7_75t_L g4745 ( 
.A1(n_4035),
.A2(n_4038),
.B(n_3969),
.Y(n_4745)
);

INVx3_ASAP7_75t_L g4746 ( 
.A(n_4070),
.Y(n_4746)
);

OAI21x1_ASAP7_75t_L g4747 ( 
.A1(n_3798),
.A2(n_3806),
.B(n_3804),
.Y(n_4747)
);

OAI21x1_ASAP7_75t_L g4748 ( 
.A1(n_3804),
.A2(n_3807),
.B(n_3806),
.Y(n_4748)
);

AO21x2_ASAP7_75t_L g4749 ( 
.A1(n_3968),
.A2(n_3980),
.B(n_3979),
.Y(n_4749)
);

OAI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_3764),
.A2(n_4145),
.B(n_4139),
.Y(n_4750)
);

NOR2x1_ASAP7_75t_L g4751 ( 
.A(n_3797),
.B(n_3856),
.Y(n_4751)
);

AOI22xp33_ASAP7_75t_L g4752 ( 
.A1(n_3882),
.A2(n_3890),
.B1(n_4124),
.B2(n_3992),
.Y(n_4752)
);

AO31x2_ASAP7_75t_L g4753 ( 
.A1(n_3804),
.A2(n_3807),
.A3(n_3812),
.B(n_3806),
.Y(n_4753)
);

OAI221xp5_ASAP7_75t_L g4754 ( 
.A1(n_3797),
.A2(n_3856),
.B1(n_3922),
.B2(n_3923),
.C(n_3895),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_3807),
.Y(n_4755)
);

OA21x2_ASAP7_75t_L g4756 ( 
.A1(n_4035),
.A2(n_3980),
.B(n_3979),
.Y(n_4756)
);

AND2x4_ASAP7_75t_L g4757 ( 
.A(n_4119),
.B(n_3829),
.Y(n_4757)
);

OR2x6_ASAP7_75t_L g4758 ( 
.A(n_4119),
.B(n_3802),
.Y(n_4758)
);

INVx4_ASAP7_75t_L g4759 ( 
.A(n_4392),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4756),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4345),
.B(n_3726),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4201),
.Y(n_4762)
);

BUFx4_ASAP7_75t_R g4763 ( 
.A(n_4226),
.Y(n_4763)
);

BUFx2_ASAP7_75t_L g4764 ( 
.A(n_4758),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4743),
.B(n_4110),
.Y(n_4765)
);

OAI22xp5_ASAP7_75t_L g4766 ( 
.A1(n_4206),
.A2(n_3930),
.B1(n_4174),
.B2(n_3942),
.Y(n_4766)
);

NAND2x1p5_ASAP7_75t_L g4767 ( 
.A(n_4751),
.B(n_4073),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4201),
.Y(n_4768)
);

INVx2_ASAP7_75t_L g4769 ( 
.A(n_4756),
.Y(n_4769)
);

AOI22xp33_ASAP7_75t_SL g4770 ( 
.A1(n_4221),
.A2(n_3879),
.B1(n_4066),
.B2(n_3801),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4213),
.Y(n_4771)
);

NOR2xp33_ASAP7_75t_L g4772 ( 
.A(n_4409),
.B(n_3882),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4213),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4756),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4488),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4756),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4488),
.Y(n_4777)
);

AND2x2_ASAP7_75t_L g4778 ( 
.A(n_4345),
.B(n_3726),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4756),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4490),
.Y(n_4780)
);

AND2x2_ASAP7_75t_L g4781 ( 
.A(n_4345),
.B(n_3728),
.Y(n_4781)
);

CKINVDCx11_ASAP7_75t_R g4782 ( 
.A(n_4324),
.Y(n_4782)
);

INVx6_ASAP7_75t_L g4783 ( 
.A(n_4364),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4224),
.B(n_3728),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4745),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4490),
.Y(n_4786)
);

AOI22xp33_ASAP7_75t_L g4787 ( 
.A1(n_4207),
.A2(n_3890),
.B1(n_3879),
.B2(n_3801),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4491),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4745),
.Y(n_4789)
);

BUFx3_ASAP7_75t_L g4790 ( 
.A(n_4392),
.Y(n_4790)
);

INVx2_ASAP7_75t_SL g4791 ( 
.A(n_4621),
.Y(n_4791)
);

OR2x6_ASAP7_75t_L g4792 ( 
.A(n_4295),
.B(n_3802),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4745),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4491),
.Y(n_4794)
);

OAI22xp5_ASAP7_75t_L g4795 ( 
.A1(n_4219),
.A2(n_3942),
.B1(n_3906),
.B2(n_4085),
.Y(n_4795)
);

OAI22xp5_ASAP7_75t_L g4796 ( 
.A1(n_4259),
.A2(n_4085),
.B1(n_3954),
.B2(n_3687),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4502),
.Y(n_4797)
);

OA21x2_ASAP7_75t_L g4798 ( 
.A1(n_4361),
.A2(n_3885),
.B(n_3781),
.Y(n_4798)
);

OAI22xp5_ASAP7_75t_L g4799 ( 
.A1(n_4306),
.A2(n_3954),
.B1(n_3687),
.B2(n_4162),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4502),
.Y(n_4800)
);

AOI22xp33_ASAP7_75t_SL g4801 ( 
.A1(n_4221),
.A2(n_4320),
.B1(n_4207),
.B2(n_4203),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4509),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4745),
.Y(n_4803)
);

OAI22xp5_ASAP7_75t_L g4804 ( 
.A1(n_4229),
.A2(n_3954),
.B1(n_3687),
.B2(n_4193),
.Y(n_4804)
);

OAI22xp5_ASAP7_75t_L g4805 ( 
.A1(n_4229),
.A2(n_3687),
.B1(n_4088),
.B2(n_4084),
.Y(n_4805)
);

HB1xp67_ASAP7_75t_L g4806 ( 
.A(n_4394),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4509),
.Y(n_4807)
);

INVx2_ASAP7_75t_SL g4808 ( 
.A(n_4621),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4518),
.Y(n_4809)
);

OAI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4232),
.A2(n_3911),
.B(n_3905),
.Y(n_4810)
);

AOI22xp5_ASAP7_75t_L g4811 ( 
.A1(n_4257),
.A2(n_4127),
.B1(n_3879),
.B2(n_4066),
.Y(n_4811)
);

BUFx12f_ASAP7_75t_L g4812 ( 
.A(n_4392),
.Y(n_4812)
);

AO21x2_ASAP7_75t_L g4813 ( 
.A1(n_4291),
.A2(n_3815),
.B(n_3812),
.Y(n_4813)
);

INVx4_ASAP7_75t_L g4814 ( 
.A(n_4422),
.Y(n_4814)
);

INVx2_ASAP7_75t_L g4815 ( 
.A(n_4745),
.Y(n_4815)
);

AOI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_4257),
.A2(n_3879),
.B1(n_4066),
.B2(n_3801),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4742),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4742),
.Y(n_4818)
);

AOI22xp33_ASAP7_75t_L g4819 ( 
.A1(n_4323),
.A2(n_3879),
.B1(n_4066),
.B2(n_3801),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4742),
.Y(n_4820)
);

OA21x2_ASAP7_75t_L g4821 ( 
.A1(n_4361),
.A2(n_3885),
.B(n_3781),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4518),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4743),
.B(n_4110),
.Y(n_4823)
);

AO21x1_ASAP7_75t_L g4824 ( 
.A1(n_4292),
.A2(n_3900),
.B(n_3844),
.Y(n_4824)
);

BUFx8_ASAP7_75t_SL g4825 ( 
.A(n_4476),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4530),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4694),
.Y(n_4827)
);

NOR2xp33_ASAP7_75t_L g4828 ( 
.A(n_4539),
.B(n_3928),
.Y(n_4828)
);

NOR2xp67_ASAP7_75t_SL g4829 ( 
.A(n_4657),
.B(n_3675),
.Y(n_4829)
);

OAI21x1_ASAP7_75t_L g4830 ( 
.A1(n_4351),
.A2(n_4361),
.B(n_4424),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4530),
.Y(n_4831)
);

AOI22xp5_ASAP7_75t_L g4832 ( 
.A1(n_4262),
.A2(n_4278),
.B1(n_4329),
.B2(n_4323),
.Y(n_4832)
);

BUFx2_ASAP7_75t_L g4833 ( 
.A(n_4758),
.Y(n_4833)
);

AND2x2_ASAP7_75t_L g4834 ( 
.A(n_4224),
.B(n_4687),
.Y(n_4834)
);

INVx3_ASAP7_75t_SL g4835 ( 
.A(n_4415),
.Y(n_4835)
);

BUFx12f_ASAP7_75t_L g4836 ( 
.A(n_4422),
.Y(n_4836)
);

OAI21x1_ASAP7_75t_L g4837 ( 
.A1(n_4351),
.A2(n_3941),
.B(n_3935),
.Y(n_4837)
);

INVx2_ASAP7_75t_L g4838 ( 
.A(n_4694),
.Y(n_4838)
);

INVx2_ASAP7_75t_L g4839 ( 
.A(n_4694),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4544),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4544),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4563),
.Y(n_4842)
);

INVx2_ASAP7_75t_L g4843 ( 
.A(n_4694),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4694),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4563),
.Y(n_4845)
);

HB1xp67_ASAP7_75t_L g4846 ( 
.A(n_4595),
.Y(n_4846)
);

AOI21x1_ASAP7_75t_L g4847 ( 
.A1(n_4291),
.A2(n_3957),
.B(n_3876),
.Y(n_4847)
);

BUFx8_ASAP7_75t_L g4848 ( 
.A(n_4422),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4224),
.B(n_4043),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4687),
.B(n_3921),
.Y(n_4850)
);

OAI22xp5_ASAP7_75t_L g4851 ( 
.A1(n_4335),
.A2(n_4148),
.B1(n_4062),
.B2(n_3879),
.Y(n_4851)
);

INVx4_ASAP7_75t_L g4852 ( 
.A(n_4574),
.Y(n_4852)
);

INVx3_ASAP7_75t_L g4853 ( 
.A(n_4602),
.Y(n_4853)
);

BUFx12f_ASAP7_75t_L g4854 ( 
.A(n_4574),
.Y(n_4854)
);

OAI22xp5_ASAP7_75t_L g4855 ( 
.A1(n_4335),
.A2(n_4148),
.B1(n_4066),
.B2(n_3801),
.Y(n_4855)
);

OAI21x1_ASAP7_75t_L g4856 ( 
.A1(n_4424),
.A2(n_3941),
.B(n_3935),
.Y(n_4856)
);

AND2x4_ASAP7_75t_L g4857 ( 
.A(n_4758),
.B(n_4119),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4579),
.Y(n_4858)
);

OAI22xp5_ASAP7_75t_L g4859 ( 
.A1(n_4319),
.A2(n_4148),
.B1(n_4066),
.B2(n_3900),
.Y(n_4859)
);

OAI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_4383),
.A2(n_3844),
.B1(n_3711),
.B2(n_3730),
.Y(n_4860)
);

BUFx3_ASAP7_75t_L g4861 ( 
.A(n_4574),
.Y(n_4861)
);

BUFx4_ASAP7_75t_SL g4862 ( 
.A(n_4735),
.Y(n_4862)
);

AOI22xp33_ASAP7_75t_L g4863 ( 
.A1(n_4203),
.A2(n_4234),
.B1(n_4320),
.B2(n_4329),
.Y(n_4863)
);

CKINVDCx20_ASAP7_75t_R g4864 ( 
.A(n_4469),
.Y(n_4864)
);

AOI22xp33_ASAP7_75t_L g4865 ( 
.A1(n_4234),
.A2(n_4278),
.B1(n_4262),
.B2(n_4211),
.Y(n_4865)
);

BUFx12f_ASAP7_75t_L g4866 ( 
.A(n_4606),
.Y(n_4866)
);

BUFx12f_ASAP7_75t_L g4867 ( 
.A(n_4606),
.Y(n_4867)
);

AOI22xp33_ASAP7_75t_L g4868 ( 
.A1(n_4211),
.A2(n_3974),
.B1(n_3975),
.B2(n_3896),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4750),
.B(n_4114),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4579),
.Y(n_4870)
);

BUFx8_ASAP7_75t_L g4871 ( 
.A(n_4606),
.Y(n_4871)
);

BUFx8_ASAP7_75t_L g4872 ( 
.A(n_4399),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4580),
.Y(n_4873)
);

HB1xp67_ASAP7_75t_L g4874 ( 
.A(n_4615),
.Y(n_4874)
);

INVx3_ASAP7_75t_L g4875 ( 
.A(n_4602),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4580),
.Y(n_4876)
);

HB1xp67_ASAP7_75t_L g4877 ( 
.A(n_4624),
.Y(n_4877)
);

OAI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4383),
.A2(n_3711),
.B1(n_3730),
.B2(n_3992),
.Y(n_4878)
);

BUFx10_ASAP7_75t_L g4879 ( 
.A(n_4662),
.Y(n_4879)
);

AOI21x1_ASAP7_75t_L g4880 ( 
.A1(n_4204),
.A2(n_3957),
.B(n_3876),
.Y(n_4880)
);

NAND2x1p5_ASAP7_75t_L g4881 ( 
.A(n_4751),
.B(n_4073),
.Y(n_4881)
);

OAI21x1_ASAP7_75t_L g4882 ( 
.A1(n_4336),
.A2(n_4353),
.B(n_4349),
.Y(n_4882)
);

OAI22xp5_ASAP7_75t_L g4883 ( 
.A1(n_4347),
.A2(n_3711),
.B1(n_3730),
.B2(n_3905),
.Y(n_4883)
);

BUFx12f_ASAP7_75t_L g4884 ( 
.A(n_4682),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4581),
.Y(n_4885)
);

NAND2x1p5_ASAP7_75t_L g4886 ( 
.A(n_4223),
.B(n_4073),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4581),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_4753),
.Y(n_4888)
);

CKINVDCx20_ASAP7_75t_R g4889 ( 
.A(n_4233),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4582),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_4582),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4585),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4585),
.Y(n_4893)
);

AOI22xp33_ASAP7_75t_L g4894 ( 
.A1(n_4239),
.A2(n_3975),
.B1(n_3974),
.B2(n_3896),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4590),
.Y(n_4895)
);

BUFx3_ASAP7_75t_L g4896 ( 
.A(n_4341),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4750),
.B(n_4114),
.Y(n_4897)
);

INVx3_ASAP7_75t_L g4898 ( 
.A(n_4602),
.Y(n_4898)
);

BUFx6f_ASAP7_75t_L g4899 ( 
.A(n_4473),
.Y(n_4899)
);

INVx4_ASAP7_75t_L g4900 ( 
.A(n_4341),
.Y(n_4900)
);

CKINVDCx6p67_ASAP7_75t_R g4901 ( 
.A(n_4415),
.Y(n_4901)
);

AOI22xp33_ASAP7_75t_SL g4902 ( 
.A1(n_4296),
.A2(n_4107),
.B1(n_3713),
.B2(n_4124),
.Y(n_4902)
);

OAI21x1_ASAP7_75t_L g4903 ( 
.A1(n_4336),
.A2(n_3973),
.B(n_3949),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4407),
.B(n_3860),
.Y(n_4904)
);

OR2x6_ASAP7_75t_L g4905 ( 
.A(n_4295),
.B(n_4529),
.Y(n_4905)
);

CKINVDCx6p67_ASAP7_75t_R g4906 ( 
.A(n_4415),
.Y(n_4906)
);

HB1xp67_ASAP7_75t_L g4907 ( 
.A(n_4634),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4407),
.B(n_3860),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_4590),
.Y(n_4909)
);

INVx3_ASAP7_75t_L g4910 ( 
.A(n_4602),
.Y(n_4910)
);

BUFx8_ASAP7_75t_L g4911 ( 
.A(n_4399),
.Y(n_4911)
);

OAI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4239),
.A2(n_3911),
.B(n_3905),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4598),
.Y(n_4913)
);

HB1xp67_ASAP7_75t_L g4914 ( 
.A(n_4634),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4753),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4598),
.Y(n_4916)
);

OAI22xp33_ASAP7_75t_L g4917 ( 
.A1(n_4347),
.A2(n_3770),
.B1(n_3787),
.B2(n_3756),
.Y(n_4917)
);

BUFx6f_ASAP7_75t_SL g4918 ( 
.A(n_4399),
.Y(n_4918)
);

NAND2x1p5_ASAP7_75t_L g4919 ( 
.A(n_4223),
.B(n_4073),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4607),
.Y(n_4920)
);

BUFx2_ASAP7_75t_L g4921 ( 
.A(n_4758),
.Y(n_4921)
);

CKINVDCx11_ASAP7_75t_R g4922 ( 
.A(n_4737),
.Y(n_4922)
);

OAI22xp5_ASAP7_75t_L g4923 ( 
.A1(n_4296),
.A2(n_3730),
.B1(n_3970),
.B2(n_3911),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4607),
.Y(n_4924)
);

CKINVDCx11_ASAP7_75t_R g4925 ( 
.A(n_4341),
.Y(n_4925)
);

INVx2_ASAP7_75t_L g4926 ( 
.A(n_4753),
.Y(n_4926)
);

CKINVDCx11_ASAP7_75t_R g4927 ( 
.A(n_4341),
.Y(n_4927)
);

HB1xp67_ASAP7_75t_L g4928 ( 
.A(n_4712),
.Y(n_4928)
);

INVxp67_ASAP7_75t_L g4929 ( 
.A(n_4717),
.Y(n_4929)
);

AOI22xp33_ASAP7_75t_L g4930 ( 
.A1(n_4332),
.A2(n_3975),
.B1(n_3974),
.B2(n_3896),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4408),
.B(n_3895),
.Y(n_4931)
);

HB1xp67_ASAP7_75t_L g4932 ( 
.A(n_4712),
.Y(n_4932)
);

AOI22xp33_ASAP7_75t_L g4933 ( 
.A1(n_4332),
.A2(n_3975),
.B1(n_3974),
.B2(n_3896),
.Y(n_4933)
);

OAI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4281),
.A2(n_3730),
.B1(n_3970),
.B2(n_3911),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4408),
.B(n_3923),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4613),
.Y(n_4936)
);

NAND2x1p5_ASAP7_75t_L g4937 ( 
.A(n_4223),
.B(n_4073),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4613),
.Y(n_4938)
);

BUFx8_ASAP7_75t_L g4939 ( 
.A(n_4471),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4617),
.Y(n_4940)
);

NAND2x1p5_ASAP7_75t_L g4941 ( 
.A(n_4223),
.B(n_4073),
.Y(n_4941)
);

BUFx6f_ASAP7_75t_SL g4942 ( 
.A(n_4471),
.Y(n_4942)
);

NAND2x1p5_ASAP7_75t_L g4943 ( 
.A(n_4223),
.B(n_4108),
.Y(n_4943)
);

OAI22xp33_ASAP7_75t_L g4944 ( 
.A1(n_4437),
.A2(n_3770),
.B1(n_3787),
.B2(n_3756),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4617),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4753),
.Y(n_4946)
);

AOI22xp5_ASAP7_75t_L g4947 ( 
.A1(n_4215),
.A2(n_3675),
.B1(n_3838),
.B2(n_3831),
.Y(n_4947)
);

BUFx12f_ASAP7_75t_L g4948 ( 
.A(n_4692),
.Y(n_4948)
);

INVx2_ASAP7_75t_SL g4949 ( 
.A(n_4621),
.Y(n_4949)
);

INVx2_ASAP7_75t_SL g4950 ( 
.A(n_4621),
.Y(n_4950)
);

BUFx2_ASAP7_75t_SL g4951 ( 
.A(n_4657),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4436),
.B(n_3943),
.Y(n_4952)
);

AOI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_4242),
.A2(n_3831),
.B1(n_3847),
.B2(n_3838),
.Y(n_4953)
);

AO21x1_ASAP7_75t_L g4954 ( 
.A1(n_4448),
.A2(n_4094),
.B(n_4097),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4625),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4753),
.Y(n_4956)
);

INVx2_ASAP7_75t_L g4957 ( 
.A(n_4753),
.Y(n_4957)
);

CKINVDCx5p33_ASAP7_75t_R g4958 ( 
.A(n_4420),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4753),
.Y(n_4959)
);

INVx6_ASAP7_75t_SL g4960 ( 
.A(n_4758),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4625),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4747),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4747),
.Y(n_4963)
);

BUFx2_ASAP7_75t_L g4964 ( 
.A(n_4758),
.Y(n_4964)
);

INVx2_ASAP7_75t_SL g4965 ( 
.A(n_4757),
.Y(n_4965)
);

NOR2x1_ASAP7_75t_SL g4966 ( 
.A(n_4475),
.B(n_3871),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4630),
.Y(n_4967)
);

AOI22xp33_ASAP7_75t_L g4968 ( 
.A1(n_4359),
.A2(n_3975),
.B1(n_3974),
.B2(n_3896),
.Y(n_4968)
);

AOI22xp33_ASAP7_75t_L g4969 ( 
.A1(n_4359),
.A2(n_3974),
.B1(n_3975),
.B2(n_3713),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4687),
.B(n_4227),
.Y(n_4970)
);

INVx1_ASAP7_75t_SL g4971 ( 
.A(n_4691),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4630),
.Y(n_4972)
);

OAI21x1_ASAP7_75t_L g4973 ( 
.A1(n_4336),
.A2(n_3973),
.B(n_3949),
.Y(n_4973)
);

OAI21x1_ASAP7_75t_L g4974 ( 
.A1(n_4349),
.A2(n_3973),
.B(n_3949),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4747),
.Y(n_4975)
);

BUFx3_ASAP7_75t_L g4976 ( 
.A(n_4341),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4436),
.B(n_3943),
.Y(n_4977)
);

BUFx4f_ASAP7_75t_L g4978 ( 
.A(n_4341),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4651),
.Y(n_4979)
);

OAI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4204),
.A2(n_3994),
.B(n_3970),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4748),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4651),
.Y(n_4982)
);

BUFx8_ASAP7_75t_L g4983 ( 
.A(n_4471),
.Y(n_4983)
);

INVx2_ASAP7_75t_L g4984 ( 
.A(n_4748),
.Y(n_4984)
);

INVx3_ASAP7_75t_SL g4985 ( 
.A(n_4435),
.Y(n_4985)
);

BUFx2_ASAP7_75t_R g4986 ( 
.A(n_4287),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4652),
.Y(n_4987)
);

INVx2_ASAP7_75t_L g4988 ( 
.A(n_4748),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4652),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_4707),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4707),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4444),
.B(n_3951),
.Y(n_4992)
);

OAI22xp5_ASAP7_75t_L g4993 ( 
.A1(n_4346),
.A2(n_4437),
.B1(n_4202),
.B2(n_4432),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4653),
.Y(n_4994)
);

INVx3_ASAP7_75t_L g4995 ( 
.A(n_4602),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4653),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4227),
.B(n_3921),
.Y(n_4997)
);

HB1xp67_ASAP7_75t_L g4998 ( 
.A(n_4712),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4655),
.Y(n_4999)
);

NOR2xp33_ASAP7_75t_L g5000 ( 
.A(n_4539),
.B(n_4450),
.Y(n_5000)
);

INVx3_ASAP7_75t_L g5001 ( 
.A(n_4602),
.Y(n_5001)
);

HB1xp67_ASAP7_75t_L g5002 ( 
.A(n_4691),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4227),
.B(n_3921),
.Y(n_5003)
);

BUFx3_ASAP7_75t_L g5004 ( 
.A(n_4430),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4444),
.B(n_3951),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4655),
.Y(n_5006)
);

AOI21x1_ASAP7_75t_L g5007 ( 
.A1(n_4616),
.A2(n_3815),
.B(n_3812),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4656),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4656),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4659),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4720),
.Y(n_5011)
);

OAI22x1_ASAP7_75t_SL g5012 ( 
.A1(n_4199),
.A2(n_3707),
.B1(n_3811),
.B2(n_3718),
.Y(n_5012)
);

BUFx2_ASAP7_75t_SL g5013 ( 
.A(n_4657),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4659),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4664),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4664),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4669),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4669),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4279),
.B(n_3772),
.Y(n_5019)
);

INVx2_ASAP7_75t_SL g5020 ( 
.A(n_4757),
.Y(n_5020)
);

INVx3_ASAP7_75t_L g5021 ( 
.A(n_4602),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4674),
.Y(n_5022)
);

INVx5_ASAP7_75t_L g5023 ( 
.A(n_4556),
.Y(n_5023)
);

AOI22xp33_ASAP7_75t_L g5024 ( 
.A1(n_4547),
.A2(n_3974),
.B1(n_3975),
.B2(n_3713),
.Y(n_5024)
);

BUFx2_ASAP7_75t_L g5025 ( 
.A(n_4498),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4674),
.Y(n_5026)
);

BUFx10_ASAP7_75t_L g5027 ( 
.A(n_4217),
.Y(n_5027)
);

BUFx2_ASAP7_75t_SL g5028 ( 
.A(n_4283),
.Y(n_5028)
);

INVx2_ASAP7_75t_L g5029 ( 
.A(n_4720),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4279),
.B(n_3772),
.Y(n_5030)
);

INVx1_ASAP7_75t_SL g5031 ( 
.A(n_4723),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4738),
.Y(n_5032)
);

CKINVDCx6p67_ASAP7_75t_R g5033 ( 
.A(n_4481),
.Y(n_5033)
);

OAI22xp33_ASAP7_75t_L g5034 ( 
.A1(n_4432),
.A2(n_3770),
.B1(n_3787),
.B2(n_3756),
.Y(n_5034)
);

AND2x2_ASAP7_75t_L g5035 ( 
.A(n_4722),
.B(n_3921),
.Y(n_5035)
);

BUFx6f_ASAP7_75t_L g5036 ( 
.A(n_4473),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_4722),
.B(n_3921),
.Y(n_5037)
);

AOI22xp33_ASAP7_75t_L g5038 ( 
.A1(n_4547),
.A2(n_3713),
.B1(n_3720),
.B2(n_4107),
.Y(n_5038)
);

INVx2_ASAP7_75t_L g5039 ( 
.A(n_4738),
.Y(n_5039)
);

INVx2_ASAP7_75t_L g5040 ( 
.A(n_4749),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_4749),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4680),
.Y(n_5042)
);

BUFx3_ASAP7_75t_L g5043 ( 
.A(n_4430),
.Y(n_5043)
);

AOI21x1_ASAP7_75t_L g5044 ( 
.A1(n_4616),
.A2(n_3825),
.B(n_3805),
.Y(n_5044)
);

CKINVDCx8_ASAP7_75t_R g5045 ( 
.A(n_4287),
.Y(n_5045)
);

BUFx3_ASAP7_75t_L g5046 ( 
.A(n_4430),
.Y(n_5046)
);

AO21x1_ASAP7_75t_L g5047 ( 
.A1(n_4448),
.A2(n_4094),
.B(n_4097),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4680),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4683),
.Y(n_5049)
);

AOI22xp5_ASAP7_75t_L g5050 ( 
.A1(n_4276),
.A2(n_3847),
.B1(n_3828),
.B2(n_4124),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_4749),
.Y(n_5051)
);

AO21x1_ASAP7_75t_SL g5052 ( 
.A1(n_4504),
.A2(n_3867),
.B(n_3865),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4683),
.Y(n_5053)
);

OAI22xp5_ASAP7_75t_L g5054 ( 
.A1(n_4346),
.A2(n_3970),
.B1(n_3994),
.B2(n_3828),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4749),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4526),
.B(n_3796),
.Y(n_5056)
);

BUFx4f_ASAP7_75t_L g5057 ( 
.A(n_4430),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_4198),
.Y(n_5058)
);

BUFx3_ASAP7_75t_L g5059 ( 
.A(n_4430),
.Y(n_5059)
);

OR2x2_ASAP7_75t_L g5060 ( 
.A(n_4723),
.B(n_4018),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4688),
.Y(n_5061)
);

INVx6_ASAP7_75t_L g5062 ( 
.A(n_4364),
.Y(n_5062)
);

AOI22xp33_ASAP7_75t_L g5063 ( 
.A1(n_4547),
.A2(n_3713),
.B1(n_3720),
.B2(n_4107),
.Y(n_5063)
);

AND2x2_ASAP7_75t_SL g5064 ( 
.A(n_4398),
.B(n_3679),
.Y(n_5064)
);

BUFx3_ASAP7_75t_L g5065 ( 
.A(n_4430),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4198),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4688),
.Y(n_5067)
);

OAI21x1_ASAP7_75t_L g5068 ( 
.A1(n_4349),
.A2(n_3973),
.B(n_3949),
.Y(n_5068)
);

INVx3_ASAP7_75t_L g5069 ( 
.A(n_4648),
.Y(n_5069)
);

INVxp67_ASAP7_75t_L g5070 ( 
.A(n_4290),
.Y(n_5070)
);

CKINVDCx20_ASAP7_75t_R g5071 ( 
.A(n_4516),
.Y(n_5071)
);

OAI22xp33_ASAP7_75t_L g5072 ( 
.A1(n_4672),
.A2(n_3770),
.B1(n_3787),
.B2(n_3756),
.Y(n_5072)
);

BUFx3_ASAP7_75t_L g5073 ( 
.A(n_4481),
.Y(n_5073)
);

INVx3_ASAP7_75t_L g5074 ( 
.A(n_4648),
.Y(n_5074)
);

BUFx2_ASAP7_75t_L g5075 ( 
.A(n_4498),
.Y(n_5075)
);

AOI22xp33_ASAP7_75t_L g5076 ( 
.A1(n_4348),
.A2(n_3720),
.B1(n_4107),
.B2(n_3822),
.Y(n_5076)
);

INVxp67_ASAP7_75t_L g5077 ( 
.A(n_4647),
.Y(n_5077)
);

HB1xp67_ASAP7_75t_L g5078 ( 
.A(n_4271),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4526),
.B(n_3796),
.Y(n_5079)
);

CKINVDCx8_ASAP7_75t_R g5080 ( 
.A(n_4199),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4451),
.B(n_4031),
.Y(n_5081)
);

BUFx3_ASAP7_75t_L g5082 ( 
.A(n_4481),
.Y(n_5082)
);

INVx2_ASAP7_75t_SL g5083 ( 
.A(n_4757),
.Y(n_5083)
);

OAI21xp5_ASAP7_75t_L g5084 ( 
.A1(n_4244),
.A2(n_3994),
.B(n_3881),
.Y(n_5084)
);

INVx1_ASAP7_75t_SL g5085 ( 
.A(n_4271),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4693),
.Y(n_5086)
);

OAI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4210),
.A2(n_3994),
.B1(n_3828),
.B2(n_3880),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4693),
.Y(n_5088)
);

AOI22xp33_ASAP7_75t_L g5089 ( 
.A1(n_4348),
.A2(n_3720),
.B1(n_4107),
.B2(n_3822),
.Y(n_5089)
);

AOI22xp33_ASAP7_75t_L g5090 ( 
.A1(n_4375),
.A2(n_3822),
.B1(n_3830),
.B2(n_3809),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4697),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4697),
.Y(n_5092)
);

AOI21x1_ASAP7_75t_L g5093 ( 
.A1(n_4439),
.A2(n_3825),
.B(n_3805),
.Y(n_5093)
);

INVxp67_ASAP7_75t_SL g5094 ( 
.A(n_4706),
.Y(n_5094)
);

BUFx6f_ASAP7_75t_L g5095 ( 
.A(n_4473),
.Y(n_5095)
);

CKINVDCx11_ASAP7_75t_R g5096 ( 
.A(n_4521),
.Y(n_5096)
);

OAI22xp33_ASAP7_75t_L g5097 ( 
.A1(n_4460),
.A2(n_3822),
.B1(n_3830),
.B2(n_3809),
.Y(n_5097)
);

INVx3_ASAP7_75t_L g5098 ( 
.A(n_4648),
.Y(n_5098)
);

BUFx2_ASAP7_75t_L g5099 ( 
.A(n_4519),
.Y(n_5099)
);

NAND2x1p5_ASAP7_75t_L g5100 ( 
.A(n_4223),
.B(n_4108),
.Y(n_5100)
);

BUFx10_ASAP7_75t_L g5101 ( 
.A(n_4248),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4698),
.Y(n_5102)
);

INVx2_ASAP7_75t_L g5103 ( 
.A(n_4198),
.Y(n_5103)
);

INVx2_ASAP7_75t_L g5104 ( 
.A(n_4212),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4698),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4702),
.Y(n_5106)
);

INVx2_ASAP7_75t_L g5107 ( 
.A(n_4212),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4702),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_4212),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4703),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_4703),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_4722),
.B(n_3982),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4705),
.Y(n_5113)
);

BUFx12f_ASAP7_75t_L g5114 ( 
.A(n_4521),
.Y(n_5114)
);

CKINVDCx14_ASAP7_75t_R g5115 ( 
.A(n_4282),
.Y(n_5115)
);

INVx2_ASAP7_75t_L g5116 ( 
.A(n_4214),
.Y(n_5116)
);

AO21x1_ASAP7_75t_L g5117 ( 
.A1(n_4457),
.A2(n_4007),
.B(n_4003),
.Y(n_5117)
);

OAI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_4286),
.A2(n_3881),
.B(n_3955),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4705),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_4708),
.Y(n_5120)
);

INVx2_ASAP7_75t_L g5121 ( 
.A(n_4214),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4708),
.Y(n_5122)
);

INVx2_ASAP7_75t_L g5123 ( 
.A(n_4214),
.Y(n_5123)
);

CKINVDCx20_ASAP7_75t_R g5124 ( 
.A(n_4521),
.Y(n_5124)
);

BUFx4f_ASAP7_75t_SL g5125 ( 
.A(n_4589),
.Y(n_5125)
);

HB1xp67_ASAP7_75t_L g5126 ( 
.A(n_4277),
.Y(n_5126)
);

AOI22xp33_ASAP7_75t_SL g5127 ( 
.A1(n_4457),
.A2(n_4124),
.B1(n_3880),
.B2(n_3899),
.Y(n_5127)
);

CKINVDCx6p67_ASAP7_75t_R g5128 ( 
.A(n_4589),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4710),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_4710),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_4711),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4711),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4725),
.Y(n_5133)
);

BUFx2_ASAP7_75t_L g5134 ( 
.A(n_4519),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4725),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4732),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_4732),
.Y(n_5137)
);

OAI21x1_ASAP7_75t_L g5138 ( 
.A1(n_4302),
.A2(n_3977),
.B(n_3983),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4218),
.Y(n_5139)
);

BUFx2_ASAP7_75t_R g5140 ( 
.A(n_4226),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4218),
.Y(n_5141)
);

INVx1_ASAP7_75t_SL g5142 ( 
.A(n_4277),
.Y(n_5142)
);

INVx2_ASAP7_75t_L g5143 ( 
.A(n_4249),
.Y(n_5143)
);

INVxp33_ASAP7_75t_L g5144 ( 
.A(n_4643),
.Y(n_5144)
);

AO21x1_ASAP7_75t_SL g5145 ( 
.A1(n_4479),
.A2(n_3867),
.B(n_3865),
.Y(n_5145)
);

INVx2_ASAP7_75t_L g5146 ( 
.A(n_4249),
.Y(n_5146)
);

INVx2_ASAP7_75t_L g5147 ( 
.A(n_4249),
.Y(n_5147)
);

BUFx6f_ASAP7_75t_L g5148 ( 
.A(n_4473),
.Y(n_5148)
);

NAND2x1p5_ASAP7_75t_L g5149 ( 
.A(n_4223),
.B(n_4108),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4235),
.Y(n_5150)
);

NAND2x1p5_ASAP7_75t_L g5151 ( 
.A(n_4402),
.B(n_4108),
.Y(n_5151)
);

AND2x4_ASAP7_75t_L g5152 ( 
.A(n_4364),
.B(n_4083),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4235),
.Y(n_5153)
);

AOI22xp33_ASAP7_75t_L g5154 ( 
.A1(n_4375),
.A2(n_3830),
.B1(n_3910),
.B2(n_3809),
.Y(n_5154)
);

AO21x1_ASAP7_75t_SL g5155 ( 
.A1(n_4479),
.A2(n_4131),
.B(n_4128),
.Y(n_5155)
);

AND2x2_ASAP7_75t_L g5156 ( 
.A(n_4728),
.B(n_3982),
.Y(n_5156)
);

BUFx2_ASAP7_75t_L g5157 ( 
.A(n_4536),
.Y(n_5157)
);

OAI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4244),
.A2(n_3679),
.B(n_3955),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4236),
.Y(n_5159)
);

OAI21xp5_ASAP7_75t_L g5160 ( 
.A1(n_4398),
.A2(n_4360),
.B(n_4381),
.Y(n_5160)
);

OAI21x1_ASAP7_75t_L g5161 ( 
.A1(n_4302),
.A2(n_3977),
.B(n_3983),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_4254),
.Y(n_5162)
);

INVx2_ASAP7_75t_L g5163 ( 
.A(n_4254),
.Y(n_5163)
);

AOI22xp33_ASAP7_75t_SL g5164 ( 
.A1(n_4209),
.A2(n_3899),
.B1(n_3917),
.B2(n_3871),
.Y(n_5164)
);

AND2x2_ASAP7_75t_L g5165 ( 
.A(n_4728),
.B(n_3982),
.Y(n_5165)
);

AOI21x1_ASAP7_75t_L g5166 ( 
.A1(n_4439),
.A2(n_3827),
.B(n_3805),
.Y(n_5166)
);

OAI21x1_ASAP7_75t_L g5167 ( 
.A1(n_4302),
.A2(n_3993),
.B(n_3983),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_4254),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4236),
.Y(n_5169)
);

AOI22xp33_ASAP7_75t_L g5170 ( 
.A1(n_4385),
.A2(n_3830),
.B1(n_3910),
.B2(n_3809),
.Y(n_5170)
);

AOI22xp33_ASAP7_75t_L g5171 ( 
.A1(n_4385),
.A2(n_3918),
.B1(n_3931),
.B2(n_3910),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_4728),
.B(n_3982),
.Y(n_5172)
);

INVx2_ASAP7_75t_L g5173 ( 
.A(n_4258),
.Y(n_5173)
);

AND2x2_ASAP7_75t_L g5174 ( 
.A(n_4704),
.B(n_4228),
.Y(n_5174)
);

INVx3_ASAP7_75t_L g5175 ( 
.A(n_4648),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4238),
.Y(n_5176)
);

OAI21x1_ASAP7_75t_L g5177 ( 
.A1(n_4309),
.A2(n_4014),
.B(n_3993),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_4238),
.Y(n_5178)
);

BUFx8_ASAP7_75t_SL g5179 ( 
.A(n_4589),
.Y(n_5179)
);

CKINVDCx11_ASAP7_75t_R g5180 ( 
.A(n_4604),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_4253),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_4253),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4255),
.Y(n_5183)
);

OAI22xp5_ASAP7_75t_L g5184 ( 
.A1(n_4505),
.A2(n_3960),
.B1(n_3963),
.B2(n_3917),
.Y(n_5184)
);

BUFx2_ASAP7_75t_L g5185 ( 
.A(n_4536),
.Y(n_5185)
);

BUFx2_ASAP7_75t_L g5186 ( 
.A(n_4587),
.Y(n_5186)
);

INVx2_ASAP7_75t_SL g5187 ( 
.A(n_4757),
.Y(n_5187)
);

BUFx4f_ASAP7_75t_SL g5188 ( 
.A(n_4604),
.Y(n_5188)
);

NOR2x1_ASAP7_75t_R g5189 ( 
.A(n_4604),
.B(n_3724),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4255),
.Y(n_5190)
);

BUFx6f_ASAP7_75t_L g5191 ( 
.A(n_4700),
.Y(n_5191)
);

OAI22xp5_ASAP7_75t_SL g5192 ( 
.A1(n_4754),
.A2(n_4689),
.B1(n_4362),
.B2(n_4417),
.Y(n_5192)
);

CKINVDCx20_ASAP7_75t_R g5193 ( 
.A(n_4226),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4260),
.Y(n_5194)
);

BUFx3_ASAP7_75t_L g5195 ( 
.A(n_4435),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4260),
.Y(n_5196)
);

NOR2xp67_ASAP7_75t_SL g5197 ( 
.A(n_4307),
.B(n_3690),
.Y(n_5197)
);

OAI22xp5_ASAP7_75t_L g5198 ( 
.A1(n_4462),
.A2(n_3963),
.B1(n_3971),
.B2(n_3960),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_4284),
.Y(n_5199)
);

OAI22xp5_ASAP7_75t_L g5200 ( 
.A1(n_4496),
.A2(n_4024),
.B1(n_4030),
.B2(n_3971),
.Y(n_5200)
);

OAI21xp5_ASAP7_75t_L g5201 ( 
.A1(n_4360),
.A2(n_3679),
.B(n_3976),
.Y(n_5201)
);

INVx3_ASAP7_75t_L g5202 ( 
.A(n_4648),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4284),
.Y(n_5203)
);

AOI22xp33_ASAP7_75t_L g5204 ( 
.A1(n_4285),
.A2(n_3918),
.B1(n_3931),
.B2(n_3910),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_4300),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4300),
.Y(n_5206)
);

AOI22xp33_ASAP7_75t_L g5207 ( 
.A1(n_4285),
.A2(n_3931),
.B1(n_3947),
.B2(n_3918),
.Y(n_5207)
);

BUFx3_ASAP7_75t_L g5208 ( 
.A(n_4435),
.Y(n_5208)
);

OAI22xp5_ASAP7_75t_L g5209 ( 
.A1(n_4443),
.A2(n_4030),
.B1(n_4024),
.B2(n_3780),
.Y(n_5209)
);

INVx3_ASAP7_75t_L g5210 ( 
.A(n_4648),
.Y(n_5210)
);

HB1xp67_ASAP7_75t_L g5211 ( 
.A(n_4343),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_4258),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_4314),
.Y(n_5213)
);

HB1xp67_ASAP7_75t_L g5214 ( 
.A(n_4343),
.Y(n_5214)
);

AOI22xp33_ASAP7_75t_L g5215 ( 
.A1(n_4286),
.A2(n_4419),
.B1(n_4352),
.B2(n_4403),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_4258),
.Y(n_5216)
);

OR2x2_ASAP7_75t_L g5217 ( 
.A(n_4451),
.B(n_4018),
.Y(n_5217)
);

BUFx2_ASAP7_75t_R g5218 ( 
.A(n_4307),
.Y(n_5218)
);

BUFx2_ASAP7_75t_SL g5219 ( 
.A(n_4283),
.Y(n_5219)
);

HB1xp67_ASAP7_75t_L g5220 ( 
.A(n_4378),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_4314),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4318),
.Y(n_5222)
);

AOI22xp5_ASAP7_75t_L g5223 ( 
.A1(n_4428),
.A2(n_3931),
.B1(n_3947),
.B2(n_3918),
.Y(n_5223)
);

AOI21xp5_ASAP7_75t_L g5224 ( 
.A1(n_4405),
.A2(n_3901),
.B(n_3802),
.Y(n_5224)
);

BUFx2_ASAP7_75t_L g5225 ( 
.A(n_4587),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4318),
.Y(n_5226)
);

HB1xp67_ASAP7_75t_L g5227 ( 
.A(n_4378),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_4241),
.B(n_4256),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_4325),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4325),
.Y(n_5230)
);

OAI22xp5_ASAP7_75t_L g5231 ( 
.A1(n_4696),
.A2(n_4477),
.B1(n_4535),
.B2(n_4381),
.Y(n_5231)
);

AO21x2_ASAP7_75t_L g5232 ( 
.A1(n_4545),
.A2(n_4189),
.B(n_4007),
.Y(n_5232)
);

BUFx3_ASAP7_75t_L g5233 ( 
.A(n_4584),
.Y(n_5233)
);

BUFx2_ASAP7_75t_L g5234 ( 
.A(n_4632),
.Y(n_5234)
);

INVx4_ASAP7_75t_SL g5235 ( 
.A(n_4584),
.Y(n_5235)
);

INVx5_ASAP7_75t_L g5236 ( 
.A(n_4556),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_4263),
.Y(n_5237)
);

OAI21x1_ASAP7_75t_L g5238 ( 
.A1(n_4309),
.A2(n_4014),
.B(n_3993),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_4263),
.Y(n_5239)
);

OAI21x1_ASAP7_75t_L g5240 ( 
.A1(n_4309),
.A2(n_4014),
.B(n_3993),
.Y(n_5240)
);

AND2x2_ASAP7_75t_L g5241 ( 
.A(n_4704),
.B(n_3982),
.Y(n_5241)
);

INVxp67_ASAP7_75t_L g5242 ( 
.A(n_4658),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_4326),
.Y(n_5243)
);

INVx2_ASAP7_75t_SL g5244 ( 
.A(n_4648),
.Y(n_5244)
);

OAI21x1_ASAP7_75t_L g5245 ( 
.A1(n_4312),
.A2(n_4017),
.B(n_4014),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_4326),
.Y(n_5246)
);

BUFx2_ASAP7_75t_L g5247 ( 
.A(n_4632),
.Y(n_5247)
);

INVx4_ASAP7_75t_L g5248 ( 
.A(n_4584),
.Y(n_5248)
);

INVx2_ASAP7_75t_L g5249 ( 
.A(n_4263),
.Y(n_5249)
);

OAI22x1_ASAP7_75t_SL g5250 ( 
.A1(n_4643),
.A2(n_3854),
.B1(n_3811),
.B2(n_3732),
.Y(n_5250)
);

BUFx3_ASAP7_75t_L g5251 ( 
.A(n_4671),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_4264),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4241),
.B(n_4031),
.Y(n_5253)
);

AOI21xp5_ASAP7_75t_L g5254 ( 
.A1(n_4405),
.A2(n_4486),
.B(n_4418),
.Y(n_5254)
);

INVx2_ASAP7_75t_SL g5255 ( 
.A(n_4482),
.Y(n_5255)
);

HB1xp67_ASAP7_75t_L g5256 ( 
.A(n_4414),
.Y(n_5256)
);

NOR2x1_ASAP7_75t_SL g5257 ( 
.A(n_4475),
.B(n_3892),
.Y(n_5257)
);

OAI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_4696),
.A2(n_3780),
.B1(n_3766),
.B2(n_3702),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_4334),
.Y(n_5259)
);

INVxp67_ASAP7_75t_L g5260 ( 
.A(n_4548),
.Y(n_5260)
);

OAI22xp33_ASAP7_75t_L g5261 ( 
.A1(n_4460),
.A2(n_4000),
.B1(n_4002),
.B2(n_3947),
.Y(n_5261)
);

INVx3_ASAP7_75t_SL g5262 ( 
.A(n_4364),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4334),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_4354),
.Y(n_5264)
);

AND2x2_ASAP7_75t_L g5265 ( 
.A(n_4704),
.B(n_4023),
.Y(n_5265)
);

INVx2_ASAP7_75t_SL g5266 ( 
.A(n_4482),
.Y(n_5266)
);

INVx3_ASAP7_75t_L g5267 ( 
.A(n_4247),
.Y(n_5267)
);

NAND2x1p5_ASAP7_75t_L g5268 ( 
.A(n_4402),
.B(n_4108),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_4256),
.B(n_4033),
.Y(n_5269)
);

OAI22xp5_ASAP7_75t_L g5270 ( 
.A1(n_4376),
.A2(n_4427),
.B1(n_4752),
.B2(n_4403),
.Y(n_5270)
);

AND2x2_ASAP7_75t_L g5271 ( 
.A(n_4228),
.B(n_4023),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_4354),
.Y(n_5272)
);

INVx2_ASAP7_75t_L g5273 ( 
.A(n_4264),
.Y(n_5273)
);

INVx2_ASAP7_75t_L g5274 ( 
.A(n_4264),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_4355),
.Y(n_5275)
);

OAI22xp33_ASAP7_75t_L g5276 ( 
.A1(n_4679),
.A2(n_4000),
.B1(n_4002),
.B2(n_3947),
.Y(n_5276)
);

BUFx6f_ASAP7_75t_L g5277 ( 
.A(n_4700),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4355),
.Y(n_5278)
);

BUFx2_ASAP7_75t_L g5279 ( 
.A(n_4724),
.Y(n_5279)
);

AND2x2_ASAP7_75t_L g5280 ( 
.A(n_4228),
.B(n_4023),
.Y(n_5280)
);

INVx4_ASAP7_75t_SL g5281 ( 
.A(n_4556),
.Y(n_5281)
);

INVx2_ASAP7_75t_L g5282 ( 
.A(n_4266),
.Y(n_5282)
);

AND2x2_ASAP7_75t_L g5283 ( 
.A(n_4272),
.B(n_4023),
.Y(n_5283)
);

AOI21x1_ASAP7_75t_L g5284 ( 
.A1(n_4456),
.A2(n_3842),
.B(n_3827),
.Y(n_5284)
);

OAI22xp5_ASAP7_75t_L g5285 ( 
.A1(n_4546),
.A2(n_4515),
.B1(n_4718),
.B2(n_4654),
.Y(n_5285)
);

OAI22xp33_ASAP7_75t_L g5286 ( 
.A1(n_4679),
.A2(n_4002),
.B1(n_4000),
.B2(n_3790),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_4369),
.Y(n_5287)
);

AOI22xp33_ASAP7_75t_L g5288 ( 
.A1(n_4419),
.A2(n_4002),
.B1(n_4000),
.B2(n_3850),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_4266),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_4414),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_4369),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_4266),
.Y(n_5292)
);

AOI21x1_ASAP7_75t_L g5293 ( 
.A1(n_4456),
.A2(n_3842),
.B(n_3827),
.Y(n_5293)
);

CKINVDCx20_ASAP7_75t_R g5294 ( 
.A(n_4307),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4371),
.Y(n_5295)
);

BUFx2_ASAP7_75t_L g5296 ( 
.A(n_4724),
.Y(n_5296)
);

INVx4_ASAP7_75t_L g5297 ( 
.A(n_4310),
.Y(n_5297)
);

INVx2_ASAP7_75t_SL g5298 ( 
.A(n_4482),
.Y(n_5298)
);

OAI21x1_ASAP7_75t_L g5299 ( 
.A1(n_4312),
.A2(n_4048),
.B(n_4017),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_4371),
.Y(n_5300)
);

BUFx12f_ASAP7_75t_L g5301 ( 
.A(n_4700),
.Y(n_5301)
);

INVx3_ASAP7_75t_L g5302 ( 
.A(n_4247),
.Y(n_5302)
);

AOI22xp33_ASAP7_75t_L g5303 ( 
.A1(n_4339),
.A2(n_3850),
.B1(n_3861),
.B2(n_3849),
.Y(n_5303)
);

AOI22xp33_ASAP7_75t_L g5304 ( 
.A1(n_4339),
.A2(n_3850),
.B1(n_3861),
.B2(n_3849),
.Y(n_5304)
);

HB1xp67_ASAP7_75t_L g5305 ( 
.A(n_4454),
.Y(n_5305)
);

INVx2_ASAP7_75t_L g5306 ( 
.A(n_4740),
.Y(n_5306)
);

BUFx3_ASAP7_75t_L g5307 ( 
.A(n_4671),
.Y(n_5307)
);

HB1xp67_ASAP7_75t_L g5308 ( 
.A(n_4454),
.Y(n_5308)
);

AND2x2_ASAP7_75t_L g5309 ( 
.A(n_4272),
.B(n_4274),
.Y(n_5309)
);

HB1xp67_ASAP7_75t_L g5310 ( 
.A(n_4489),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4384),
.Y(n_5311)
);

AO21x2_ASAP7_75t_L g5312 ( 
.A1(n_4545),
.A2(n_4189),
.B(n_4012),
.Y(n_5312)
);

BUFx6f_ASAP7_75t_L g5313 ( 
.A(n_4700),
.Y(n_5313)
);

BUFx3_ASAP7_75t_L g5314 ( 
.A(n_4671),
.Y(n_5314)
);

CKINVDCx11_ASAP7_75t_R g5315 ( 
.A(n_4548),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_4384),
.Y(n_5316)
);

AND2x2_ASAP7_75t_L g5317 ( 
.A(n_4272),
.B(n_4023),
.Y(n_5317)
);

INVx4_ASAP7_75t_L g5318 ( 
.A(n_4310),
.Y(n_5318)
);

AOI21x1_ASAP7_75t_L g5319 ( 
.A1(n_4524),
.A2(n_3862),
.B(n_3842),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_4274),
.B(n_4047),
.Y(n_5320)
);

BUFx6f_ASAP7_75t_L g5321 ( 
.A(n_4739),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_4740),
.Y(n_5322)
);

INVx2_ASAP7_75t_SL g5323 ( 
.A(n_4713),
.Y(n_5323)
);

INVxp67_ASAP7_75t_SL g5324 ( 
.A(n_4706),
.Y(n_5324)
);

AND2x4_ASAP7_75t_L g5325 ( 
.A(n_4364),
.B(n_4372),
.Y(n_5325)
);

INVx1_ASAP7_75t_SL g5326 ( 
.A(n_4489),
.Y(n_5326)
);

OAI21xp5_ASAP7_75t_SL g5327 ( 
.A1(n_4484),
.A2(n_3837),
.B(n_3829),
.Y(n_5327)
);

INVx3_ASAP7_75t_L g5328 ( 
.A(n_4247),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_4388),
.Y(n_5329)
);

INVx4_ASAP7_75t_L g5330 ( 
.A(n_4310),
.Y(n_5330)
);

NAND2x1p5_ASAP7_75t_L g5331 ( 
.A(n_4402),
.B(n_4115),
.Y(n_5331)
);

INVx2_ASAP7_75t_L g5332 ( 
.A(n_4740),
.Y(n_5332)
);

AOI21x1_ASAP7_75t_L g5333 ( 
.A1(n_4524),
.A2(n_3862),
.B(n_4189),
.Y(n_5333)
);

INVx2_ASAP7_75t_L g5334 ( 
.A(n_4275),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4388),
.Y(n_5335)
);

BUFx6f_ASAP7_75t_L g5336 ( 
.A(n_4739),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_4275),
.Y(n_5337)
);

AOI22xp33_ASAP7_75t_L g5338 ( 
.A1(n_4466),
.A2(n_3861),
.B1(n_3863),
.B2(n_3849),
.Y(n_5338)
);

HB1xp67_ASAP7_75t_L g5339 ( 
.A(n_4495),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_4389),
.Y(n_5340)
);

AOI22xp33_ASAP7_75t_SL g5341 ( 
.A1(n_4486),
.A2(n_3854),
.B1(n_3766),
.B2(n_3863),
.Y(n_5341)
);

AOI22xp33_ASAP7_75t_L g5342 ( 
.A1(n_4466),
.A2(n_3866),
.B1(n_3870),
.B2(n_3863),
.Y(n_5342)
);

AOI22xp33_ASAP7_75t_L g5343 ( 
.A1(n_4447),
.A2(n_3870),
.B1(n_3866),
.B2(n_3913),
.Y(n_5343)
);

AOI21x1_ASAP7_75t_L g5344 ( 
.A1(n_4365),
.A2(n_4719),
.B(n_4733),
.Y(n_5344)
);

INVx1_ASAP7_75t_SL g5345 ( 
.A(n_4495),
.Y(n_5345)
);

AOI22xp33_ASAP7_75t_L g5346 ( 
.A1(n_4447),
.A2(n_4418),
.B1(n_4423),
.B2(n_4387),
.Y(n_5346)
);

NOR2xp67_ASAP7_75t_SL g5347 ( 
.A(n_4321),
.B(n_3693),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_4389),
.Y(n_5348)
);

BUFx2_ASAP7_75t_L g5349 ( 
.A(n_4372),
.Y(n_5349)
);

CKINVDCx20_ASAP7_75t_R g5350 ( 
.A(n_4321),
.Y(n_5350)
);

HB1xp67_ASAP7_75t_L g5351 ( 
.A(n_4305),
.Y(n_5351)
);

INVx6_ASAP7_75t_L g5352 ( 
.A(n_4372),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_4275),
.Y(n_5353)
);

BUFx3_ASAP7_75t_L g5354 ( 
.A(n_4713),
.Y(n_5354)
);

OAI21x1_ASAP7_75t_L g5355 ( 
.A1(n_4312),
.A2(n_4048),
.B(n_4017),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_4288),
.Y(n_5356)
);

AND2x2_ASAP7_75t_L g5357 ( 
.A(n_4274),
.B(n_4047),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_4288),
.Y(n_5358)
);

OAI22xp5_ASAP7_75t_L g5359 ( 
.A1(n_4654),
.A2(n_3702),
.B1(n_3717),
.B2(n_3693),
.Y(n_5359)
);

CKINVDCx20_ASAP7_75t_R g5360 ( 
.A(n_4321),
.Y(n_5360)
);

AOI22xp33_ASAP7_75t_L g5361 ( 
.A1(n_4447),
.A2(n_3870),
.B1(n_3866),
.B2(n_3913),
.Y(n_5361)
);

AOI22xp33_ASAP7_75t_L g5362 ( 
.A1(n_4447),
.A2(n_3924),
.B1(n_3953),
.B2(n_3913),
.Y(n_5362)
);

OAI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_4689),
.A2(n_3702),
.B1(n_3717),
.B2(n_3693),
.Y(n_5363)
);

INVx2_ASAP7_75t_SL g5364 ( 
.A(n_4713),
.Y(n_5364)
);

BUFx12f_ASAP7_75t_L g5365 ( 
.A(n_4338),
.Y(n_5365)
);

INVx2_ASAP7_75t_L g5366 ( 
.A(n_4288),
.Y(n_5366)
);

HB1xp67_ASAP7_75t_L g5367 ( 
.A(n_4305),
.Y(n_5367)
);

AOI22xp33_ASAP7_75t_L g5368 ( 
.A1(n_4447),
.A2(n_3953),
.B1(n_3962),
.B2(n_3924),
.Y(n_5368)
);

AOI22xp33_ASAP7_75t_L g5369 ( 
.A1(n_4387),
.A2(n_3953),
.B1(n_3962),
.B2(n_3924),
.Y(n_5369)
);

AND2x2_ASAP7_75t_L g5370 ( 
.A(n_4467),
.B(n_4047),
.Y(n_5370)
);

AOI22xp5_ASAP7_75t_SL g5371 ( 
.A1(n_4484),
.A2(n_3719),
.B1(n_3722),
.B2(n_3717),
.Y(n_5371)
);

OAI21x1_ASAP7_75t_SL g5372 ( 
.A1(n_4506),
.A2(n_3684),
.B(n_3683),
.Y(n_5372)
);

INVx3_ASAP7_75t_SL g5373 ( 
.A(n_4372),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_4555),
.B(n_4033),
.Y(n_5374)
);

AOI22xp33_ASAP7_75t_L g5375 ( 
.A1(n_4423),
.A2(n_3978),
.B1(n_3988),
.B2(n_3962),
.Y(n_5375)
);

BUFx2_ASAP7_75t_SL g5376 ( 
.A(n_4283),
.Y(n_5376)
);

OAI21xp5_ASAP7_75t_SL g5377 ( 
.A1(n_4501),
.A2(n_3837),
.B(n_3829),
.Y(n_5377)
);

OAI22xp33_ASAP7_75t_L g5378 ( 
.A1(n_4402),
.A2(n_3790),
.B1(n_3793),
.B2(n_3776),
.Y(n_5378)
);

AOI22xp33_ASAP7_75t_SL g5379 ( 
.A1(n_4501),
.A2(n_4402),
.B1(n_4431),
.B2(n_4410),
.Y(n_5379)
);

OAI21xp5_ASAP7_75t_L g5380 ( 
.A1(n_4330),
.A2(n_3998),
.B(n_3976),
.Y(n_5380)
);

INVx4_ASAP7_75t_L g5381 ( 
.A(n_4338),
.Y(n_5381)
);

NOR2xp33_ASAP7_75t_L g5382 ( 
.A(n_4661),
.B(n_3724),
.Y(n_5382)
);

INVx3_ASAP7_75t_SL g5383 ( 
.A(n_4372),
.Y(n_5383)
);

HB1xp67_ASAP7_75t_L g5384 ( 
.A(n_4331),
.Y(n_5384)
);

BUFx12f_ASAP7_75t_L g5385 ( 
.A(n_4338),
.Y(n_5385)
);

INVx1_ASAP7_75t_SL g5386 ( 
.A(n_4555),
.Y(n_5386)
);

INVx3_ASAP7_75t_L g5387 ( 
.A(n_4247),
.Y(n_5387)
);

OAI22xp33_ASAP7_75t_L g5388 ( 
.A1(n_4402),
.A2(n_3790),
.B1(n_3793),
.B2(n_3776),
.Y(n_5388)
);

HB1xp67_ASAP7_75t_L g5389 ( 
.A(n_4331),
.Y(n_5389)
);

BUFx4f_ASAP7_75t_SL g5390 ( 
.A(n_4564),
.Y(n_5390)
);

INVx2_ASAP7_75t_SL g5391 ( 
.A(n_4622),
.Y(n_5391)
);

AND2x2_ASAP7_75t_L g5392 ( 
.A(n_4467),
.B(n_4533),
.Y(n_5392)
);

BUFx2_ASAP7_75t_L g5393 ( 
.A(n_4412),
.Y(n_5393)
);

AO21x1_ASAP7_75t_SL g5394 ( 
.A1(n_4575),
.A2(n_4131),
.B(n_4128),
.Y(n_5394)
);

OAI22xp5_ASAP7_75t_L g5395 ( 
.A1(n_4549),
.A2(n_3722),
.B1(n_3736),
.B2(n_3719),
.Y(n_5395)
);

AOI21x1_ASAP7_75t_L g5396 ( 
.A1(n_4365),
.A2(n_3862),
.B(n_4189),
.Y(n_5396)
);

BUFx2_ASAP7_75t_R g5397 ( 
.A(n_4665),
.Y(n_5397)
);

BUFx2_ASAP7_75t_L g5398 ( 
.A(n_4412),
.Y(n_5398)
);

BUFx6f_ASAP7_75t_L g5399 ( 
.A(n_4739),
.Y(n_5399)
);

BUFx8_ASAP7_75t_L g5400 ( 
.A(n_4425),
.Y(n_5400)
);

BUFx3_ASAP7_75t_L g5401 ( 
.A(n_4506),
.Y(n_5401)
);

AND2x2_ASAP7_75t_L g5402 ( 
.A(n_4467),
.B(n_4533),
.Y(n_5402)
);

INVx4_ASAP7_75t_L g5403 ( 
.A(n_4412),
.Y(n_5403)
);

AO21x2_ASAP7_75t_L g5404 ( 
.A1(n_4497),
.A2(n_4189),
.B(n_4012),
.Y(n_5404)
);

AOI21x1_ASAP7_75t_L g5405 ( 
.A1(n_4719),
.A2(n_4733),
.B(n_4216),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4438),
.Y(n_5406)
);

HB1xp67_ASAP7_75t_L g5407 ( 
.A(n_4350),
.Y(n_5407)
);

NAND2xp5_ASAP7_75t_L g5408 ( 
.A(n_4564),
.B(n_4036),
.Y(n_5408)
);

OAI21xp5_ASAP7_75t_L g5409 ( 
.A1(n_4508),
.A2(n_3998),
.B(n_4016),
.Y(n_5409)
);

INVx3_ASAP7_75t_L g5410 ( 
.A(n_4270),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_4445),
.Y(n_5411)
);

OA21x2_ASAP7_75t_L g5412 ( 
.A1(n_4400),
.A2(n_4015),
.B(n_4003),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_4363),
.Y(n_5413)
);

INVx4_ASAP7_75t_L g5414 ( 
.A(n_4412),
.Y(n_5414)
);

AOI21x1_ASAP7_75t_L g5415 ( 
.A1(n_4197),
.A2(n_4142),
.B(n_4137),
.Y(n_5415)
);

BUFx3_ASAP7_75t_L g5416 ( 
.A(n_4739),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_4445),
.Y(n_5417)
);

AOI22xp33_ASAP7_75t_L g5418 ( 
.A1(n_4431),
.A2(n_3988),
.B1(n_3991),
.B2(n_3978),
.Y(n_5418)
);

AND2x4_ASAP7_75t_L g5419 ( 
.A(n_4412),
.B(n_4472),
.Y(n_5419)
);

AOI22xp33_ASAP7_75t_L g5420 ( 
.A1(n_4577),
.A2(n_3988),
.B1(n_3991),
.B2(n_3978),
.Y(n_5420)
);

OAI22xp33_ASAP7_75t_L g5421 ( 
.A1(n_4402),
.A2(n_3793),
.B1(n_3995),
.B2(n_3991),
.Y(n_5421)
);

HB1xp67_ASAP7_75t_L g5422 ( 
.A(n_4350),
.Y(n_5422)
);

AND2x2_ASAP7_75t_L g5423 ( 
.A(n_4467),
.B(n_4047),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_4446),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_4446),
.Y(n_5425)
);

AOI22xp5_ASAP7_75t_L g5426 ( 
.A1(n_4511),
.A2(n_3722),
.B1(n_3736),
.B2(n_3719),
.Y(n_5426)
);

NAND2xp5_ASAP7_75t_L g5427 ( 
.A(n_4566),
.B(n_4036),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_4458),
.Y(n_5428)
);

AOI22xp33_ASAP7_75t_L g5429 ( 
.A1(n_4577),
.A2(n_3999),
.B1(n_4001),
.B2(n_3995),
.Y(n_5429)
);

AOI22xp33_ASAP7_75t_L g5430 ( 
.A1(n_4434),
.A2(n_3999),
.B1(n_4001),
.B2(n_3995),
.Y(n_5430)
);

BUFx3_ASAP7_75t_L g5431 ( 
.A(n_4675),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_4775),
.Y(n_5432)
);

INVx2_ASAP7_75t_SL g5433 ( 
.A(n_4783),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_4775),
.Y(n_5434)
);

INVx3_ASAP7_75t_L g5435 ( 
.A(n_5325),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_4777),
.Y(n_5436)
);

HB1xp67_ASAP7_75t_L g5437 ( 
.A(n_4907),
.Y(n_5437)
);

AND2x2_ASAP7_75t_L g5438 ( 
.A(n_4834),
.B(n_4304),
.Y(n_5438)
);

INVx2_ASAP7_75t_L g5439 ( 
.A(n_4785),
.Y(n_5439)
);

INVx2_ASAP7_75t_SL g5440 ( 
.A(n_4783),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_L g5441 ( 
.A(n_5056),
.B(n_4566),
.Y(n_5441)
);

INVx2_ASAP7_75t_SL g5442 ( 
.A(n_4783),
.Y(n_5442)
);

INVx2_ASAP7_75t_SL g5443 ( 
.A(n_4783),
.Y(n_5443)
);

HB1xp67_ASAP7_75t_L g5444 ( 
.A(n_4914),
.Y(n_5444)
);

BUFx2_ASAP7_75t_L g5445 ( 
.A(n_4960),
.Y(n_5445)
);

INVx2_ASAP7_75t_L g5446 ( 
.A(n_4785),
.Y(n_5446)
);

AND2x4_ASAP7_75t_L g5447 ( 
.A(n_5281),
.B(n_4472),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_4777),
.Y(n_5448)
);

INVx3_ASAP7_75t_L g5449 ( 
.A(n_5325),
.Y(n_5449)
);

INVx2_ASAP7_75t_L g5450 ( 
.A(n_4785),
.Y(n_5450)
);

OR2x2_ASAP7_75t_L g5451 ( 
.A(n_4971),
.B(n_4441),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_4780),
.Y(n_5452)
);

INVxp67_ASAP7_75t_L g5453 ( 
.A(n_5079),
.Y(n_5453)
);

INVxp67_ASAP7_75t_L g5454 ( 
.A(n_5078),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_4780),
.Y(n_5455)
);

NAND2xp5_ASAP7_75t_L g5456 ( 
.A(n_5228),
.B(n_4583),
.Y(n_5456)
);

INVx2_ASAP7_75t_SL g5457 ( 
.A(n_4783),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_4789),
.Y(n_5458)
);

INVx3_ASAP7_75t_L g5459 ( 
.A(n_5325),
.Y(n_5459)
);

INVx2_ASAP7_75t_L g5460 ( 
.A(n_4789),
.Y(n_5460)
);

INVx2_ASAP7_75t_L g5461 ( 
.A(n_4789),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_4793),
.Y(n_5462)
);

INVx2_ASAP7_75t_L g5463 ( 
.A(n_4793),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_4786),
.Y(n_5464)
);

INVx3_ASAP7_75t_L g5465 ( 
.A(n_5325),
.Y(n_5465)
);

OAI21x1_ASAP7_75t_L g5466 ( 
.A1(n_5333),
.A2(n_4553),
.B(n_4562),
.Y(n_5466)
);

BUFx3_ASAP7_75t_L g5467 ( 
.A(n_4848),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_4786),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_4788),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_4788),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_4793),
.Y(n_5471)
);

INVxp67_ASAP7_75t_L g5472 ( 
.A(n_5126),
.Y(n_5472)
);

BUFx2_ASAP7_75t_L g5473 ( 
.A(n_4960),
.Y(n_5473)
);

INVx2_ASAP7_75t_L g5474 ( 
.A(n_4803),
.Y(n_5474)
);

OAI21xp5_ASAP7_75t_L g5475 ( 
.A1(n_4801),
.A2(n_4508),
.B(n_4730),
.Y(n_5475)
);

INVx3_ASAP7_75t_L g5476 ( 
.A(n_5419),
.Y(n_5476)
);

OA21x2_ASAP7_75t_L g5477 ( 
.A1(n_4830),
.A2(n_4380),
.B(n_4453),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_4794),
.Y(n_5478)
);

INVx8_ASAP7_75t_L g5479 ( 
.A(n_4812),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_4794),
.Y(n_5480)
);

NAND2xp5_ASAP7_75t_L g5481 ( 
.A(n_5077),
.B(n_4583),
.Y(n_5481)
);

OAI21x1_ASAP7_75t_L g5482 ( 
.A1(n_5333),
.A2(n_4553),
.B(n_4562),
.Y(n_5482)
);

OAI21x1_ASAP7_75t_L g5483 ( 
.A1(n_5319),
.A2(n_4553),
.B(n_4562),
.Y(n_5483)
);

INVxp67_ASAP7_75t_L g5484 ( 
.A(n_5211),
.Y(n_5484)
);

INVx2_ASAP7_75t_L g5485 ( 
.A(n_4803),
.Y(n_5485)
);

AO21x2_ASAP7_75t_L g5486 ( 
.A1(n_4847),
.A2(n_4497),
.B(n_4273),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_4797),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_4803),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_4797),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_4800),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_4815),
.Y(n_5491)
);

AO21x2_ASAP7_75t_L g5492 ( 
.A1(n_4847),
.A2(n_4273),
.B(n_4243),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_4800),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_4815),
.Y(n_5494)
);

INVx2_ASAP7_75t_L g5495 ( 
.A(n_4815),
.Y(n_5495)
);

NAND2x1p5_ASAP7_75t_L g5496 ( 
.A(n_5023),
.B(n_4289),
.Y(n_5496)
);

INVx2_ASAP7_75t_L g5497 ( 
.A(n_4760),
.Y(n_5497)
);

INVx3_ASAP7_75t_L g5498 ( 
.A(n_5419),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_4802),
.Y(n_5499)
);

BUFx2_ASAP7_75t_L g5500 ( 
.A(n_4960),
.Y(n_5500)
);

CKINVDCx5p33_ASAP7_75t_R g5501 ( 
.A(n_4825),
.Y(n_5501)
);

BUFx3_ASAP7_75t_L g5502 ( 
.A(n_4848),
.Y(n_5502)
);

INVx3_ASAP7_75t_L g5503 ( 
.A(n_5419),
.Y(n_5503)
);

INVx1_ASAP7_75t_L g5504 ( 
.A(n_4802),
.Y(n_5504)
);

AO21x2_ASAP7_75t_L g5505 ( 
.A1(n_4880),
.A2(n_4243),
.B(n_4673),
.Y(n_5505)
);

OR2x2_ASAP7_75t_L g5506 ( 
.A(n_4971),
.B(n_4441),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_4807),
.Y(n_5507)
);

INVx2_ASAP7_75t_L g5508 ( 
.A(n_4760),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_4807),
.Y(n_5509)
);

AO21x2_ASAP7_75t_L g5510 ( 
.A1(n_4880),
.A2(n_4673),
.B(n_4543),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_5242),
.B(n_4636),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_4760),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_4809),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_4809),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_4769),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_4822),
.Y(n_5516)
);

INVx1_ASAP7_75t_SL g5517 ( 
.A(n_4986),
.Y(n_5517)
);

OR2x2_ASAP7_75t_L g5518 ( 
.A(n_5031),
.B(n_4441),
.Y(n_5518)
);

INVx3_ASAP7_75t_L g5519 ( 
.A(n_5419),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_4769),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_4822),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_4826),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_4826),
.Y(n_5523)
);

AND2x2_ASAP7_75t_L g5524 ( 
.A(n_4834),
.B(n_4970),
.Y(n_5524)
);

AND2x2_ASAP7_75t_L g5525 ( 
.A(n_4970),
.B(n_4304),
.Y(n_5525)
);

OR2x2_ASAP7_75t_L g5526 ( 
.A(n_5031),
.B(n_4441),
.Y(n_5526)
);

INVx3_ASAP7_75t_L g5527 ( 
.A(n_4960),
.Y(n_5527)
);

OR2x2_ASAP7_75t_L g5528 ( 
.A(n_5002),
.B(n_4222),
.Y(n_5528)
);

INVx2_ASAP7_75t_SL g5529 ( 
.A(n_5062),
.Y(n_5529)
);

O2A1O1Ixp33_ASAP7_75t_L g5530 ( 
.A1(n_5160),
.A2(n_4754),
.B(n_4514),
.C(n_4565),
.Y(n_5530)
);

INVx2_ASAP7_75t_L g5531 ( 
.A(n_4769),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_4831),
.Y(n_5532)
);

BUFx6f_ASAP7_75t_L g5533 ( 
.A(n_4812),
.Y(n_5533)
);

AOI22xp5_ASAP7_75t_L g5534 ( 
.A1(n_4832),
.A2(n_4623),
.B1(n_4619),
.B2(n_4523),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_4831),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_4840),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_4840),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_4841),
.Y(n_5538)
);

INVxp67_ASAP7_75t_SL g5539 ( 
.A(n_4824),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_4841),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_4774),
.Y(n_5541)
);

HB1xp67_ASAP7_75t_L g5542 ( 
.A(n_4806),
.Y(n_5542)
);

BUFx3_ASAP7_75t_L g5543 ( 
.A(n_4848),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_4842),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_4774),
.Y(n_5545)
);

OR2x2_ASAP7_75t_L g5546 ( 
.A(n_5094),
.B(n_5324),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_4774),
.Y(n_5547)
);

OAI22xp5_ASAP7_75t_L g5548 ( 
.A1(n_4863),
.A2(n_4865),
.B1(n_4832),
.B2(n_5050),
.Y(n_5548)
);

BUFx2_ASAP7_75t_R g5549 ( 
.A(n_5080),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_4776),
.Y(n_5550)
);

OAI21x1_ASAP7_75t_L g5551 ( 
.A1(n_5319),
.A2(n_5293),
.B(n_5284),
.Y(n_5551)
);

INVx2_ASAP7_75t_L g5552 ( 
.A(n_4776),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4842),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_4845),
.Y(n_5554)
);

NOR2xp33_ASAP7_75t_L g5555 ( 
.A(n_4759),
.B(n_3682),
.Y(n_5555)
);

AND2x2_ASAP7_75t_L g5556 ( 
.A(n_4850),
.B(n_4304),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4845),
.Y(n_5557)
);

CKINVDCx8_ASAP7_75t_R g5558 ( 
.A(n_4951),
.Y(n_5558)
);

INVx2_ASAP7_75t_L g5559 ( 
.A(n_4776),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4858),
.Y(n_5560)
);

NAND2xp5_ASAP7_75t_L g5561 ( 
.A(n_4765),
.B(n_4823),
.Y(n_5561)
);

AND2x2_ASAP7_75t_L g5562 ( 
.A(n_4850),
.B(n_4311),
.Y(n_5562)
);

BUFx6f_ASAP7_75t_L g5563 ( 
.A(n_4812),
.Y(n_5563)
);

OAI21x1_ASAP7_75t_L g5564 ( 
.A1(n_5284),
.A2(n_4576),
.B(n_4453),
.Y(n_5564)
);

OAI21x1_ASAP7_75t_L g5565 ( 
.A1(n_5293),
.A2(n_4576),
.B(n_4453),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_4858),
.Y(n_5566)
);

AND2x2_ASAP7_75t_L g5567 ( 
.A(n_5392),
.B(n_4311),
.Y(n_5567)
);

BUFx2_ASAP7_75t_L g5568 ( 
.A(n_5349),
.Y(n_5568)
);

INVx2_ASAP7_75t_SL g5569 ( 
.A(n_5062),
.Y(n_5569)
);

AND2x2_ASAP7_75t_L g5570 ( 
.A(n_5392),
.B(n_4311),
.Y(n_5570)
);

OAI21x1_ASAP7_75t_L g5571 ( 
.A1(n_5044),
.A2(n_4576),
.B(n_4510),
.Y(n_5571)
);

CKINVDCx5p33_ASAP7_75t_R g5572 ( 
.A(n_4782),
.Y(n_5572)
);

BUFx2_ASAP7_75t_L g5573 ( 
.A(n_5349),
.Y(n_5573)
);

AND2x6_ASAP7_75t_L g5574 ( 
.A(n_5223),
.B(n_4499),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_4870),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_4779),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_4779),
.Y(n_5577)
);

INVx2_ASAP7_75t_L g5578 ( 
.A(n_4779),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_L g5579 ( 
.A(n_4869),
.B(n_4897),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_4870),
.Y(n_5580)
);

INVx2_ASAP7_75t_L g5581 ( 
.A(n_5058),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_4873),
.Y(n_5582)
);

INVx2_ASAP7_75t_L g5583 ( 
.A(n_5058),
.Y(n_5583)
);

AO21x2_ASAP7_75t_L g5584 ( 
.A1(n_5117),
.A2(n_4543),
.B(n_4605),
.Y(n_5584)
);

AND2x2_ASAP7_75t_L g5585 ( 
.A(n_5402),
.B(n_4337),
.Y(n_5585)
);

BUFx12f_ASAP7_75t_L g5586 ( 
.A(n_4848),
.Y(n_5586)
);

AND2x2_ASAP7_75t_L g5587 ( 
.A(n_5402),
.B(n_4337),
.Y(n_5587)
);

INVx2_ASAP7_75t_L g5588 ( 
.A(n_5058),
.Y(n_5588)
);

INVx2_ASAP7_75t_L g5589 ( 
.A(n_5066),
.Y(n_5589)
);

BUFx3_ASAP7_75t_L g5590 ( 
.A(n_4871),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_4873),
.Y(n_5591)
);

OAI21xp5_ASAP7_75t_L g5592 ( 
.A1(n_5160),
.A2(n_4730),
.B(n_4216),
.Y(n_5592)
);

OAI22xp5_ASAP7_75t_L g5593 ( 
.A1(n_5050),
.A2(n_4612),
.B1(n_4644),
.B2(n_4550),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_4876),
.Y(n_5594)
);

NOR2x1_ASAP7_75t_R g5595 ( 
.A(n_4922),
.B(n_3724),
.Y(n_5595)
);

HB1xp67_ASAP7_75t_L g5596 ( 
.A(n_4846),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_4876),
.Y(n_5597)
);

BUFx12f_ASAP7_75t_L g5598 ( 
.A(n_4871),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5066),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_4885),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5260),
.B(n_4636),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_4885),
.Y(n_5602)
);

OAI21x1_ASAP7_75t_L g5603 ( 
.A1(n_5044),
.A2(n_4510),
.B(n_4731),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_4887),
.Y(n_5604)
);

INVx2_ASAP7_75t_L g5605 ( 
.A(n_5066),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_4887),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_4890),
.Y(n_5607)
);

AOI21x1_ASAP7_75t_L g5608 ( 
.A1(n_4829),
.A2(n_4755),
.B(n_4677),
.Y(n_5608)
);

INVx2_ASAP7_75t_L g5609 ( 
.A(n_5103),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_4890),
.Y(n_5610)
);

INVx2_ASAP7_75t_L g5611 ( 
.A(n_5103),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5103),
.Y(n_5612)
);

HB1xp67_ASAP7_75t_L g5613 ( 
.A(n_4874),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_5104),
.Y(n_5614)
);

AND2x4_ASAP7_75t_L g5615 ( 
.A(n_5281),
.B(n_4472),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_4891),
.Y(n_5616)
);

INVx2_ASAP7_75t_L g5617 ( 
.A(n_5104),
.Y(n_5617)
);

AOI22xp33_ASAP7_75t_L g5618 ( 
.A1(n_4993),
.A2(n_4410),
.B1(n_4523),
.B2(n_4434),
.Y(n_5618)
);

OR2x2_ASAP7_75t_L g5619 ( 
.A(n_5217),
.B(n_4222),
.Y(n_5619)
);

AND2x2_ASAP7_75t_L g5620 ( 
.A(n_5174),
.B(n_4337),
.Y(n_5620)
);

BUFx2_ASAP7_75t_L g5621 ( 
.A(n_5393),
.Y(n_5621)
);

INVx2_ASAP7_75t_SL g5622 ( 
.A(n_5062),
.Y(n_5622)
);

OR2x2_ASAP7_75t_L g5623 ( 
.A(n_5217),
.B(n_4449),
.Y(n_5623)
);

AND2x2_ASAP7_75t_L g5624 ( 
.A(n_5174),
.B(n_4357),
.Y(n_5624)
);

BUFx2_ASAP7_75t_L g5625 ( 
.A(n_5393),
.Y(n_5625)
);

OAI21x1_ASAP7_75t_L g5626 ( 
.A1(n_5093),
.A2(n_4510),
.B(n_4731),
.Y(n_5626)
);

OAI21x1_ASAP7_75t_L g5627 ( 
.A1(n_5093),
.A2(n_4736),
.B(n_4731),
.Y(n_5627)
);

INVx2_ASAP7_75t_L g5628 ( 
.A(n_5104),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5107),
.Y(n_5629)
);

INVx3_ASAP7_75t_L g5630 ( 
.A(n_5062),
.Y(n_5630)
);

OR2x2_ASAP7_75t_L g5631 ( 
.A(n_5060),
.B(n_4449),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_4891),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_5107),
.Y(n_5633)
);

NAND2xp5_ASAP7_75t_L g5634 ( 
.A(n_4929),
.B(n_4646),
.Y(n_5634)
);

AND2x2_ASAP7_75t_L g5635 ( 
.A(n_5370),
.B(n_4357),
.Y(n_5635)
);

AND2x2_ASAP7_75t_L g5636 ( 
.A(n_5370),
.B(n_4357),
.Y(n_5636)
);

HB1xp67_ASAP7_75t_L g5637 ( 
.A(n_4877),
.Y(n_5637)
);

AND2x2_ASAP7_75t_L g5638 ( 
.A(n_5423),
.B(n_4374),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_4892),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_4892),
.Y(n_5640)
);

HB1xp67_ASAP7_75t_L g5641 ( 
.A(n_5214),
.Y(n_5641)
);

OAI21xp5_ASAP7_75t_L g5642 ( 
.A1(n_5254),
.A2(n_4197),
.B(n_4265),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_4893),
.Y(n_5643)
);

OAI21x1_ASAP7_75t_L g5644 ( 
.A1(n_5166),
.A2(n_4736),
.B(n_4380),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_5107),
.Y(n_5645)
);

INVx2_ASAP7_75t_L g5646 ( 
.A(n_5109),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_5109),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_4893),
.Y(n_5648)
);

HB1xp67_ASAP7_75t_L g5649 ( 
.A(n_5220),
.Y(n_5649)
);

AND2x2_ASAP7_75t_L g5650 ( 
.A(n_5423),
.B(n_4965),
.Y(n_5650)
);

AO21x2_ASAP7_75t_L g5651 ( 
.A1(n_5117),
.A2(n_4605),
.B(n_4301),
.Y(n_5651)
);

INVx2_ASAP7_75t_SL g5652 ( 
.A(n_5062),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_4895),
.Y(n_5653)
);

INVx5_ASAP7_75t_L g5654 ( 
.A(n_4836),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_4895),
.Y(n_5655)
);

NAND2xp5_ASAP7_75t_L g5656 ( 
.A(n_5386),
.B(n_4646),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_4909),
.Y(n_5657)
);

INVx2_ASAP7_75t_L g5658 ( 
.A(n_4827),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_4909),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_4827),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_4827),
.Y(n_5661)
);

HB1xp67_ASAP7_75t_L g5662 ( 
.A(n_5227),
.Y(n_5662)
);

INVx1_ASAP7_75t_SL g5663 ( 
.A(n_5315),
.Y(n_5663)
);

INVx2_ASAP7_75t_L g5664 ( 
.A(n_4838),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_4913),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_4913),
.Y(n_5666)
);

HB1xp67_ASAP7_75t_L g5667 ( 
.A(n_5256),
.Y(n_5667)
);

OAI22xp5_ASAP7_75t_L g5668 ( 
.A1(n_5426),
.A2(n_4554),
.B1(n_4593),
.B2(n_4600),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_4838),
.Y(n_5669)
);

CKINVDCx14_ASAP7_75t_R g5670 ( 
.A(n_5115),
.Y(n_5670)
);

AND2x2_ASAP7_75t_L g5671 ( 
.A(n_4965),
.B(n_4374),
.Y(n_5671)
);

HB1xp67_ASAP7_75t_L g5672 ( 
.A(n_5290),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_4838),
.Y(n_5673)
);

NAND2x1p5_ASAP7_75t_L g5674 ( 
.A(n_5023),
.B(n_4289),
.Y(n_5674)
);

BUFx2_ASAP7_75t_L g5675 ( 
.A(n_5398),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_4916),
.Y(n_5676)
);

BUFx2_ASAP7_75t_L g5677 ( 
.A(n_5398),
.Y(n_5677)
);

INVx3_ASAP7_75t_L g5678 ( 
.A(n_5352),
.Y(n_5678)
);

BUFx2_ASAP7_75t_L g5679 ( 
.A(n_5400),
.Y(n_5679)
);

INVx2_ASAP7_75t_L g5680 ( 
.A(n_4839),
.Y(n_5680)
);

CKINVDCx5p33_ASAP7_75t_R g5681 ( 
.A(n_4864),
.Y(n_5681)
);

OR2x2_ASAP7_75t_L g5682 ( 
.A(n_5060),
.B(n_4534),
.Y(n_5682)
);

AND2x2_ASAP7_75t_L g5683 ( 
.A(n_5020),
.B(n_4374),
.Y(n_5683)
);

HB1xp67_ASAP7_75t_L g5684 ( 
.A(n_5305),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_4916),
.Y(n_5685)
);

OAI21xp5_ASAP7_75t_L g5686 ( 
.A1(n_5346),
.A2(n_4293),
.B(n_4265),
.Y(n_5686)
);

AND2x2_ASAP7_75t_L g5687 ( 
.A(n_5020),
.B(n_4379),
.Y(n_5687)
);

INVx2_ASAP7_75t_L g5688 ( 
.A(n_4839),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_4920),
.Y(n_5689)
);

INVxp67_ASAP7_75t_L g5690 ( 
.A(n_5308),
.Y(n_5690)
);

INVx2_ASAP7_75t_L g5691 ( 
.A(n_4839),
.Y(n_5691)
);

INVx2_ASAP7_75t_L g5692 ( 
.A(n_4843),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_4920),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_4924),
.Y(n_5694)
);

AND2x4_ASAP7_75t_L g5695 ( 
.A(n_5281),
.B(n_4472),
.Y(n_5695)
);

HB1xp67_ASAP7_75t_L g5696 ( 
.A(n_5310),
.Y(n_5696)
);

INVx2_ASAP7_75t_L g5697 ( 
.A(n_4843),
.Y(n_5697)
);

AND2x4_ASAP7_75t_L g5698 ( 
.A(n_5281),
.B(n_4472),
.Y(n_5698)
);

AOI22xp5_ASAP7_75t_L g5699 ( 
.A1(n_5231),
.A2(n_4623),
.B1(n_4619),
.B2(n_4410),
.Y(n_5699)
);

INVxp67_ASAP7_75t_SL g5700 ( 
.A(n_4824),
.Y(n_5700)
);

INVx2_ASAP7_75t_L g5701 ( 
.A(n_4843),
.Y(n_5701)
);

INVx3_ASAP7_75t_L g5702 ( 
.A(n_5352),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_4924),
.Y(n_5703)
);

BUFx3_ASAP7_75t_L g5704 ( 
.A(n_4871),
.Y(n_5704)
);

NAND2x1_ASAP7_75t_L g5705 ( 
.A(n_5372),
.B(n_4631),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_4936),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_L g5707 ( 
.A(n_5386),
.B(n_4663),
.Y(n_5707)
);

HB1xp67_ASAP7_75t_L g5708 ( 
.A(n_5339),
.Y(n_5708)
);

INVx2_ASAP7_75t_L g5709 ( 
.A(n_4844),
.Y(n_5709)
);

INVx3_ASAP7_75t_L g5710 ( 
.A(n_5352),
.Y(n_5710)
);

BUFx2_ASAP7_75t_L g5711 ( 
.A(n_5400),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_4844),
.Y(n_5712)
);

INVx2_ASAP7_75t_L g5713 ( 
.A(n_4844),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_4936),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_4938),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_4938),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_4940),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5412),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_4940),
.Y(n_5719)
);

INVx2_ASAP7_75t_SL g5720 ( 
.A(n_5352),
.Y(n_5720)
);

OAI21xp5_ASAP7_75t_L g5721 ( 
.A1(n_4953),
.A2(n_4328),
.B(n_4293),
.Y(n_5721)
);

AND2x4_ASAP7_75t_L g5722 ( 
.A(n_5281),
.B(n_4289),
.Y(n_5722)
);

INVx2_ASAP7_75t_L g5723 ( 
.A(n_5412),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_4945),
.Y(n_5724)
);

INVx2_ASAP7_75t_L g5725 ( 
.A(n_5412),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_4945),
.Y(n_5726)
);

AO21x1_ASAP7_75t_L g5727 ( 
.A1(n_5380),
.A2(n_4716),
.B(n_4686),
.Y(n_5727)
);

INVx3_ASAP7_75t_L g5728 ( 
.A(n_5352),
.Y(n_5728)
);

AOI22xp33_ASAP7_75t_L g5729 ( 
.A1(n_5400),
.A2(n_4410),
.B1(n_4356),
.B2(n_4541),
.Y(n_5729)
);

OAI21x1_ASAP7_75t_L g5730 ( 
.A1(n_5166),
.A2(n_4736),
.B(n_4380),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_5412),
.Y(n_5731)
);

OR2x2_ASAP7_75t_L g5732 ( 
.A(n_4928),
.B(n_4534),
.Y(n_5732)
);

INVx2_ASAP7_75t_SL g5733 ( 
.A(n_5101),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_4955),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_5007),
.Y(n_5735)
);

AOI21x1_ASAP7_75t_L g5736 ( 
.A1(n_4829),
.A2(n_4755),
.B(n_4677),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_5109),
.Y(n_5737)
);

BUFx3_ASAP7_75t_L g5738 ( 
.A(n_4871),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_4955),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_4961),
.Y(n_5740)
);

OAI21x1_ASAP7_75t_L g5741 ( 
.A1(n_5396),
.A2(n_4470),
.B(n_4594),
.Y(n_5741)
);

INVx1_ASAP7_75t_L g5742 ( 
.A(n_4961),
.Y(n_5742)
);

OAI21x1_ASAP7_75t_L g5743 ( 
.A1(n_5396),
.A2(n_4470),
.B(n_4594),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5116),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_4967),
.Y(n_5745)
);

OA21x2_ASAP7_75t_L g5746 ( 
.A1(n_4830),
.A2(n_4299),
.B(n_4298),
.Y(n_5746)
);

INVx2_ASAP7_75t_L g5747 ( 
.A(n_5116),
.Y(n_5747)
);

NAND2xp5_ASAP7_75t_L g5748 ( 
.A(n_4904),
.B(n_4663),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5116),
.Y(n_5749)
);

HB1xp67_ASAP7_75t_L g5750 ( 
.A(n_5085),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5121),
.Y(n_5751)
);

HB1xp67_ASAP7_75t_L g5752 ( 
.A(n_5085),
.Y(n_5752)
);

NOR2xp33_ASAP7_75t_L g5753 ( 
.A(n_4759),
.B(n_3682),
.Y(n_5753)
);

INVx1_ASAP7_75t_SL g5754 ( 
.A(n_5397),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_4967),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_4972),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5121),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5121),
.Y(n_5758)
);

BUFx2_ASAP7_75t_SL g5759 ( 
.A(n_5045),
.Y(n_5759)
);

AOI22xp33_ASAP7_75t_L g5760 ( 
.A1(n_5400),
.A2(n_4410),
.B1(n_4356),
.B2(n_4541),
.Y(n_5760)
);

OR2x2_ASAP7_75t_L g5761 ( 
.A(n_4932),
.B(n_4538),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5123),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_5123),
.Y(n_5763)
);

NAND2xp5_ASAP7_75t_L g5764 ( 
.A(n_4908),
.B(n_4328),
.Y(n_5764)
);

CKINVDCx5p33_ASAP7_75t_R g5765 ( 
.A(n_4862),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_4972),
.Y(n_5766)
);

AOI22xp33_ASAP7_75t_L g5767 ( 
.A1(n_5270),
.A2(n_4356),
.B1(n_4541),
.B2(n_4596),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_4979),
.Y(n_5768)
);

INVx2_ASAP7_75t_L g5769 ( 
.A(n_5123),
.Y(n_5769)
);

INVx4_ASAP7_75t_L g5770 ( 
.A(n_4836),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_4979),
.Y(n_5771)
);

CKINVDCx5p33_ASAP7_75t_R g5772 ( 
.A(n_4958),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_4982),
.Y(n_5773)
);

INVx2_ASAP7_75t_L g5774 ( 
.A(n_5143),
.Y(n_5774)
);

HB1xp67_ASAP7_75t_L g5775 ( 
.A(n_5142),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5143),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_5143),
.Y(n_5777)
);

HB1xp67_ASAP7_75t_L g5778 ( 
.A(n_5142),
.Y(n_5778)
);

OAI21x1_ASAP7_75t_L g5779 ( 
.A1(n_5007),
.A2(n_4470),
.B(n_4594),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_4982),
.Y(n_5780)
);

BUFx2_ASAP7_75t_L g5781 ( 
.A(n_5403),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_4987),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_4987),
.Y(n_5783)
);

INVx3_ASAP7_75t_L g5784 ( 
.A(n_5101),
.Y(n_5784)
);

NAND2xp5_ASAP7_75t_L g5785 ( 
.A(n_5326),
.B(n_4401),
.Y(n_5785)
);

AO21x2_ASAP7_75t_L g5786 ( 
.A1(n_4990),
.A2(n_4301),
.B(n_4294),
.Y(n_5786)
);

INVx2_ASAP7_75t_L g5787 ( 
.A(n_5146),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_5146),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5146),
.Y(n_5789)
);

AND2x4_ASAP7_75t_L g5790 ( 
.A(n_5152),
.B(n_4297),
.Y(n_5790)
);

AOI21x1_ASAP7_75t_L g5791 ( 
.A1(n_4990),
.A2(n_4529),
.B(n_4377),
.Y(n_5791)
);

OAI21x1_ASAP7_75t_SL g5792 ( 
.A1(n_5257),
.A2(n_4631),
.B(n_4627),
.Y(n_5792)
);

INVx1_ASAP7_75t_SL g5793 ( 
.A(n_5390),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_5147),
.Y(n_5794)
);

OR2x2_ASAP7_75t_L g5795 ( 
.A(n_4998),
.B(n_5351),
.Y(n_5795)
);

AO21x2_ASAP7_75t_L g5796 ( 
.A1(n_4990),
.A2(n_4301),
.B(n_4294),
.Y(n_5796)
);

AOI22xp33_ASAP7_75t_L g5797 ( 
.A1(n_5192),
.A2(n_4356),
.B1(n_4541),
.B2(n_4596),
.Y(n_5797)
);

AO21x2_ASAP7_75t_L g5798 ( 
.A1(n_4991),
.A2(n_4301),
.B(n_4294),
.Y(n_5798)
);

INVx2_ASAP7_75t_L g5799 ( 
.A(n_5147),
.Y(n_5799)
);

OAI21x1_ASAP7_75t_L g5800 ( 
.A1(n_4886),
.A2(n_4513),
.B(n_4668),
.Y(n_5800)
);

INVx3_ASAP7_75t_L g5801 ( 
.A(n_5101),
.Y(n_5801)
);

OR2x2_ASAP7_75t_L g5802 ( 
.A(n_5367),
.B(n_4538),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5083),
.B(n_4379),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_4989),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_4989),
.Y(n_5805)
);

INVx2_ASAP7_75t_L g5806 ( 
.A(n_5147),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_4994),
.Y(n_5807)
);

INVx3_ASAP7_75t_L g5808 ( 
.A(n_5101),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_4994),
.Y(n_5809)
);

INVx2_ASAP7_75t_SL g5810 ( 
.A(n_5251),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_4996),
.Y(n_5811)
);

INVx2_ASAP7_75t_L g5812 ( 
.A(n_5162),
.Y(n_5812)
);

INVx2_ASAP7_75t_L g5813 ( 
.A(n_5162),
.Y(n_5813)
);

INVx3_ASAP7_75t_L g5814 ( 
.A(n_5403),
.Y(n_5814)
);

HB1xp67_ASAP7_75t_L g5815 ( 
.A(n_5326),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_4996),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5162),
.Y(n_5817)
);

AOI22xp33_ASAP7_75t_L g5818 ( 
.A1(n_5192),
.A2(n_4356),
.B1(n_4596),
.B2(n_4569),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_4999),
.Y(n_5819)
);

INVx2_ASAP7_75t_L g5820 ( 
.A(n_5163),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_4999),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5006),
.Y(n_5822)
);

INVx3_ASAP7_75t_L g5823 ( 
.A(n_5403),
.Y(n_5823)
);

OAI21x1_ASAP7_75t_L g5824 ( 
.A1(n_4886),
.A2(n_4513),
.B(n_4668),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5006),
.Y(n_5825)
);

BUFx3_ASAP7_75t_L g5826 ( 
.A(n_5179),
.Y(n_5826)
);

HB1xp67_ASAP7_75t_L g5827 ( 
.A(n_5345),
.Y(n_5827)
);

NOR2xp67_ASAP7_75t_L g5828 ( 
.A(n_5023),
.B(n_4670),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5008),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_4888),
.Y(n_5830)
);

BUFx2_ASAP7_75t_L g5831 ( 
.A(n_5403),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5008),
.Y(n_5832)
);

AND2x4_ASAP7_75t_L g5833 ( 
.A(n_5152),
.B(n_4297),
.Y(n_5833)
);

INVx3_ASAP7_75t_L g5834 ( 
.A(n_5414),
.Y(n_5834)
);

NOR2xp33_ASAP7_75t_L g5835 ( 
.A(n_4759),
.B(n_3682),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5163),
.Y(n_5836)
);

OR2x6_ASAP7_75t_L g5837 ( 
.A(n_4951),
.B(n_4487),
.Y(n_5837)
);

INVx4_ASAP7_75t_L g5838 ( 
.A(n_4836),
.Y(n_5838)
);

INVx3_ASAP7_75t_L g5839 ( 
.A(n_5414),
.Y(n_5839)
);

BUFx3_ASAP7_75t_L g5840 ( 
.A(n_4854),
.Y(n_5840)
);

OAI21x1_ASAP7_75t_L g5841 ( 
.A1(n_4886),
.A2(n_4513),
.B(n_4668),
.Y(n_5841)
);

INVx2_ASAP7_75t_L g5842 ( 
.A(n_5163),
.Y(n_5842)
);

NAND2xp5_ASAP7_75t_L g5843 ( 
.A(n_5345),
.B(n_4401),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5009),
.Y(n_5844)
);

OAI22xp33_ASAP7_75t_L g5845 ( 
.A1(n_4953),
.A2(n_4356),
.B1(n_4596),
.B2(n_4601),
.Y(n_5845)
);

NOR2x1_ASAP7_75t_R g5846 ( 
.A(n_4854),
.B(n_3732),
.Y(n_5846)
);

NAND2xp5_ASAP7_75t_L g5847 ( 
.A(n_4931),
.B(n_4463),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5009),
.Y(n_5848)
);

OA21x2_ASAP7_75t_L g5849 ( 
.A1(n_4882),
.A2(n_4299),
.B(n_4298),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5168),
.Y(n_5850)
);

NOR2xp33_ASAP7_75t_L g5851 ( 
.A(n_4759),
.B(n_3715),
.Y(n_5851)
);

NAND2x1p5_ASAP7_75t_L g5852 ( 
.A(n_5023),
.B(n_4297),
.Y(n_5852)
);

AOI22xp33_ASAP7_75t_L g5853 ( 
.A1(n_5064),
.A2(n_4596),
.B1(n_4558),
.B2(n_4569),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5010),
.Y(n_5854)
);

AOI22xp33_ASAP7_75t_SL g5855 ( 
.A1(n_5064),
.A2(n_4442),
.B1(n_4455),
.B2(n_4452),
.Y(n_5855)
);

BUFx8_ASAP7_75t_SL g5856 ( 
.A(n_4884),
.Y(n_5856)
);

OAI21x1_ASAP7_75t_L g5857 ( 
.A1(n_4919),
.A2(n_4685),
.B(n_4695),
.Y(n_5857)
);

AND2x2_ASAP7_75t_L g5858 ( 
.A(n_5083),
.B(n_4379),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5010),
.Y(n_5859)
);

AND2x2_ASAP7_75t_L g5860 ( 
.A(n_5187),
.B(n_4791),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_5014),
.Y(n_5861)
);

HB1xp67_ASAP7_75t_L g5862 ( 
.A(n_5384),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5014),
.Y(n_5863)
);

INVxp67_ASAP7_75t_L g5864 ( 
.A(n_5027),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5015),
.Y(n_5865)
);

AO21x2_ASAP7_75t_L g5866 ( 
.A1(n_4991),
.A2(n_4294),
.B(n_4532),
.Y(n_5866)
);

INVx2_ASAP7_75t_L g5867 ( 
.A(n_5168),
.Y(n_5867)
);

OR2x6_ASAP7_75t_L g5868 ( 
.A(n_5013),
.B(n_4487),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5015),
.Y(n_5869)
);

AND2x2_ASAP7_75t_L g5870 ( 
.A(n_5187),
.B(n_4442),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5016),
.Y(n_5871)
);

INVxp67_ASAP7_75t_L g5872 ( 
.A(n_5027),
.Y(n_5872)
);

NAND2xp5_ASAP7_75t_L g5873 ( 
.A(n_4935),
.B(n_4463),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5168),
.Y(n_5874)
);

INVx2_ASAP7_75t_L g5875 ( 
.A(n_5173),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5016),
.Y(n_5876)
);

OR2x2_ASAP7_75t_L g5877 ( 
.A(n_5389),
.B(n_4483),
.Y(n_5877)
);

OAI21x1_ASAP7_75t_L g5878 ( 
.A1(n_4919),
.A2(n_4685),
.B(n_4695),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5017),
.Y(n_5879)
);

INVx2_ASAP7_75t_L g5880 ( 
.A(n_5173),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_5017),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5018),
.Y(n_5882)
);

HB1xp67_ASAP7_75t_L g5883 ( 
.A(n_5407),
.Y(n_5883)
);

INVx3_ASAP7_75t_L g5884 ( 
.A(n_5414),
.Y(n_5884)
);

INVx2_ASAP7_75t_L g5885 ( 
.A(n_5173),
.Y(n_5885)
);

INVxp67_ASAP7_75t_L g5886 ( 
.A(n_5027),
.Y(n_5886)
);

HB1xp67_ASAP7_75t_L g5887 ( 
.A(n_5422),
.Y(n_5887)
);

HB1xp67_ASAP7_75t_L g5888 ( 
.A(n_5415),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5212),
.Y(n_5889)
);

INVx3_ASAP7_75t_SL g5890 ( 
.A(n_4901),
.Y(n_5890)
);

AOI21xp5_ASAP7_75t_L g5891 ( 
.A1(n_5200),
.A2(n_4440),
.B(n_4333),
.Y(n_5891)
);

OAI221xp5_ASAP7_75t_L g5892 ( 
.A1(n_5379),
.A2(n_4485),
.B1(n_4726),
.B2(n_4561),
.C(n_4568),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5018),
.Y(n_5893)
);

HB1xp67_ASAP7_75t_L g5894 ( 
.A(n_5415),
.Y(n_5894)
);

INVx2_ASAP7_75t_L g5895 ( 
.A(n_5212),
.Y(n_5895)
);

INVx2_ASAP7_75t_L g5896 ( 
.A(n_5212),
.Y(n_5896)
);

HB1xp67_ASAP7_75t_L g5897 ( 
.A(n_4762),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5022),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5022),
.Y(n_5899)
);

CKINVDCx5p33_ASAP7_75t_R g5900 ( 
.A(n_4889),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_4888),
.Y(n_5901)
);

NOR2xp33_ASAP7_75t_L g5902 ( 
.A(n_4814),
.B(n_3715),
.Y(n_5902)
);

INVx2_ASAP7_75t_L g5903 ( 
.A(n_4888),
.Y(n_5903)
);

INVx2_ASAP7_75t_SL g5904 ( 
.A(n_5251),
.Y(n_5904)
);

BUFx6f_ASAP7_75t_L g5905 ( 
.A(n_4854),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5026),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5026),
.Y(n_5907)
);

OR2x2_ASAP7_75t_L g5908 ( 
.A(n_5081),
.B(n_4483),
.Y(n_5908)
);

INVx2_ASAP7_75t_L g5909 ( 
.A(n_4915),
.Y(n_5909)
);

OR2x2_ASAP7_75t_L g5910 ( 
.A(n_5253),
.B(n_4507),
.Y(n_5910)
);

AO21x2_ASAP7_75t_L g5911 ( 
.A1(n_4991),
.A2(n_4532),
.B(n_4485),
.Y(n_5911)
);

INVx2_ASAP7_75t_L g5912 ( 
.A(n_4915),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_4915),
.Y(n_5913)
);

AND2x2_ASAP7_75t_L g5914 ( 
.A(n_4791),
.B(n_4442),
.Y(n_5914)
);

AO31x2_ASAP7_75t_L g5915 ( 
.A1(n_4954),
.A2(n_4681),
.A3(n_4701),
.B(n_4507),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_4808),
.B(n_4452),
.Y(n_5916)
);

INVx2_ASAP7_75t_SL g5917 ( 
.A(n_5251),
.Y(n_5917)
);

OAI21xp33_ASAP7_75t_SL g5918 ( 
.A1(n_5380),
.A2(n_4455),
.B(n_4452),
.Y(n_5918)
);

INVx2_ASAP7_75t_L g5919 ( 
.A(n_4926),
.Y(n_5919)
);

OAI21x1_ASAP7_75t_L g5920 ( 
.A1(n_4919),
.A2(n_4685),
.B(n_4695),
.Y(n_5920)
);

BUFx3_ASAP7_75t_L g5921 ( 
.A(n_4866),
.Y(n_5921)
);

AND2x2_ASAP7_75t_L g5922 ( 
.A(n_4808),
.B(n_4455),
.Y(n_5922)
);

NAND2x1p5_ASAP7_75t_L g5923 ( 
.A(n_5023),
.B(n_4393),
.Y(n_5923)
);

INVx3_ASAP7_75t_L g5924 ( 
.A(n_5414),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5042),
.Y(n_5925)
);

BUFx6f_ASAP7_75t_SL g5926 ( 
.A(n_4790),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5042),
.Y(n_5927)
);

AND2x2_ASAP7_75t_L g5928 ( 
.A(n_4949),
.B(n_4528),
.Y(n_5928)
);

NOR2xp33_ASAP7_75t_R g5929 ( 
.A(n_5080),
.B(n_3732),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5048),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5048),
.Y(n_5931)
);

INVx2_ASAP7_75t_L g5932 ( 
.A(n_4926),
.Y(n_5932)
);

HB1xp67_ASAP7_75t_L g5933 ( 
.A(n_4762),
.Y(n_5933)
);

INVx3_ASAP7_75t_L g5934 ( 
.A(n_5152),
.Y(n_5934)
);

INVx2_ASAP7_75t_L g5935 ( 
.A(n_4926),
.Y(n_5935)
);

OAI22xp5_ASAP7_75t_L g5936 ( 
.A1(n_5426),
.A2(n_4609),
.B1(n_4729),
.B2(n_4561),
.Y(n_5936)
);

INVx1_ASAP7_75t_L g5937 ( 
.A(n_5049),
.Y(n_5937)
);

AND2x2_ASAP7_75t_L g5938 ( 
.A(n_4949),
.B(n_4528),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_4946),
.Y(n_5939)
);

INVx2_ASAP7_75t_L g5940 ( 
.A(n_4946),
.Y(n_5940)
);

INVx1_ASAP7_75t_SL g5941 ( 
.A(n_5140),
.Y(n_5941)
);

INVx2_ASAP7_75t_L g5942 ( 
.A(n_4946),
.Y(n_5942)
);

INVx1_ASAP7_75t_SL g5943 ( 
.A(n_5218),
.Y(n_5943)
);

INVx2_ASAP7_75t_L g5944 ( 
.A(n_5216),
.Y(n_5944)
);

OAI21xp5_ASAP7_75t_L g5945 ( 
.A1(n_5215),
.A2(n_4440),
.B(n_4494),
.Y(n_5945)
);

AOI21x1_ASAP7_75t_L g5946 ( 
.A1(n_5011),
.A2(n_4377),
.B(n_4373),
.Y(n_5946)
);

NAND2xp5_ASAP7_75t_L g5947 ( 
.A(n_4952),
.B(n_4608),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_5216),
.Y(n_5948)
);

INVx1_ASAP7_75t_L g5949 ( 
.A(n_5049),
.Y(n_5949)
);

INVx2_ASAP7_75t_L g5950 ( 
.A(n_5216),
.Y(n_5950)
);

CKINVDCx5p33_ASAP7_75t_R g5951 ( 
.A(n_5012),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5053),
.Y(n_5952)
);

NAND2xp5_ASAP7_75t_L g5953 ( 
.A(n_4977),
.B(n_4608),
.Y(n_5953)
);

NAND2xp5_ASAP7_75t_L g5954 ( 
.A(n_4992),
.B(n_5005),
.Y(n_5954)
);

INVx1_ASAP7_75t_L g5955 ( 
.A(n_5053),
.Y(n_5955)
);

HB1xp67_ASAP7_75t_L g5956 ( 
.A(n_4768),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5061),
.Y(n_5957)
);

INVx2_ASAP7_75t_L g5958 ( 
.A(n_5237),
.Y(n_5958)
);

HB1xp67_ASAP7_75t_L g5959 ( 
.A(n_4768),
.Y(n_5959)
);

HB1xp67_ASAP7_75t_SL g5960 ( 
.A(n_5045),
.Y(n_5960)
);

AOI22xp33_ASAP7_75t_L g5961 ( 
.A1(n_5064),
.A2(n_4596),
.B1(n_4569),
.B2(n_4558),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5061),
.Y(n_5962)
);

INVx2_ASAP7_75t_L g5963 ( 
.A(n_5237),
.Y(n_5963)
);

OR2x6_ASAP7_75t_L g5964 ( 
.A(n_5013),
.B(n_4540),
.Y(n_5964)
);

AOI21x1_ASAP7_75t_L g5965 ( 
.A1(n_5011),
.A2(n_4377),
.B(n_4373),
.Y(n_5965)
);

NOR2xp33_ASAP7_75t_L g5966 ( 
.A(n_4814),
.B(n_4852),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5067),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5067),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5086),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5086),
.Y(n_5970)
);

HB1xp67_ASAP7_75t_L g5971 ( 
.A(n_4771),
.Y(n_5971)
);

INVx1_ASAP7_75t_L g5972 ( 
.A(n_5088),
.Y(n_5972)
);

HB1xp67_ASAP7_75t_L g5973 ( 
.A(n_4771),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5237),
.Y(n_5974)
);

AND2x2_ASAP7_75t_L g5975 ( 
.A(n_4950),
.B(n_4528),
.Y(n_5975)
);

INVx2_ASAP7_75t_L g5976 ( 
.A(n_5239),
.Y(n_5976)
);

BUFx3_ASAP7_75t_L g5977 ( 
.A(n_4866),
.Y(n_5977)
);

OAI21xp5_ASAP7_75t_L g5978 ( 
.A1(n_4947),
.A2(n_4494),
.B(n_4527),
.Y(n_5978)
);

BUFx6f_ASAP7_75t_L g5979 ( 
.A(n_4866),
.Y(n_5979)
);

AND2x2_ASAP7_75t_L g5980 ( 
.A(n_4950),
.B(n_5241),
.Y(n_5980)
);

INVx2_ASAP7_75t_L g5981 ( 
.A(n_5239),
.Y(n_5981)
);

INVx2_ASAP7_75t_L g5982 ( 
.A(n_5239),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5088),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5091),
.Y(n_5984)
);

INVx6_ASAP7_75t_L g5985 ( 
.A(n_4872),
.Y(n_5985)
);

BUFx2_ASAP7_75t_SL g5986 ( 
.A(n_5071),
.Y(n_5986)
);

OAI22xp5_ASAP7_75t_L g5987 ( 
.A1(n_4947),
.A2(n_4499),
.B1(n_4660),
.B2(n_4552),
.Y(n_5987)
);

CKINVDCx5p33_ASAP7_75t_R g5988 ( 
.A(n_5012),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5091),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5092),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5092),
.Y(n_5991)
);

INVx1_ASAP7_75t_L g5992 ( 
.A(n_5102),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5102),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5241),
.B(n_4558),
.Y(n_5994)
);

INVx3_ASAP7_75t_L g5995 ( 
.A(n_5152),
.Y(n_5995)
);

INVxp67_ASAP7_75t_L g5996 ( 
.A(n_5027),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5105),
.Y(n_5997)
);

OR2x2_ASAP7_75t_L g5998 ( 
.A(n_5269),
.B(n_4512),
.Y(n_5998)
);

INVxp33_ASAP7_75t_SL g5999 ( 
.A(n_5189),
.Y(n_5999)
);

INVx2_ASAP7_75t_L g6000 ( 
.A(n_5249),
.Y(n_6000)
);

AOI22xp33_ASAP7_75t_L g6001 ( 
.A1(n_5285),
.A2(n_4611),
.B1(n_4649),
.B2(n_4633),
.Y(n_6001)
);

BUFx12f_ASAP7_75t_L g6002 ( 
.A(n_4867),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5105),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5106),
.Y(n_6004)
);

INVx1_ASAP7_75t_L g6005 ( 
.A(n_5106),
.Y(n_6005)
);

OAI21x1_ASAP7_75t_L g6006 ( 
.A1(n_4937),
.A2(n_4941),
.B(n_4882),
.Y(n_6006)
);

HB1xp67_ASAP7_75t_L g6007 ( 
.A(n_4773),
.Y(n_6007)
);

AOI21x1_ASAP7_75t_L g6008 ( 
.A1(n_5011),
.A2(n_4390),
.B(n_4373),
.Y(n_6008)
);

OA21x2_ASAP7_75t_L g6009 ( 
.A1(n_4856),
.A2(n_4299),
.B(n_4298),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5108),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5108),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5249),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5110),
.Y(n_6013)
);

NOR2xp33_ASAP7_75t_L g6014 ( 
.A(n_4814),
.B(n_3715),
.Y(n_6014)
);

HB1xp67_ASAP7_75t_L g6015 ( 
.A(n_4773),
.Y(n_6015)
);

INVx2_ASAP7_75t_L g6016 ( 
.A(n_5249),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5110),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5111),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5111),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5252),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5113),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5113),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5119),
.Y(n_6023)
);

AND2x2_ASAP7_75t_L g6024 ( 
.A(n_5265),
.B(n_4611),
.Y(n_6024)
);

AND2x4_ASAP7_75t_L g6025 ( 
.A(n_5023),
.B(n_4393),
.Y(n_6025)
);

AND2x2_ASAP7_75t_L g6026 ( 
.A(n_5265),
.B(n_4611),
.Y(n_6026)
);

AND2x4_ASAP7_75t_L g6027 ( 
.A(n_5236),
.B(n_4393),
.Y(n_6027)
);

AND2x4_ASAP7_75t_L g6028 ( 
.A(n_5236),
.B(n_4406),
.Y(n_6028)
);

AND2x2_ASAP7_75t_L g6029 ( 
.A(n_5391),
.B(n_4571),
.Y(n_6029)
);

HB1xp67_ASAP7_75t_L g6030 ( 
.A(n_5119),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5120),
.Y(n_6031)
);

HB1xp67_ASAP7_75t_L g6032 ( 
.A(n_5120),
.Y(n_6032)
);

AND2x4_ASAP7_75t_L g6033 ( 
.A(n_5236),
.B(n_4406),
.Y(n_6033)
);

NAND2xp5_ASAP7_75t_L g6034 ( 
.A(n_5019),
.B(n_4734),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5122),
.Y(n_6035)
);

INVx4_ASAP7_75t_SL g6036 ( 
.A(n_5250),
.Y(n_6036)
);

AO21x2_ASAP7_75t_L g6037 ( 
.A1(n_5029),
.A2(n_4532),
.B(n_4618),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_5252),
.Y(n_6038)
);

INVx2_ASAP7_75t_L g6039 ( 
.A(n_5252),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5122),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5391),
.B(n_4571),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5309),
.B(n_4571),
.Y(n_6042)
);

AO21x2_ASAP7_75t_L g6043 ( 
.A1(n_5029),
.A2(n_4532),
.B(n_4618),
.Y(n_6043)
);

BUFx6f_ASAP7_75t_L g6044 ( 
.A(n_4867),
.Y(n_6044)
);

HB1xp67_ASAP7_75t_L g6045 ( 
.A(n_5129),
.Y(n_6045)
);

AND2x6_ASAP7_75t_L g6046 ( 
.A(n_5223),
.B(n_4499),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5129),
.Y(n_6047)
);

INVx3_ASAP7_75t_L g6048 ( 
.A(n_5321),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5273),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5130),
.Y(n_6050)
);

AND2x2_ASAP7_75t_L g6051 ( 
.A(n_5309),
.B(n_4571),
.Y(n_6051)
);

INVx2_ASAP7_75t_L g6052 ( 
.A(n_5273),
.Y(n_6052)
);

INVx3_ASAP7_75t_L g6053 ( 
.A(n_5321),
.Y(n_6053)
);

OAI21x1_ASAP7_75t_L g6054 ( 
.A1(n_4937),
.A2(n_4599),
.B(n_4468),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5130),
.Y(n_6055)
);

OAI21xp5_ASAP7_75t_L g6056 ( 
.A1(n_5118),
.A2(n_4527),
.B(n_4670),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5131),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5131),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_5132),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5132),
.Y(n_6060)
);

NOR2x1_ASAP7_75t_SL g6061 ( 
.A(n_5155),
.B(n_4641),
.Y(n_6061)
);

BUFx3_ASAP7_75t_L g6062 ( 
.A(n_4867),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5133),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5133),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5135),
.Y(n_6065)
);

AOI22xp33_ASAP7_75t_SL g6066 ( 
.A1(n_5371),
.A2(n_4633),
.B1(n_4649),
.B2(n_4499),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5135),
.Y(n_6067)
);

INVx2_ASAP7_75t_SL g6068 ( 
.A(n_5307),
.Y(n_6068)
);

BUFx3_ASAP7_75t_L g6069 ( 
.A(n_4872),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5273),
.Y(n_6070)
);

INVx4_ASAP7_75t_L g6071 ( 
.A(n_4835),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5136),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5136),
.Y(n_6073)
);

OAI21xp5_ASAP7_75t_L g6074 ( 
.A1(n_4811),
.A2(n_4333),
.B(n_4316),
.Y(n_6074)
);

OAI21x1_ASAP7_75t_L g6075 ( 
.A1(n_4937),
.A2(n_4599),
.B(n_4468),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5137),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_4764),
.B(n_4586),
.Y(n_6077)
);

BUFx6f_ASAP7_75t_L g6078 ( 
.A(n_4835),
.Y(n_6078)
);

HB1xp67_ASAP7_75t_L g6079 ( 
.A(n_5750),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_5432),
.Y(n_6080)
);

OA21x2_ASAP7_75t_L g6081 ( 
.A1(n_5539),
.A2(n_5041),
.B(n_5040),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_5432),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5434),
.Y(n_6083)
);

INVx3_ASAP7_75t_L g6084 ( 
.A(n_5558),
.Y(n_6084)
);

AO21x2_ASAP7_75t_L g6085 ( 
.A1(n_5700),
.A2(n_5047),
.B(n_4954),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_5453),
.B(n_5070),
.Y(n_6086)
);

AO21x2_ASAP7_75t_L g6087 ( 
.A1(n_5475),
.A2(n_5047),
.B(n_5032),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5946),
.Y(n_6088)
);

OR2x2_ASAP7_75t_L g6089 ( 
.A(n_5546),
.B(n_5409),
.Y(n_6089)
);

OR2x2_ASAP7_75t_L g6090 ( 
.A(n_5546),
.B(n_5409),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5434),
.Y(n_6091)
);

INVx2_ASAP7_75t_L g6092 ( 
.A(n_5946),
.Y(n_6092)
);

OAI21x1_ASAP7_75t_L g6093 ( 
.A1(n_5551),
.A2(n_5405),
.B(n_5344),
.Y(n_6093)
);

OR2x6_ASAP7_75t_L g6094 ( 
.A(n_5759),
.B(n_5248),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5436),
.Y(n_6095)
);

HB1xp67_ASAP7_75t_L g6096 ( 
.A(n_5752),
.Y(n_6096)
);

HB1xp67_ASAP7_75t_L g6097 ( 
.A(n_5775),
.Y(n_6097)
);

AND2x2_ASAP7_75t_L g6098 ( 
.A(n_5679),
.B(n_4764),
.Y(n_6098)
);

INVx2_ASAP7_75t_L g6099 ( 
.A(n_5965),
.Y(n_6099)
);

OR2x2_ASAP7_75t_L g6100 ( 
.A(n_5910),
.B(n_5374),
.Y(n_6100)
);

INVx2_ASAP7_75t_L g6101 ( 
.A(n_5965),
.Y(n_6101)
);

INVx5_ASAP7_75t_SL g6102 ( 
.A(n_5533),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_5436),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5448),
.Y(n_6104)
);

AND2x2_ASAP7_75t_L g6105 ( 
.A(n_5679),
.B(n_4833),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_5448),
.Y(n_6106)
);

OAI21xp5_ASAP7_75t_L g6107 ( 
.A1(n_6056),
.A2(n_4811),
.B(n_4816),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_5452),
.Y(n_6108)
);

NAND2xp5_ASAP7_75t_L g6109 ( 
.A(n_5592),
.B(n_5030),
.Y(n_6109)
);

AND2x4_ASAP7_75t_L g6110 ( 
.A(n_5447),
.B(n_4792),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5452),
.Y(n_6111)
);

INVx2_ASAP7_75t_L g6112 ( 
.A(n_6008),
.Y(n_6112)
);

NAND2xp5_ASAP7_75t_L g6113 ( 
.A(n_5642),
.B(n_5073),
.Y(n_6113)
);

INVx2_ASAP7_75t_L g6114 ( 
.A(n_6008),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_5711),
.B(n_4833),
.Y(n_6115)
);

BUFx6f_ASAP7_75t_L g6116 ( 
.A(n_5586),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5581),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5455),
.Y(n_6118)
);

INVx2_ASAP7_75t_SL g6119 ( 
.A(n_5435),
.Y(n_6119)
);

NOR2x1_ASAP7_75t_SL g6120 ( 
.A(n_5759),
.B(n_5155),
.Y(n_6120)
);

AND2x2_ASAP7_75t_L g6121 ( 
.A(n_5711),
.B(n_4921),
.Y(n_6121)
);

INVx2_ASAP7_75t_L g6122 ( 
.A(n_5581),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5455),
.Y(n_6123)
);

OAI21xp5_ASAP7_75t_L g6124 ( 
.A1(n_5978),
.A2(n_4816),
.B(n_5201),
.Y(n_6124)
);

NOR2xp33_ASAP7_75t_L g6125 ( 
.A(n_5595),
.B(n_4814),
.Y(n_6125)
);

AND2x2_ASAP7_75t_L g6126 ( 
.A(n_5524),
.B(n_4921),
.Y(n_6126)
);

INVx1_ASAP7_75t_SL g6127 ( 
.A(n_5549),
.Y(n_6127)
);

NOR2xp33_ASAP7_75t_L g6128 ( 
.A(n_5595),
.B(n_5951),
.Y(n_6128)
);

INVx2_ASAP7_75t_SL g6129 ( 
.A(n_5435),
.Y(n_6129)
);

OR2x2_ASAP7_75t_L g6130 ( 
.A(n_5910),
.B(n_5998),
.Y(n_6130)
);

AO21x2_ASAP7_75t_L g6131 ( 
.A1(n_5828),
.A2(n_5894),
.B(n_5888),
.Y(n_6131)
);

AND2x2_ASAP7_75t_L g6132 ( 
.A(n_5524),
.B(n_4964),
.Y(n_6132)
);

INVx2_ASAP7_75t_L g6133 ( 
.A(n_5583),
.Y(n_6133)
);

BUFx6f_ASAP7_75t_L g6134 ( 
.A(n_5586),
.Y(n_6134)
);

INVx2_ASAP7_75t_SL g6135 ( 
.A(n_5435),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_5464),
.Y(n_6136)
);

AND2x2_ASAP7_75t_L g6137 ( 
.A(n_5435),
.B(n_4964),
.Y(n_6137)
);

AND2x2_ASAP7_75t_L g6138 ( 
.A(n_5449),
.B(n_4857),
.Y(n_6138)
);

BUFx3_ASAP7_75t_L g6139 ( 
.A(n_5826),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_5583),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5464),
.Y(n_6141)
);

INVx2_ASAP7_75t_L g6142 ( 
.A(n_5588),
.Y(n_6142)
);

AND2x4_ASAP7_75t_L g6143 ( 
.A(n_5447),
.B(n_4792),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_5449),
.B(n_4857),
.Y(n_6144)
);

OAI21x1_ASAP7_75t_L g6145 ( 
.A1(n_5551),
.A2(n_5405),
.B(n_5344),
.Y(n_6145)
);

NAND2xp5_ASAP7_75t_L g6146 ( 
.A(n_5561),
.B(n_5073),
.Y(n_6146)
);

INVx2_ASAP7_75t_SL g6147 ( 
.A(n_5449),
.Y(n_6147)
);

OR2x2_ASAP7_75t_L g6148 ( 
.A(n_5998),
.B(n_5408),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_5468),
.Y(n_6149)
);

CKINVDCx5p33_ASAP7_75t_R g6150 ( 
.A(n_5856),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_5468),
.Y(n_6151)
);

HB1xp67_ASAP7_75t_L g6152 ( 
.A(n_5778),
.Y(n_6152)
);

INVx2_ASAP7_75t_L g6153 ( 
.A(n_5588),
.Y(n_6153)
);

BUFx6f_ASAP7_75t_L g6154 ( 
.A(n_5598),
.Y(n_6154)
);

HB1xp67_ASAP7_75t_L g6155 ( 
.A(n_5815),
.Y(n_6155)
);

BUFx3_ASAP7_75t_L g6156 ( 
.A(n_5826),
.Y(n_6156)
);

INVx3_ASAP7_75t_L g6157 ( 
.A(n_5558),
.Y(n_6157)
);

OR2x2_ASAP7_75t_L g6158 ( 
.A(n_5908),
.B(n_5623),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_5469),
.Y(n_6159)
);

INVxp67_ASAP7_75t_L g6160 ( 
.A(n_5960),
.Y(n_6160)
);

INVx1_ASAP7_75t_L g6161 ( 
.A(n_5469),
.Y(n_6161)
);

OAI221xp5_ASAP7_75t_L g6162 ( 
.A1(n_6001),
.A2(n_5327),
.B1(n_5377),
.B2(n_5000),
.C(n_4902),
.Y(n_6162)
);

AND2x2_ASAP7_75t_L g6163 ( 
.A(n_5449),
.B(n_4857),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5470),
.Y(n_6164)
);

NAND2xp5_ASAP7_75t_L g6165 ( 
.A(n_5579),
.B(n_5073),
.Y(n_6165)
);

AO21x2_ASAP7_75t_L g6166 ( 
.A1(n_5828),
.A2(n_5032),
.B(n_5029),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5470),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5478),
.Y(n_6168)
);

INVx2_ASAP7_75t_L g6169 ( 
.A(n_5589),
.Y(n_6169)
);

HB1xp67_ASAP7_75t_L g6170 ( 
.A(n_5827),
.Y(n_6170)
);

AOI21x1_ASAP7_75t_L g6171 ( 
.A1(n_5568),
.A2(n_5075),
.B(n_5025),
.Y(n_6171)
);

INVx2_ASAP7_75t_L g6172 ( 
.A(n_5589),
.Y(n_6172)
);

HB1xp67_ASAP7_75t_L g6173 ( 
.A(n_5641),
.Y(n_6173)
);

INVx2_ASAP7_75t_L g6174 ( 
.A(n_5599),
.Y(n_6174)
);

INVx2_ASAP7_75t_L g6175 ( 
.A(n_5599),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_5459),
.B(n_4857),
.Y(n_6176)
);

HB1xp67_ASAP7_75t_L g6177 ( 
.A(n_5649),
.Y(n_6177)
);

INVx2_ASAP7_75t_L g6178 ( 
.A(n_5605),
.Y(n_6178)
);

AND2x2_ASAP7_75t_L g6179 ( 
.A(n_5459),
.B(n_4997),
.Y(n_6179)
);

INVx2_ASAP7_75t_SL g6180 ( 
.A(n_5459),
.Y(n_6180)
);

AO21x2_ASAP7_75t_L g6181 ( 
.A1(n_5651),
.A2(n_5039),
.B(n_5032),
.Y(n_6181)
);

INVx2_ASAP7_75t_L g6182 ( 
.A(n_5605),
.Y(n_6182)
);

AND2x4_ASAP7_75t_L g6183 ( 
.A(n_5447),
.B(n_4792),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5478),
.Y(n_6184)
);

AND2x2_ASAP7_75t_L g6185 ( 
.A(n_5459),
.B(n_4997),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5480),
.Y(n_6186)
);

OR2x6_ASAP7_75t_L g6187 ( 
.A(n_5985),
.B(n_5248),
.Y(n_6187)
);

INVx3_ASAP7_75t_L g6188 ( 
.A(n_5447),
.Y(n_6188)
);

NOR2xp33_ASAP7_75t_L g6189 ( 
.A(n_5988),
.B(n_5670),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5480),
.Y(n_6190)
);

INVx2_ASAP7_75t_SL g6191 ( 
.A(n_5465),
.Y(n_6191)
);

AO31x2_ASAP7_75t_L g6192 ( 
.A1(n_5727),
.A2(n_5257),
.A3(n_5039),
.B(n_5248),
.Y(n_6192)
);

INVx2_ASAP7_75t_L g6193 ( 
.A(n_5609),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_5609),
.Y(n_6194)
);

INVx2_ASAP7_75t_L g6195 ( 
.A(n_5611),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5487),
.Y(n_6196)
);

OR2x2_ASAP7_75t_L g6197 ( 
.A(n_5908),
.B(n_5427),
.Y(n_6197)
);

INVx2_ASAP7_75t_SL g6198 ( 
.A(n_5465),
.Y(n_6198)
);

OR2x6_ASAP7_75t_L g6199 ( 
.A(n_5985),
.B(n_5248),
.Y(n_6199)
);

INVx3_ASAP7_75t_L g6200 ( 
.A(n_5615),
.Y(n_6200)
);

NOR2xp33_ASAP7_75t_L g6201 ( 
.A(n_5598),
.B(n_6002),
.Y(n_6201)
);

BUFx6f_ASAP7_75t_L g6202 ( 
.A(n_6002),
.Y(n_6202)
);

AO21x2_ASAP7_75t_L g6203 ( 
.A1(n_5651),
.A2(n_5039),
.B(n_5040),
.Y(n_6203)
);

OA21x2_ASAP7_75t_L g6204 ( 
.A1(n_5718),
.A2(n_5041),
.B(n_5040),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_5487),
.Y(n_6205)
);

AND2x2_ASAP7_75t_L g6206 ( 
.A(n_5465),
.B(n_5003),
.Y(n_6206)
);

AND2x2_ASAP7_75t_L g6207 ( 
.A(n_5465),
.B(n_5003),
.Y(n_6207)
);

AND2x2_ASAP7_75t_L g6208 ( 
.A(n_5476),
.B(n_5271),
.Y(n_6208)
);

NOR2xp33_ASAP7_75t_L g6209 ( 
.A(n_5770),
.B(n_4852),
.Y(n_6209)
);

OA21x2_ASAP7_75t_L g6210 ( 
.A1(n_5718),
.A2(n_5051),
.B(n_5041),
.Y(n_6210)
);

INVx3_ASAP7_75t_L g6211 ( 
.A(n_5615),
.Y(n_6211)
);

AND2x4_ASAP7_75t_L g6212 ( 
.A(n_5615),
.B(n_4792),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_5489),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_5611),
.Y(n_6214)
);

OA21x2_ASAP7_75t_L g6215 ( 
.A1(n_5718),
.A2(n_5055),
.B(n_5051),
.Y(n_6215)
);

INVx2_ASAP7_75t_L g6216 ( 
.A(n_5612),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_5476),
.B(n_5498),
.Y(n_6217)
);

INVx3_ASAP7_75t_L g6218 ( 
.A(n_5615),
.Y(n_6218)
);

INVx3_ASAP7_75t_SL g6219 ( 
.A(n_5572),
.Y(n_6219)
);

OA21x2_ASAP7_75t_L g6220 ( 
.A1(n_5723),
.A2(n_5055),
.B(n_5051),
.Y(n_6220)
);

INVx1_ASAP7_75t_L g6221 ( 
.A(n_5489),
.Y(n_6221)
);

OR2x6_ASAP7_75t_L g6222 ( 
.A(n_5985),
.B(n_5365),
.Y(n_6222)
);

INVx2_ASAP7_75t_SL g6223 ( 
.A(n_5476),
.Y(n_6223)
);

AND2x2_ASAP7_75t_L g6224 ( 
.A(n_5476),
.B(n_5271),
.Y(n_6224)
);

OAI21x1_ASAP7_75t_L g6225 ( 
.A1(n_5466),
.A2(n_4881),
.B(n_4767),
.Y(n_6225)
);

OAI21x1_ASAP7_75t_L g6226 ( 
.A1(n_5466),
.A2(n_4881),
.B(n_4767),
.Y(n_6226)
);

INVx2_ASAP7_75t_L g6227 ( 
.A(n_5612),
.Y(n_6227)
);

OAI21x1_ASAP7_75t_L g6228 ( 
.A1(n_5482),
.A2(n_4881),
.B(n_4767),
.Y(n_6228)
);

INVx3_ASAP7_75t_L g6229 ( 
.A(n_5695),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5490),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5490),
.Y(n_6231)
);

AO21x2_ASAP7_75t_L g6232 ( 
.A1(n_5651),
.A2(n_5055),
.B(n_5372),
.Y(n_6232)
);

HB1xp67_ASAP7_75t_L g6233 ( 
.A(n_5662),
.Y(n_6233)
);

AOI22xp33_ASAP7_75t_SL g6234 ( 
.A1(n_5892),
.A2(n_5548),
.B1(n_5945),
.B2(n_5987),
.Y(n_6234)
);

AO21x2_ASAP7_75t_L g6235 ( 
.A1(n_5510),
.A2(n_4957),
.B(n_4956),
.Y(n_6235)
);

OA21x2_ASAP7_75t_L g6236 ( 
.A1(n_5723),
.A2(n_4957),
.B(n_4956),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_5493),
.Y(n_6237)
);

BUFx6f_ASAP7_75t_L g6238 ( 
.A(n_5826),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_5493),
.Y(n_6239)
);

OA21x2_ASAP7_75t_L g6240 ( 
.A1(n_5723),
.A2(n_4957),
.B(n_4956),
.Y(n_6240)
);

OAI21xp5_ASAP7_75t_L g6241 ( 
.A1(n_5530),
.A2(n_5201),
.B(n_4878),
.Y(n_6241)
);

NAND2xp5_ASAP7_75t_L g6242 ( 
.A(n_5441),
.B(n_5082),
.Y(n_6242)
);

OAI21x1_ASAP7_75t_L g6243 ( 
.A1(n_5482),
.A2(n_5161),
.B(n_5138),
.Y(n_6243)
);

OR2x6_ASAP7_75t_L g6244 ( 
.A(n_5985),
.B(n_5365),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5499),
.Y(n_6245)
);

AND2x2_ASAP7_75t_L g6246 ( 
.A(n_5498),
.B(n_5280),
.Y(n_6246)
);

AO21x2_ASAP7_75t_L g6247 ( 
.A1(n_5510),
.A2(n_4959),
.B(n_5306),
.Y(n_6247)
);

OA21x2_ASAP7_75t_L g6248 ( 
.A1(n_5725),
.A2(n_4959),
.B(n_5138),
.Y(n_6248)
);

OA21x2_ASAP7_75t_L g6249 ( 
.A1(n_5725),
.A2(n_5731),
.B(n_5627),
.Y(n_6249)
);

OR2x2_ASAP7_75t_L g6250 ( 
.A(n_5623),
.B(n_4512),
.Y(n_6250)
);

CKINVDCx5p33_ASAP7_75t_R g6251 ( 
.A(n_5986),
.Y(n_6251)
);

INVx2_ASAP7_75t_L g6252 ( 
.A(n_5614),
.Y(n_6252)
);

INVx2_ASAP7_75t_L g6253 ( 
.A(n_5614),
.Y(n_6253)
);

INVx1_ASAP7_75t_L g6254 ( 
.A(n_5499),
.Y(n_6254)
);

INVx2_ASAP7_75t_L g6255 ( 
.A(n_5617),
.Y(n_6255)
);

AO21x2_ASAP7_75t_L g6256 ( 
.A1(n_5510),
.A2(n_4959),
.B(n_5306),
.Y(n_6256)
);

OR2x2_ASAP7_75t_L g6257 ( 
.A(n_5619),
.B(n_4522),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5504),
.Y(n_6258)
);

INVx2_ASAP7_75t_L g6259 ( 
.A(n_5617),
.Y(n_6259)
);

AND2x2_ASAP7_75t_L g6260 ( 
.A(n_5498),
.B(n_5280),
.Y(n_6260)
);

INVxp67_ASAP7_75t_L g6261 ( 
.A(n_5986),
.Y(n_6261)
);

INVx2_ASAP7_75t_SL g6262 ( 
.A(n_5498),
.Y(n_6262)
);

BUFx4f_ASAP7_75t_SL g6263 ( 
.A(n_5890),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_5504),
.Y(n_6264)
);

AND2x2_ASAP7_75t_L g6265 ( 
.A(n_5503),
.B(n_5371),
.Y(n_6265)
);

INVxp67_ASAP7_75t_L g6266 ( 
.A(n_5542),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_5507),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_5507),
.Y(n_6268)
);

OR2x2_ASAP7_75t_L g6269 ( 
.A(n_5619),
.B(n_4522),
.Y(n_6269)
);

OR2x2_ASAP7_75t_L g6270 ( 
.A(n_5877),
.B(n_4531),
.Y(n_6270)
);

AND2x2_ASAP7_75t_L g6271 ( 
.A(n_5503),
.B(n_5035),
.Y(n_6271)
);

HB1xp67_ASAP7_75t_L g6272 ( 
.A(n_5667),
.Y(n_6272)
);

OR2x2_ASAP7_75t_L g6273 ( 
.A(n_5877),
.B(n_5631),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5509),
.Y(n_6274)
);

AO21x2_ASAP7_75t_L g6275 ( 
.A1(n_5505),
.A2(n_5322),
.B(n_5306),
.Y(n_6275)
);

INVx2_ASAP7_75t_L g6276 ( 
.A(n_5628),
.Y(n_6276)
);

NOR2x1_ASAP7_75t_SL g6277 ( 
.A(n_5837),
.B(n_5394),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_5509),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_5628),
.Y(n_6279)
);

OR2x2_ASAP7_75t_L g6280 ( 
.A(n_5631),
.B(n_4531),
.Y(n_6280)
);

INVx2_ASAP7_75t_L g6281 ( 
.A(n_5629),
.Y(n_6281)
);

NAND2xp5_ASAP7_75t_L g6282 ( 
.A(n_5947),
.B(n_5082),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_5513),
.Y(n_6283)
);

BUFx2_ASAP7_75t_L g6284 ( 
.A(n_5695),
.Y(n_6284)
);

INVx2_ASAP7_75t_L g6285 ( 
.A(n_5629),
.Y(n_6285)
);

OR2x2_ASAP7_75t_L g6286 ( 
.A(n_5682),
.B(n_5528),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_5503),
.B(n_5035),
.Y(n_6287)
);

BUFx2_ASAP7_75t_L g6288 ( 
.A(n_5695),
.Y(n_6288)
);

OAI221xp5_ASAP7_75t_SL g6289 ( 
.A1(n_5618),
.A2(n_5377),
.B1(n_5420),
.B2(n_5429),
.C(n_5327),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_5633),
.Y(n_6290)
);

OAI21x1_ASAP7_75t_L g6291 ( 
.A1(n_5483),
.A2(n_5167),
.B(n_5161),
.Y(n_6291)
);

BUFx3_ASAP7_75t_L g6292 ( 
.A(n_5890),
.Y(n_6292)
);

AND2x2_ASAP7_75t_L g6293 ( 
.A(n_5503),
.B(n_5037),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_5513),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_5519),
.B(n_5037),
.Y(n_6295)
);

HB1xp67_ASAP7_75t_L g6296 ( 
.A(n_5672),
.Y(n_6296)
);

NAND2xp5_ASAP7_75t_L g6297 ( 
.A(n_5953),
.B(n_5082),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_5519),
.B(n_5934),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_5514),
.Y(n_6299)
);

HB1xp67_ASAP7_75t_L g6300 ( 
.A(n_5684),
.Y(n_6300)
);

NOR2xp33_ASAP7_75t_L g6301 ( 
.A(n_5770),
.B(n_4852),
.Y(n_6301)
);

NOR2xp33_ASAP7_75t_L g6302 ( 
.A(n_5770),
.B(n_4852),
.Y(n_6302)
);

AND2x4_ASAP7_75t_L g6303 ( 
.A(n_5695),
.B(n_4792),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5514),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_5633),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_5516),
.Y(n_6306)
);

INVx2_ASAP7_75t_L g6307 ( 
.A(n_5645),
.Y(n_6307)
);

AND2x4_ASAP7_75t_L g6308 ( 
.A(n_5698),
.B(n_5236),
.Y(n_6308)
);

AO21x2_ASAP7_75t_L g6309 ( 
.A1(n_5505),
.A2(n_5332),
.B(n_5322),
.Y(n_6309)
);

AO21x2_ASAP7_75t_L g6310 ( 
.A1(n_5505),
.A2(n_5332),
.B(n_5322),
.Y(n_6310)
);

HB1xp67_ASAP7_75t_L g6311 ( 
.A(n_5696),
.Y(n_6311)
);

OR2x2_ASAP7_75t_L g6312 ( 
.A(n_5682),
.B(n_4734),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5516),
.Y(n_6313)
);

NAND2xp5_ASAP7_75t_L g6314 ( 
.A(n_5686),
.B(n_5283),
.Y(n_6314)
);

BUFx6f_ASAP7_75t_L g6315 ( 
.A(n_5533),
.Y(n_6315)
);

AO21x2_ASAP7_75t_L g6316 ( 
.A1(n_5735),
.A2(n_5332),
.B(n_4963),
.Y(n_6316)
);

AND2x2_ASAP7_75t_L g6317 ( 
.A(n_5519),
.B(n_5112),
.Y(n_6317)
);

NAND3xp33_ASAP7_75t_SL g6318 ( 
.A(n_5727),
.B(n_5127),
.C(n_5341),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_5519),
.B(n_5112),
.Y(n_6319)
);

AO21x2_ASAP7_75t_L g6320 ( 
.A1(n_5735),
.A2(n_6074),
.B(n_6043),
.Y(n_6320)
);

AND2x4_ASAP7_75t_L g6321 ( 
.A(n_5698),
.B(n_5236),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5521),
.Y(n_6322)
);

OR2x2_ASAP7_75t_L g6323 ( 
.A(n_5528),
.B(n_4744),
.Y(n_6323)
);

INVx2_ASAP7_75t_L g6324 ( 
.A(n_5645),
.Y(n_6324)
);

INVx3_ASAP7_75t_L g6325 ( 
.A(n_5698),
.Y(n_6325)
);

OR2x6_ASAP7_75t_L g6326 ( 
.A(n_6071),
.B(n_5365),
.Y(n_6326)
);

INVx2_ASAP7_75t_SL g6327 ( 
.A(n_6078),
.Y(n_6327)
);

OR2x2_ASAP7_75t_L g6328 ( 
.A(n_5795),
.B(n_4744),
.Y(n_6328)
);

INVxp67_ASAP7_75t_SL g6329 ( 
.A(n_5708),
.Y(n_6329)
);

AND2x2_ASAP7_75t_L g6330 ( 
.A(n_5934),
.B(n_5156),
.Y(n_6330)
);

OR2x6_ASAP7_75t_L g6331 ( 
.A(n_6071),
.B(n_5385),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_5646),
.Y(n_6332)
);

OAI21xp5_ASAP7_75t_L g6333 ( 
.A1(n_5891),
.A2(n_4766),
.B(n_4860),
.Y(n_6333)
);

BUFx3_ASAP7_75t_L g6334 ( 
.A(n_5890),
.Y(n_6334)
);

BUFx2_ASAP7_75t_L g6335 ( 
.A(n_5698),
.Y(n_6335)
);

AO21x2_ASAP7_75t_L g6336 ( 
.A1(n_5735),
.A2(n_4963),
.B(n_4962),
.Y(n_6336)
);

AO21x2_ASAP7_75t_L g6337 ( 
.A1(n_6037),
.A2(n_4963),
.B(n_4962),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_5646),
.Y(n_6338)
);

AND2x2_ASAP7_75t_L g6339 ( 
.A(n_5934),
.B(n_5156),
.Y(n_6339)
);

NAND2xp5_ASAP7_75t_L g6340 ( 
.A(n_5721),
.B(n_5283),
.Y(n_6340)
);

OA21x2_ASAP7_75t_L g6341 ( 
.A1(n_5725),
.A2(n_5177),
.B(n_5167),
.Y(n_6341)
);

OA21x2_ASAP7_75t_L g6342 ( 
.A1(n_5731),
.A2(n_5238),
.B(n_5177),
.Y(n_6342)
);

NAND2xp5_ASAP7_75t_L g6343 ( 
.A(n_5454),
.B(n_5317),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_5521),
.Y(n_6344)
);

OA21x2_ASAP7_75t_L g6345 ( 
.A1(n_5731),
.A2(n_5240),
.B(n_5238),
.Y(n_6345)
);

INVx2_ASAP7_75t_L g6346 ( 
.A(n_5647),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_5522),
.Y(n_6347)
);

INVx8_ASAP7_75t_L g6348 ( 
.A(n_5479),
.Y(n_6348)
);

OR2x6_ASAP7_75t_L g6349 ( 
.A(n_6071),
.B(n_5385),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_5647),
.Y(n_6350)
);

AO21x2_ASAP7_75t_L g6351 ( 
.A1(n_6037),
.A2(n_4975),
.B(n_4962),
.Y(n_6351)
);

OA21x2_ASAP7_75t_L g6352 ( 
.A1(n_5627),
.A2(n_5245),
.B(n_5240),
.Y(n_6352)
);

AO21x2_ASAP7_75t_L g6353 ( 
.A1(n_6037),
.A2(n_4981),
.B(n_4975),
.Y(n_6353)
);

INVx1_ASAP7_75t_L g6354 ( 
.A(n_5522),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_5523),
.Y(n_6355)
);

OR2x2_ASAP7_75t_L g6356 ( 
.A(n_5795),
.B(n_4433),
.Y(n_6356)
);

INVx3_ASAP7_75t_L g6357 ( 
.A(n_5496),
.Y(n_6357)
);

OR2x6_ASAP7_75t_L g6358 ( 
.A(n_6071),
.B(n_5385),
.Y(n_6358)
);

OA21x2_ASAP7_75t_L g6359 ( 
.A1(n_5644),
.A2(n_5299),
.B(n_5245),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_5523),
.Y(n_6360)
);

AND2x2_ASAP7_75t_L g6361 ( 
.A(n_5934),
.B(n_5165),
.Y(n_6361)
);

AND2x2_ASAP7_75t_L g6362 ( 
.A(n_5995),
.B(n_5165),
.Y(n_6362)
);

NAND2xp5_ASAP7_75t_L g6363 ( 
.A(n_5472),
.B(n_5317),
.Y(n_6363)
);

AND2x4_ASAP7_75t_L g6364 ( 
.A(n_5630),
.B(n_5236),
.Y(n_6364)
);

INVx2_ASAP7_75t_L g6365 ( 
.A(n_5737),
.Y(n_6365)
);

OR2x6_ASAP7_75t_L g6366 ( 
.A(n_6078),
.B(n_5301),
.Y(n_6366)
);

INVx2_ASAP7_75t_L g6367 ( 
.A(n_5737),
.Y(n_6367)
);

AO21x2_ASAP7_75t_L g6368 ( 
.A1(n_6043),
.A2(n_5792),
.B(n_5911),
.Y(n_6368)
);

BUFx3_ASAP7_75t_L g6369 ( 
.A(n_5467),
.Y(n_6369)
);

CKINVDCx20_ASAP7_75t_R g6370 ( 
.A(n_5681),
.Y(n_6370)
);

AND2x2_ASAP7_75t_L g6371 ( 
.A(n_5995),
.B(n_5172),
.Y(n_6371)
);

AOI22xp33_ASAP7_75t_L g6372 ( 
.A1(n_5855),
.A2(n_4804),
.B1(n_4799),
.B2(n_5054),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_5995),
.B(n_5172),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_5532),
.Y(n_6374)
);

AO21x2_ASAP7_75t_L g6375 ( 
.A1(n_6043),
.A2(n_4981),
.B(n_4975),
.Y(n_6375)
);

CKINVDCx5p33_ASAP7_75t_R g6376 ( 
.A(n_5501),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_5532),
.Y(n_6377)
);

INVx3_ASAP7_75t_L g6378 ( 
.A(n_5496),
.Y(n_6378)
);

AO21x2_ASAP7_75t_L g6379 ( 
.A1(n_5792),
.A2(n_5911),
.B(n_5584),
.Y(n_6379)
);

AND2x4_ASAP7_75t_L g6380 ( 
.A(n_5630),
.B(n_5235),
.Y(n_6380)
);

HB1xp67_ASAP7_75t_L g6381 ( 
.A(n_5596),
.Y(n_6381)
);

INVx3_ASAP7_75t_L g6382 ( 
.A(n_5496),
.Y(n_6382)
);

BUFx6f_ASAP7_75t_L g6383 ( 
.A(n_5533),
.Y(n_6383)
);

INVx2_ASAP7_75t_SL g6384 ( 
.A(n_6078),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_5535),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_5535),
.Y(n_6386)
);

CKINVDCx5p33_ASAP7_75t_R g6387 ( 
.A(n_5929),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5536),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_5536),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_5995),
.B(n_5320),
.Y(n_6390)
);

INVx2_ASAP7_75t_L g6391 ( 
.A(n_5744),
.Y(n_6391)
);

NAND2xp5_ASAP7_75t_L g6392 ( 
.A(n_5484),
.B(n_5320),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_5537),
.Y(n_6393)
);

OR2x6_ASAP7_75t_L g6394 ( 
.A(n_6078),
.B(n_5301),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_5537),
.Y(n_6395)
);

AND2x2_ASAP7_75t_L g6396 ( 
.A(n_5438),
.B(n_5357),
.Y(n_6396)
);

INVx2_ASAP7_75t_L g6397 ( 
.A(n_5744),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_5438),
.B(n_5357),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_5538),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_5538),
.Y(n_6400)
);

OA21x2_ASAP7_75t_L g6401 ( 
.A1(n_5644),
.A2(n_5355),
.B(n_5299),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_5540),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_5747),
.Y(n_6403)
);

INVx2_ASAP7_75t_L g6404 ( 
.A(n_5747),
.Y(n_6404)
);

AO21x2_ASAP7_75t_L g6405 ( 
.A1(n_5911),
.A2(n_4984),
.B(n_4981),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_5540),
.Y(n_6406)
);

AND2x4_ASAP7_75t_L g6407 ( 
.A(n_5630),
.B(n_5235),
.Y(n_6407)
);

AOI21x1_ASAP7_75t_L g6408 ( 
.A1(n_5568),
.A2(n_5075),
.B(n_5025),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_5544),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5544),
.Y(n_6410)
);

INVx3_ASAP7_75t_L g6411 ( 
.A(n_5674),
.Y(n_6411)
);

INVx2_ASAP7_75t_L g6412 ( 
.A(n_5749),
.Y(n_6412)
);

HB1xp67_ASAP7_75t_L g6413 ( 
.A(n_5613),
.Y(n_6413)
);

INVx2_ASAP7_75t_L g6414 ( 
.A(n_5749),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_5553),
.Y(n_6415)
);

HB1xp67_ASAP7_75t_L g6416 ( 
.A(n_5637),
.Y(n_6416)
);

INVx1_ASAP7_75t_SL g6417 ( 
.A(n_5517),
.Y(n_6417)
);

AND2x2_ASAP7_75t_L g6418 ( 
.A(n_5630),
.B(n_5099),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_5553),
.Y(n_6419)
);

AND2x2_ASAP7_75t_L g6420 ( 
.A(n_5678),
.B(n_5099),
.Y(n_6420)
);

NOR2x1_ASAP7_75t_R g6421 ( 
.A(n_5654),
.B(n_4884),
.Y(n_6421)
);

OAI21x1_ASAP7_75t_L g6422 ( 
.A1(n_5483),
.A2(n_5355),
.B(n_4837),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_5751),
.Y(n_6423)
);

INVx2_ASAP7_75t_L g6424 ( 
.A(n_5751),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_5554),
.Y(n_6425)
);

NAND2x1_ASAP7_75t_L g6426 ( 
.A(n_5678),
.B(n_5702),
.Y(n_6426)
);

NAND2xp5_ASAP7_75t_L g6427 ( 
.A(n_5690),
.B(n_4784),
.Y(n_6427)
);

BUFx6f_ASAP7_75t_L g6428 ( 
.A(n_5533),
.Y(n_6428)
);

AND2x2_ASAP7_75t_L g6429 ( 
.A(n_5678),
.B(n_5134),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_5554),
.Y(n_6430)
);

AO21x2_ASAP7_75t_L g6431 ( 
.A1(n_5584),
.A2(n_4988),
.B(n_4984),
.Y(n_6431)
);

INVx2_ASAP7_75t_L g6432 ( 
.A(n_5757),
.Y(n_6432)
);

OAI22xp33_ASAP7_75t_L g6433 ( 
.A1(n_5699),
.A2(n_4883),
.B1(n_4810),
.B2(n_5087),
.Y(n_6433)
);

INVx2_ASAP7_75t_SL g6434 ( 
.A(n_6078),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_5557),
.Y(n_6435)
);

AOI21x1_ASAP7_75t_L g6436 ( 
.A1(n_5573),
.A2(n_5157),
.B(n_5134),
.Y(n_6436)
);

AND2x2_ASAP7_75t_L g6437 ( 
.A(n_5678),
.B(n_5157),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_5557),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_5560),
.Y(n_6439)
);

NAND3xp33_ASAP7_75t_L g6440 ( 
.A(n_5699),
.B(n_4933),
.C(n_4930),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_5757),
.Y(n_6441)
);

INVx2_ASAP7_75t_L g6442 ( 
.A(n_5758),
.Y(n_6442)
);

NAND2xp5_ASAP7_75t_L g6443 ( 
.A(n_5764),
.B(n_4784),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_5560),
.Y(n_6444)
);

NAND2xp5_ASAP7_75t_L g6445 ( 
.A(n_5864),
.B(n_4633),
.Y(n_6445)
);

AO21x2_ASAP7_75t_L g6446 ( 
.A1(n_5584),
.A2(n_4988),
.B(n_4984),
.Y(n_6446)
);

AO21x2_ASAP7_75t_L g6447 ( 
.A1(n_5866),
.A2(n_4988),
.B(n_4818),
.Y(n_6447)
);

AND2x4_ASAP7_75t_L g6448 ( 
.A(n_5702),
.B(n_5235),
.Y(n_6448)
);

INVx3_ASAP7_75t_L g6449 ( 
.A(n_5674),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_5566),
.Y(n_6450)
);

INVx2_ASAP7_75t_L g6451 ( 
.A(n_5758),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_5566),
.Y(n_6452)
);

INVx2_ASAP7_75t_L g6453 ( 
.A(n_5762),
.Y(n_6453)
);

NAND2xp5_ASAP7_75t_L g6454 ( 
.A(n_5872),
.B(n_4649),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_5702),
.B(n_5185),
.Y(n_6455)
);

AND2x2_ASAP7_75t_L g6456 ( 
.A(n_5702),
.B(n_5185),
.Y(n_6456)
);

OR2x6_ASAP7_75t_L g6457 ( 
.A(n_5479),
.B(n_5301),
.Y(n_6457)
);

AND2x2_ASAP7_75t_L g6458 ( 
.A(n_5710),
.B(n_5186),
.Y(n_6458)
);

INVx2_ASAP7_75t_L g6459 ( 
.A(n_5762),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_5575),
.Y(n_6460)
);

INVx1_ASAP7_75t_L g6461 ( 
.A(n_5575),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_5580),
.Y(n_6462)
);

NAND2x1p5_ASAP7_75t_L g6463 ( 
.A(n_5527),
.B(n_5197),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_5580),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_5710),
.B(n_5186),
.Y(n_6465)
);

OR2x2_ASAP7_75t_L g6466 ( 
.A(n_5862),
.B(n_4433),
.Y(n_6466)
);

BUFx2_ASAP7_75t_L g6467 ( 
.A(n_5573),
.Y(n_6467)
);

AND2x2_ASAP7_75t_L g6468 ( 
.A(n_5710),
.B(n_5225),
.Y(n_6468)
);

INVx2_ASAP7_75t_L g6469 ( 
.A(n_5763),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_5582),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_5763),
.Y(n_6471)
);

INVx2_ASAP7_75t_L g6472 ( 
.A(n_5769),
.Y(n_6472)
);

NOR2x1_ASAP7_75t_L g6473 ( 
.A(n_5840),
.B(n_5250),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_L g6474 ( 
.A(n_5886),
.B(n_5033),
.Y(n_6474)
);

HB1xp67_ASAP7_75t_L g6475 ( 
.A(n_5437),
.Y(n_6475)
);

BUFx12f_ASAP7_75t_L g6476 ( 
.A(n_5533),
.Y(n_6476)
);

BUFx2_ASAP7_75t_L g6477 ( 
.A(n_5621),
.Y(n_6477)
);

INVx2_ASAP7_75t_L g6478 ( 
.A(n_5769),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_5582),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5591),
.Y(n_6480)
);

INVx3_ASAP7_75t_L g6481 ( 
.A(n_5674),
.Y(n_6481)
);

BUFx2_ASAP7_75t_L g6482 ( 
.A(n_5621),
.Y(n_6482)
);

HB1xp67_ASAP7_75t_L g6483 ( 
.A(n_5444),
.Y(n_6483)
);

BUFx2_ASAP7_75t_L g6484 ( 
.A(n_5625),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_5591),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_5774),
.Y(n_6486)
);

BUFx12f_ASAP7_75t_L g6487 ( 
.A(n_5563),
.Y(n_6487)
);

INVx3_ASAP7_75t_SL g6488 ( 
.A(n_6036),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_5774),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_5594),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_5594),
.Y(n_6491)
);

NOR2xp33_ASAP7_75t_SL g6492 ( 
.A(n_5846),
.B(n_5189),
.Y(n_6492)
);

OA21x2_ASAP7_75t_L g6493 ( 
.A1(n_5730),
.A2(n_4973),
.B(n_4903),
.Y(n_6493)
);

BUFx2_ASAP7_75t_L g6494 ( 
.A(n_5625),
.Y(n_6494)
);

AO21x2_ASAP7_75t_L g6495 ( 
.A1(n_5866),
.A2(n_4818),
.B(n_4817),
.Y(n_6495)
);

INVx3_ASAP7_75t_L g6496 ( 
.A(n_5852),
.Y(n_6496)
);

INVx2_ASAP7_75t_L g6497 ( 
.A(n_5776),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_5597),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_5597),
.Y(n_6499)
);

INVx2_ASAP7_75t_L g6500 ( 
.A(n_5776),
.Y(n_6500)
);

BUFx2_ASAP7_75t_L g6501 ( 
.A(n_5675),
.Y(n_6501)
);

BUFx2_ASAP7_75t_SL g6502 ( 
.A(n_5926),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_5600),
.Y(n_6503)
);

INVx2_ASAP7_75t_L g6504 ( 
.A(n_5777),
.Y(n_6504)
);

AO21x2_ASAP7_75t_L g6505 ( 
.A1(n_5866),
.A2(n_4818),
.B(n_4817),
.Y(n_6505)
);

INVx2_ASAP7_75t_L g6506 ( 
.A(n_5777),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_5787),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_5600),
.Y(n_6508)
);

AO21x2_ASAP7_75t_L g6509 ( 
.A1(n_6061),
.A2(n_4820),
.B(n_4817),
.Y(n_6509)
);

AO21x2_ASAP7_75t_L g6510 ( 
.A1(n_6061),
.A2(n_4820),
.B(n_4966),
.Y(n_6510)
);

AO21x1_ASAP7_75t_SL g6511 ( 
.A1(n_5534),
.A2(n_4912),
.B(n_4810),
.Y(n_6511)
);

INVx2_ASAP7_75t_SL g6512 ( 
.A(n_5479),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_5602),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_5602),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_5604),
.Y(n_6515)
);

INVx2_ASAP7_75t_L g6516 ( 
.A(n_5787),
.Y(n_6516)
);

INVx2_ASAP7_75t_L g6517 ( 
.A(n_5788),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_5604),
.Y(n_6518)
);

INVxp67_ASAP7_75t_L g6519 ( 
.A(n_5481),
.Y(n_6519)
);

HB1xp67_ASAP7_75t_L g6520 ( 
.A(n_5883),
.Y(n_6520)
);

AOI22xp33_ASAP7_75t_L g6521 ( 
.A1(n_5818),
.A2(n_4923),
.B1(n_4805),
.B2(n_4934),
.Y(n_6521)
);

AND2x4_ASAP7_75t_SL g6522 ( 
.A(n_5710),
.B(n_4901),
.Y(n_6522)
);

INVxp67_ASAP7_75t_SL g6523 ( 
.A(n_5996),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_5606),
.Y(n_6524)
);

INVx2_ASAP7_75t_L g6525 ( 
.A(n_5788),
.Y(n_6525)
);

INVx5_ASAP7_75t_L g6526 ( 
.A(n_5563),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_5606),
.Y(n_6527)
);

INVx2_ASAP7_75t_L g6528 ( 
.A(n_5789),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_5789),
.Y(n_6529)
);

AND2x2_ASAP7_75t_L g6530 ( 
.A(n_5728),
.B(n_5225),
.Y(n_6530)
);

HB1xp67_ASAP7_75t_L g6531 ( 
.A(n_5887),
.Y(n_6531)
);

NOR2xp33_ASAP7_75t_L g6532 ( 
.A(n_5770),
.B(n_5838),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_5607),
.Y(n_6533)
);

AOI22xp33_ASAP7_75t_L g6534 ( 
.A1(n_5936),
.A2(n_5145),
.B1(n_4770),
.B2(n_4859),
.Y(n_6534)
);

INVx2_ASAP7_75t_L g6535 ( 
.A(n_5794),
.Y(n_6535)
);

AND2x2_ASAP7_75t_L g6536 ( 
.A(n_5728),
.B(n_5234),
.Y(n_6536)
);

HB1xp67_ASAP7_75t_L g6537 ( 
.A(n_5675),
.Y(n_6537)
);

AND2x2_ASAP7_75t_L g6538 ( 
.A(n_5728),
.B(n_5234),
.Y(n_6538)
);

AND2x2_ASAP7_75t_L g6539 ( 
.A(n_5728),
.B(n_5247),
.Y(n_6539)
);

BUFx2_ASAP7_75t_L g6540 ( 
.A(n_5677),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_5607),
.Y(n_6541)
);

AND2x2_ASAP7_75t_L g6542 ( 
.A(n_5525),
.B(n_5247),
.Y(n_6542)
);

INVx8_ASAP7_75t_L g6543 ( 
.A(n_5479),
.Y(n_6543)
);

BUFx6f_ASAP7_75t_L g6544 ( 
.A(n_5563),
.Y(n_6544)
);

BUFx2_ASAP7_75t_L g6545 ( 
.A(n_5677),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_5610),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_5610),
.Y(n_6547)
);

HB1xp67_ASAP7_75t_L g6548 ( 
.A(n_5897),
.Y(n_6548)
);

OA21x2_ASAP7_75t_L g6549 ( 
.A1(n_5730),
.A2(n_4973),
.B(n_4903),
.Y(n_6549)
);

AO21x2_ASAP7_75t_L g6550 ( 
.A1(n_5786),
.A2(n_4820),
.B(n_4966),
.Y(n_6550)
);

OAI21xp5_ASAP7_75t_L g6551 ( 
.A1(n_5918),
.A2(n_5395),
.B(n_4969),
.Y(n_6551)
);

OR2x2_ASAP7_75t_L g6552 ( 
.A(n_5802),
.B(n_4433),
.Y(n_6552)
);

INVxp67_ASAP7_75t_SL g6553 ( 
.A(n_5705),
.Y(n_6553)
);

INVx2_ASAP7_75t_L g6554 ( 
.A(n_5794),
.Y(n_6554)
);

BUFx6f_ASAP7_75t_L g6555 ( 
.A(n_5563),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_5616),
.Y(n_6556)
);

INVx2_ASAP7_75t_L g6557 ( 
.A(n_5799),
.Y(n_6557)
);

INVx2_ASAP7_75t_SL g6558 ( 
.A(n_5479),
.Y(n_6558)
);

HB1xp67_ASAP7_75t_L g6559 ( 
.A(n_5933),
.Y(n_6559)
);

OR2x2_ASAP7_75t_L g6560 ( 
.A(n_5802),
.B(n_4433),
.Y(n_6560)
);

INVxp67_ASAP7_75t_R g6561 ( 
.A(n_6036),
.Y(n_6561)
);

AO21x2_ASAP7_75t_L g6562 ( 
.A1(n_5786),
.A2(n_5084),
.B(n_4813),
.Y(n_6562)
);

INVx2_ASAP7_75t_L g6563 ( 
.A(n_5799),
.Y(n_6563)
);

NAND3xp33_ASAP7_75t_L g6564 ( 
.A(n_5534),
.B(n_5304),
.C(n_5303),
.Y(n_6564)
);

INVx2_ASAP7_75t_L g6565 ( 
.A(n_5806),
.Y(n_6565)
);

NOR2xp33_ASAP7_75t_L g6566 ( 
.A(n_5838),
.B(n_5999),
.Y(n_6566)
);

INVx2_ASAP7_75t_L g6567 ( 
.A(n_5806),
.Y(n_6567)
);

OA21x2_ASAP7_75t_L g6568 ( 
.A1(n_5626),
.A2(n_5068),
.B(n_4974),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_5616),
.Y(n_6569)
);

AND2x2_ASAP7_75t_L g6570 ( 
.A(n_5525),
.B(n_5279),
.Y(n_6570)
);

AO21x2_ASAP7_75t_L g6571 ( 
.A1(n_5786),
.A2(n_5084),
.B(n_4813),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_5632),
.Y(n_6572)
);

HB1xp67_ASAP7_75t_L g6573 ( 
.A(n_5956),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_5632),
.Y(n_6574)
);

NAND2xp5_ASAP7_75t_L g6575 ( 
.A(n_5954),
.B(n_5033),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_5639),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_5567),
.B(n_5570),
.Y(n_6577)
);

AND2x2_ASAP7_75t_L g6578 ( 
.A(n_5567),
.B(n_5279),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_5639),
.Y(n_6579)
);

AND2x2_ASAP7_75t_L g6580 ( 
.A(n_5570),
.B(n_5296),
.Y(n_6580)
);

INVx1_ASAP7_75t_L g6581 ( 
.A(n_5640),
.Y(n_6581)
);

NOR2xp33_ASAP7_75t_L g6582 ( 
.A(n_5838),
.B(n_5144),
.Y(n_6582)
);

INVx2_ASAP7_75t_SL g6583 ( 
.A(n_5814),
.Y(n_6583)
);

INVx1_ASAP7_75t_L g6584 ( 
.A(n_5640),
.Y(n_6584)
);

INVx2_ASAP7_75t_L g6585 ( 
.A(n_5812),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_5643),
.Y(n_6586)
);

NAND2xp5_ASAP7_75t_L g6587 ( 
.A(n_5634),
.B(n_5128),
.Y(n_6587)
);

OAI21xp5_ASAP7_75t_L g6588 ( 
.A1(n_5918),
.A2(n_4968),
.B(n_5258),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_5643),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_5648),
.Y(n_6590)
);

INVx1_ASAP7_75t_L g6591 ( 
.A(n_5648),
.Y(n_6591)
);

HB1xp67_ASAP7_75t_L g6592 ( 
.A(n_5959),
.Y(n_6592)
);

INVx2_ASAP7_75t_L g6593 ( 
.A(n_5812),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_5653),
.Y(n_6594)
);

OAI21xp5_ASAP7_75t_L g6595 ( 
.A1(n_5797),
.A2(n_5593),
.B(n_5853),
.Y(n_6595)
);

NAND2xp5_ASAP7_75t_L g6596 ( 
.A(n_5785),
.B(n_5128),
.Y(n_6596)
);

AO21x2_ASAP7_75t_L g6597 ( 
.A1(n_5796),
.A2(n_4813),
.B(n_4980),
.Y(n_6597)
);

AND2x2_ASAP7_75t_L g6598 ( 
.A(n_5585),
.B(n_5296),
.Y(n_6598)
);

AOI22xp33_ASAP7_75t_SL g6599 ( 
.A1(n_5668),
.A2(n_4828),
.B1(n_4795),
.B2(n_4796),
.Y(n_6599)
);

OAI21xp5_ASAP7_75t_L g6600 ( 
.A1(n_5961),
.A2(n_4912),
.B(n_4819),
.Y(n_6600)
);

OR2x6_ASAP7_75t_L g6601 ( 
.A(n_5837),
.B(n_5114),
.Y(n_6601)
);

HB1xp67_ASAP7_75t_L g6602 ( 
.A(n_5971),
.Y(n_6602)
);

BUFx2_ASAP7_75t_L g6603 ( 
.A(n_5781),
.Y(n_6603)
);

OR2x6_ASAP7_75t_L g6604 ( 
.A(n_5837),
.B(n_5114),
.Y(n_6604)
);

INVx1_ASAP7_75t_L g6605 ( 
.A(n_5653),
.Y(n_6605)
);

HB1xp67_ASAP7_75t_L g6606 ( 
.A(n_5973),
.Y(n_6606)
);

INVx2_ASAP7_75t_SL g6607 ( 
.A(n_5814),
.Y(n_6607)
);

NAND2xp5_ASAP7_75t_L g6608 ( 
.A(n_5843),
.B(n_5158),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_5655),
.Y(n_6609)
);

INVx2_ASAP7_75t_L g6610 ( 
.A(n_5813),
.Y(n_6610)
);

INVx2_ASAP7_75t_SL g6611 ( 
.A(n_5814),
.Y(n_6611)
);

AOI22xp33_ASAP7_75t_L g6612 ( 
.A1(n_5837),
.A2(n_5145),
.B1(n_4868),
.B2(n_5089),
.Y(n_6612)
);

INVx2_ASAP7_75t_L g6613 ( 
.A(n_5813),
.Y(n_6613)
);

INVxp67_ASAP7_75t_L g6614 ( 
.A(n_5511),
.Y(n_6614)
);

INVx2_ASAP7_75t_L g6615 ( 
.A(n_5817),
.Y(n_6615)
);

INVx2_ASAP7_75t_SL g6616 ( 
.A(n_5814),
.Y(n_6616)
);

NAND2xp5_ASAP7_75t_L g6617 ( 
.A(n_5456),
.B(n_5158),
.Y(n_6617)
);

AO21x2_ASAP7_75t_L g6618 ( 
.A1(n_5796),
.A2(n_4813),
.B(n_4980),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_5585),
.B(n_5587),
.Y(n_6619)
);

HB1xp67_ASAP7_75t_L g6620 ( 
.A(n_6007),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6467),
.Y(n_6621)
);

OAI322xp33_ASAP7_75t_L g6622 ( 
.A1(n_6089),
.A2(n_5518),
.A3(n_5451),
.B1(n_5526),
.B2(n_5506),
.C1(n_5845),
.C2(n_5761),
.Y(n_6622)
);

HB1xp67_ASAP7_75t_L g6623 ( 
.A(n_6467),
.Y(n_6623)
);

OR2x2_ASAP7_75t_SL g6624 ( 
.A(n_6318),
.B(n_5563),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6477),
.Y(n_6625)
);

INVx2_ASAP7_75t_L g6626 ( 
.A(n_6477),
.Y(n_6626)
);

NOR2x1_ASAP7_75t_L g6627 ( 
.A(n_6084),
.B(n_5840),
.Y(n_6627)
);

BUFx2_ASAP7_75t_L g6628 ( 
.A(n_6263),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6482),
.Y(n_6629)
);

AND2x2_ASAP7_75t_L g6630 ( 
.A(n_6522),
.B(n_6098),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6522),
.B(n_6036),
.Y(n_6631)
);

HB1xp67_ASAP7_75t_L g6632 ( 
.A(n_6482),
.Y(n_6632)
);

AND2x2_ASAP7_75t_L g6633 ( 
.A(n_6098),
.B(n_6036),
.Y(n_6633)
);

BUFx3_ASAP7_75t_L g6634 ( 
.A(n_6139),
.Y(n_6634)
);

INVx2_ASAP7_75t_SL g6635 ( 
.A(n_6139),
.Y(n_6635)
);

AND2x2_ASAP7_75t_L g6636 ( 
.A(n_6105),
.B(n_6036),
.Y(n_6636)
);

HB1xp67_ASAP7_75t_L g6637 ( 
.A(n_6484),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_6484),
.Y(n_6638)
);

AND2x2_ASAP7_75t_L g6639 ( 
.A(n_6105),
.B(n_5445),
.Y(n_6639)
);

INVx2_ASAP7_75t_L g6640 ( 
.A(n_6494),
.Y(n_6640)
);

AND2x4_ASAP7_75t_L g6641 ( 
.A(n_6094),
.B(n_5823),
.Y(n_6641)
);

AND2x4_ASAP7_75t_L g6642 ( 
.A(n_6094),
.B(n_5823),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6494),
.Y(n_6643)
);

NOR2x1_ASAP7_75t_SL g6644 ( 
.A(n_6511),
.B(n_5837),
.Y(n_6644)
);

INVx1_ASAP7_75t_L g6645 ( 
.A(n_6501),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6501),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6540),
.Y(n_6647)
);

BUFx2_ASAP7_75t_L g6648 ( 
.A(n_6292),
.Y(n_6648)
);

INVx2_ASAP7_75t_L g6649 ( 
.A(n_6540),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_6545),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_6545),
.Y(n_6651)
);

AND2x2_ASAP7_75t_L g6652 ( 
.A(n_6463),
.B(n_5445),
.Y(n_6652)
);

INVx2_ASAP7_75t_L g6653 ( 
.A(n_6603),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6080),
.Y(n_6654)
);

OR2x2_ASAP7_75t_L g6655 ( 
.A(n_6089),
.B(n_5873),
.Y(n_6655)
);

AOI222xp33_ASAP7_75t_L g6656 ( 
.A1(n_6595),
.A2(n_6241),
.B1(n_6440),
.B2(n_6124),
.C1(n_6333),
.C2(n_6564),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6603),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6082),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_6166),
.Y(n_6659)
);

NAND2xp5_ASAP7_75t_L g6660 ( 
.A(n_6109),
.B(n_5810),
.Y(n_6660)
);

INVx2_ASAP7_75t_L g6661 ( 
.A(n_6166),
.Y(n_6661)
);

HB1xp67_ASAP7_75t_L g6662 ( 
.A(n_6537),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6083),
.Y(n_6663)
);

AOI21x1_ASAP7_75t_L g6664 ( 
.A1(n_6171),
.A2(n_5831),
.B(n_5781),
.Y(n_6664)
);

AND2x2_ASAP7_75t_L g6665 ( 
.A(n_6115),
.B(n_6121),
.Y(n_6665)
);

HB1xp67_ASAP7_75t_L g6666 ( 
.A(n_6079),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_6166),
.Y(n_6667)
);

AOI22xp33_ASAP7_75t_L g6668 ( 
.A1(n_6234),
.A2(n_6107),
.B1(n_6599),
.B2(n_6433),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_6091),
.Y(n_6669)
);

INVx2_ASAP7_75t_SL g6670 ( 
.A(n_6156),
.Y(n_6670)
);

OR2x2_ASAP7_75t_L g6671 ( 
.A(n_6090),
.B(n_5847),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6095),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6368),
.Y(n_6673)
);

OR2x2_ASAP7_75t_L g6674 ( 
.A(n_6090),
.B(n_6282),
.Y(n_6674)
);

BUFx4f_ASAP7_75t_L g6675 ( 
.A(n_6202),
.Y(n_6675)
);

INVx2_ASAP7_75t_L g6676 ( 
.A(n_6368),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6103),
.Y(n_6677)
);

AND2x2_ASAP7_75t_L g6678 ( 
.A(n_6115),
.B(n_5473),
.Y(n_6678)
);

INVxp67_ASAP7_75t_L g6679 ( 
.A(n_6523),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_6121),
.B(n_5473),
.Y(n_6680)
);

OR2x2_ASAP7_75t_L g6681 ( 
.A(n_6297),
.B(n_5601),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_6104),
.Y(n_6682)
);

NAND2xp5_ASAP7_75t_L g6683 ( 
.A(n_6261),
.B(n_6266),
.Y(n_6683)
);

INVx2_ASAP7_75t_L g6684 ( 
.A(n_6368),
.Y(n_6684)
);

AND2x2_ASAP7_75t_L g6685 ( 
.A(n_6110),
.B(n_5500),
.Y(n_6685)
);

INVx2_ASAP7_75t_L g6686 ( 
.A(n_6232),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6106),
.Y(n_6687)
);

INVxp33_ASAP7_75t_SL g6688 ( 
.A(n_6251),
.Y(n_6688)
);

AND2x2_ASAP7_75t_L g6689 ( 
.A(n_6110),
.B(n_5500),
.Y(n_6689)
);

OR2x2_ASAP7_75t_L g6690 ( 
.A(n_6096),
.B(n_6034),
.Y(n_6690)
);

AND2x4_ASAP7_75t_L g6691 ( 
.A(n_6094),
.B(n_5823),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_6108),
.Y(n_6692)
);

HB1xp67_ASAP7_75t_L g6693 ( 
.A(n_6097),
.Y(n_6693)
);

INVxp67_ASAP7_75t_SL g6694 ( 
.A(n_6152),
.Y(n_6694)
);

NAND2xp5_ASAP7_75t_L g6695 ( 
.A(n_6519),
.B(n_5810),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6111),
.Y(n_6696)
);

HB1xp67_ASAP7_75t_L g6697 ( 
.A(n_6155),
.Y(n_6697)
);

NAND2xp5_ASAP7_75t_L g6698 ( 
.A(n_6614),
.B(n_5904),
.Y(n_6698)
);

INVx2_ASAP7_75t_L g6699 ( 
.A(n_6232),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6118),
.Y(n_6700)
);

AND2x2_ASAP7_75t_L g6701 ( 
.A(n_6110),
.B(n_5433),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_6123),
.Y(n_6702)
);

AND2x2_ASAP7_75t_L g6703 ( 
.A(n_6143),
.B(n_5433),
.Y(n_6703)
);

AND2x2_ASAP7_75t_L g6704 ( 
.A(n_6143),
.B(n_5440),
.Y(n_6704)
);

INVx2_ASAP7_75t_SL g6705 ( 
.A(n_6156),
.Y(n_6705)
);

AND2x2_ASAP7_75t_L g6706 ( 
.A(n_6143),
.B(n_5440),
.Y(n_6706)
);

INVx4_ASAP7_75t_L g6707 ( 
.A(n_6202),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6183),
.B(n_5442),
.Y(n_6708)
);

INVx2_ASAP7_75t_L g6709 ( 
.A(n_6232),
.Y(n_6709)
);

AND2x2_ASAP7_75t_L g6710 ( 
.A(n_6183),
.B(n_6212),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6183),
.B(n_5442),
.Y(n_6711)
);

AOI22xp33_ASAP7_75t_L g6712 ( 
.A1(n_6085),
.A2(n_5868),
.B1(n_5492),
.B2(n_5767),
.Y(n_6712)
);

INVx2_ASAP7_75t_L g6713 ( 
.A(n_6542),
.Y(n_6713)
);

OR2x2_ASAP7_75t_L g6714 ( 
.A(n_6170),
.B(n_5748),
.Y(n_6714)
);

INVx2_ASAP7_75t_L g6715 ( 
.A(n_6542),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6136),
.Y(n_6716)
);

AOI22xp33_ASAP7_75t_L g6717 ( 
.A1(n_6085),
.A2(n_5868),
.B1(n_5492),
.B2(n_5502),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6570),
.Y(n_6718)
);

OAI22xp5_ASAP7_75t_L g6719 ( 
.A1(n_6372),
.A2(n_6066),
.B1(n_5760),
.B2(n_5729),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6141),
.Y(n_6720)
);

AND2x4_ASAP7_75t_L g6721 ( 
.A(n_6094),
.B(n_6284),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_L g6722 ( 
.A(n_6381),
.B(n_5904),
.Y(n_6722)
);

INVx2_ASAP7_75t_L g6723 ( 
.A(n_6570),
.Y(n_6723)
);

INVx2_ASAP7_75t_L g6724 ( 
.A(n_6408),
.Y(n_6724)
);

AND2x4_ASAP7_75t_L g6725 ( 
.A(n_6284),
.B(n_5823),
.Y(n_6725)
);

AND2x2_ASAP7_75t_L g6726 ( 
.A(n_6212),
.B(n_5443),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6149),
.Y(n_6727)
);

HB1xp67_ASAP7_75t_L g6728 ( 
.A(n_6173),
.Y(n_6728)
);

BUFx2_ASAP7_75t_L g6729 ( 
.A(n_6292),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_6436),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_6151),
.Y(n_6731)
);

AND2x2_ASAP7_75t_L g6732 ( 
.A(n_6212),
.B(n_5443),
.Y(n_6732)
);

BUFx2_ASAP7_75t_L g6733 ( 
.A(n_6334),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_6578),
.Y(n_6734)
);

INVx2_ASAP7_75t_L g6735 ( 
.A(n_6578),
.Y(n_6735)
);

INVx3_ASAP7_75t_L g6736 ( 
.A(n_6238),
.Y(n_6736)
);

INVxp67_ASAP7_75t_SL g6737 ( 
.A(n_6177),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6159),
.Y(n_6738)
);

AND2x4_ASAP7_75t_SL g6739 ( 
.A(n_6222),
.B(n_4906),
.Y(n_6739)
);

BUFx3_ASAP7_75t_L g6740 ( 
.A(n_6251),
.Y(n_6740)
);

INVx2_ASAP7_75t_L g6741 ( 
.A(n_6580),
.Y(n_6741)
);

NAND2xp5_ASAP7_75t_L g6742 ( 
.A(n_6413),
.B(n_5917),
.Y(n_6742)
);

INVx1_ASAP7_75t_L g6743 ( 
.A(n_6161),
.Y(n_6743)
);

INVx1_ASAP7_75t_L g6744 ( 
.A(n_6164),
.Y(n_6744)
);

AND2x2_ASAP7_75t_L g6745 ( 
.A(n_6303),
.B(n_5457),
.Y(n_6745)
);

AND2x2_ASAP7_75t_L g6746 ( 
.A(n_6303),
.B(n_6126),
.Y(n_6746)
);

AND2x2_ASAP7_75t_L g6747 ( 
.A(n_6303),
.B(n_5457),
.Y(n_6747)
);

BUFx3_ASAP7_75t_L g6748 ( 
.A(n_6238),
.Y(n_6748)
);

INVx1_ASAP7_75t_SL g6749 ( 
.A(n_6127),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_6126),
.B(n_5529),
.Y(n_6750)
);

AND2x2_ASAP7_75t_L g6751 ( 
.A(n_6132),
.B(n_5529),
.Y(n_6751)
);

OR2x2_ASAP7_75t_L g6752 ( 
.A(n_6329),
.B(n_5656),
.Y(n_6752)
);

INVx2_ASAP7_75t_L g6753 ( 
.A(n_6580),
.Y(n_6753)
);

AND2x2_ASAP7_75t_L g6754 ( 
.A(n_6132),
.B(n_5569),
.Y(n_6754)
);

AND2x2_ASAP7_75t_L g6755 ( 
.A(n_6222),
.B(n_5569),
.Y(n_6755)
);

INVxp67_ASAP7_75t_SL g6756 ( 
.A(n_6233),
.Y(n_6756)
);

AOI33xp33_ASAP7_75t_L g6757 ( 
.A1(n_6534),
.A2(n_5941),
.A3(n_5943),
.B1(n_5754),
.B2(n_5343),
.B3(n_5361),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_6416),
.B(n_5917),
.Y(n_6758)
);

INVx1_ASAP7_75t_L g6759 ( 
.A(n_6167),
.Y(n_6759)
);

INVx1_ASAP7_75t_L g6760 ( 
.A(n_6168),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6184),
.Y(n_6761)
);

INVx2_ASAP7_75t_L g6762 ( 
.A(n_6598),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_6598),
.Y(n_6763)
);

AND2x2_ASAP7_75t_L g6764 ( 
.A(n_6222),
.B(n_6244),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6186),
.Y(n_6765)
);

AND2x2_ASAP7_75t_L g6766 ( 
.A(n_6222),
.B(n_5622),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6086),
.B(n_6068),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_6272),
.B(n_6068),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6244),
.B(n_5622),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6244),
.B(n_5652),
.Y(n_6770)
);

NAND2xp5_ASAP7_75t_L g6771 ( 
.A(n_6296),
.B(n_5556),
.Y(n_6771)
);

INVx3_ASAP7_75t_L g6772 ( 
.A(n_6238),
.Y(n_6772)
);

AND2x2_ASAP7_75t_L g6773 ( 
.A(n_6244),
.B(n_5652),
.Y(n_6773)
);

BUFx3_ASAP7_75t_L g6774 ( 
.A(n_6238),
.Y(n_6774)
);

BUFx3_ASAP7_75t_L g6775 ( 
.A(n_6219),
.Y(n_6775)
);

INVx3_ASAP7_75t_L g6776 ( 
.A(n_6308),
.Y(n_6776)
);

AND2x4_ASAP7_75t_SL g6777 ( 
.A(n_6084),
.B(n_6157),
.Y(n_6777)
);

OR2x2_ASAP7_75t_L g6778 ( 
.A(n_6300),
.B(n_5707),
.Y(n_6778)
);

INVx2_ASAP7_75t_L g6779 ( 
.A(n_6379),
.Y(n_6779)
);

HB1xp67_ASAP7_75t_L g6780 ( 
.A(n_6311),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_6190),
.Y(n_6781)
);

BUFx3_ASAP7_75t_L g6782 ( 
.A(n_6219),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6196),
.Y(n_6783)
);

NAND2xp5_ASAP7_75t_L g6784 ( 
.A(n_6475),
.B(n_5556),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6205),
.Y(n_6785)
);

AND2x4_ASAP7_75t_L g6786 ( 
.A(n_6288),
.B(n_5834),
.Y(n_6786)
);

BUFx2_ASAP7_75t_L g6787 ( 
.A(n_6334),
.Y(n_6787)
);

INVx2_ASAP7_75t_L g6788 ( 
.A(n_6379),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6213),
.Y(n_6789)
);

INVxp67_ASAP7_75t_L g6790 ( 
.A(n_6502),
.Y(n_6790)
);

AND2x2_ASAP7_75t_L g6791 ( 
.A(n_6084),
.B(n_5720),
.Y(n_6791)
);

OR2x2_ASAP7_75t_L g6792 ( 
.A(n_6100),
.B(n_5831),
.Y(n_6792)
);

INVx2_ASAP7_75t_L g6793 ( 
.A(n_6379),
.Y(n_6793)
);

INVx2_ASAP7_75t_L g6794 ( 
.A(n_6181),
.Y(n_6794)
);

AND2x2_ASAP7_75t_L g6795 ( 
.A(n_6463),
.B(n_5527),
.Y(n_6795)
);

INVx2_ASAP7_75t_L g6796 ( 
.A(n_6181),
.Y(n_6796)
);

BUFx3_ASAP7_75t_L g6797 ( 
.A(n_6150),
.Y(n_6797)
);

AND2x2_ASAP7_75t_L g6798 ( 
.A(n_6577),
.B(n_5527),
.Y(n_6798)
);

INVx2_ASAP7_75t_L g6799 ( 
.A(n_6181),
.Y(n_6799)
);

HB1xp67_ASAP7_75t_L g6800 ( 
.A(n_6483),
.Y(n_6800)
);

NAND2xp5_ASAP7_75t_L g6801 ( 
.A(n_6520),
.B(n_6531),
.Y(n_6801)
);

INVx2_ASAP7_75t_L g6802 ( 
.A(n_6119),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_6221),
.Y(n_6803)
);

OR2x2_ASAP7_75t_L g6804 ( 
.A(n_6100),
.B(n_5527),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_L g6805 ( 
.A(n_6327),
.B(n_5562),
.Y(n_6805)
);

NAND2xp5_ASAP7_75t_L g6806 ( 
.A(n_6327),
.B(n_5562),
.Y(n_6806)
);

AOI221xp5_ASAP7_75t_L g6807 ( 
.A1(n_6289),
.A2(n_5966),
.B1(n_5926),
.B2(n_4726),
.C(n_5905),
.Y(n_6807)
);

INVxp67_ASAP7_75t_L g6808 ( 
.A(n_6157),
.Y(n_6808)
);

BUFx2_ASAP7_75t_L g6809 ( 
.A(n_6157),
.Y(n_6809)
);

INVx2_ASAP7_75t_L g6810 ( 
.A(n_6119),
.Y(n_6810)
);

INVx3_ASAP7_75t_L g6811 ( 
.A(n_6308),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6230),
.Y(n_6812)
);

AND2x2_ASAP7_75t_L g6813 ( 
.A(n_6308),
.B(n_5720),
.Y(n_6813)
);

OR2x2_ASAP7_75t_L g6814 ( 
.A(n_6148),
.B(n_5915),
.Y(n_6814)
);

AND2x2_ASAP7_75t_L g6815 ( 
.A(n_6321),
.B(n_5467),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_6321),
.B(n_5467),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6321),
.B(n_5502),
.Y(n_6817)
);

OR2x2_ASAP7_75t_L g6818 ( 
.A(n_6148),
.B(n_5915),
.Y(n_6818)
);

OAI21x1_ASAP7_75t_L g6819 ( 
.A1(n_6225),
.A2(n_5923),
.B(n_5852),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6231),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6237),
.Y(n_6821)
);

AND2x2_ASAP7_75t_L g6822 ( 
.A(n_6380),
.B(n_5502),
.Y(n_6822)
);

OR2x2_ASAP7_75t_L g6823 ( 
.A(n_6197),
.B(n_6427),
.Y(n_6823)
);

OR2x2_ASAP7_75t_L g6824 ( 
.A(n_6197),
.B(n_5915),
.Y(n_6824)
);

INVx2_ASAP7_75t_L g6825 ( 
.A(n_6129),
.Y(n_6825)
);

AND2x2_ASAP7_75t_L g6826 ( 
.A(n_6380),
.B(n_5543),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6129),
.Y(n_6827)
);

INVx2_ASAP7_75t_L g6828 ( 
.A(n_6135),
.Y(n_6828)
);

OR2x2_ASAP7_75t_L g6829 ( 
.A(n_6443),
.B(n_5915),
.Y(n_6829)
);

AND2x4_ASAP7_75t_L g6830 ( 
.A(n_6288),
.B(n_5834),
.Y(n_6830)
);

NOR2xp33_ASAP7_75t_SL g6831 ( 
.A(n_6150),
.B(n_5846),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6239),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_6245),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6380),
.B(n_5543),
.Y(n_6834)
);

OR2x2_ASAP7_75t_L g6835 ( 
.A(n_6608),
.B(n_5915),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_L g6836 ( 
.A(n_6384),
.B(n_5635),
.Y(n_6836)
);

OR2x2_ASAP7_75t_L g6837 ( 
.A(n_6340),
.B(n_6343),
.Y(n_6837)
);

OAI31xp33_ASAP7_75t_L g6838 ( 
.A1(n_6162),
.A2(n_5072),
.A3(n_6069),
.B(n_4917),
.Y(n_6838)
);

AND2x2_ASAP7_75t_L g6839 ( 
.A(n_6407),
.B(n_5543),
.Y(n_6839)
);

CKINVDCx6p67_ASAP7_75t_R g6840 ( 
.A(n_6488),
.Y(n_6840)
);

AND2x2_ASAP7_75t_L g6841 ( 
.A(n_6407),
.B(n_5590),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_6254),
.Y(n_6842)
);

NAND2xp5_ASAP7_75t_L g6843 ( 
.A(n_6384),
.B(n_5635),
.Y(n_6843)
);

INVx2_ASAP7_75t_L g6844 ( 
.A(n_6135),
.Y(n_6844)
);

INVx2_ASAP7_75t_L g6845 ( 
.A(n_6147),
.Y(n_6845)
);

AND2x4_ASAP7_75t_L g6846 ( 
.A(n_6335),
.B(n_5834),
.Y(n_6846)
);

NAND2xp5_ASAP7_75t_L g6847 ( 
.A(n_6434),
.B(n_6417),
.Y(n_6847)
);

INVx2_ASAP7_75t_L g6848 ( 
.A(n_6147),
.Y(n_6848)
);

OAI22xp5_ASAP7_75t_L g6849 ( 
.A1(n_6521),
.A2(n_4787),
.B1(n_5868),
.B2(n_6069),
.Y(n_6849)
);

INVx2_ASAP7_75t_L g6850 ( 
.A(n_6180),
.Y(n_6850)
);

NOR4xp25_ASAP7_75t_SL g6851 ( 
.A(n_6335),
.B(n_5765),
.C(n_5900),
.D(n_5772),
.Y(n_6851)
);

AND2x2_ASAP7_75t_L g6852 ( 
.A(n_6407),
.B(n_5590),
.Y(n_6852)
);

INVx2_ASAP7_75t_L g6853 ( 
.A(n_6180),
.Y(n_6853)
);

OR2x2_ASAP7_75t_L g6854 ( 
.A(n_6363),
.B(n_5915),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_6448),
.B(n_5590),
.Y(n_6855)
);

AND2x2_ASAP7_75t_L g6856 ( 
.A(n_6448),
.B(n_6265),
.Y(n_6856)
);

INVx2_ASAP7_75t_L g6857 ( 
.A(n_6191),
.Y(n_6857)
);

AND2x2_ASAP7_75t_L g6858 ( 
.A(n_6448),
.B(n_5704),
.Y(n_6858)
);

INVx1_ASAP7_75t_L g6859 ( 
.A(n_6258),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_6265),
.B(n_5704),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_L g6861 ( 
.A(n_6434),
.B(n_6369),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6369),
.B(n_5636),
.Y(n_6862)
);

AND2x2_ASAP7_75t_L g6863 ( 
.A(n_6188),
.B(n_5704),
.Y(n_6863)
);

INVx3_ASAP7_75t_L g6864 ( 
.A(n_6085),
.Y(n_6864)
);

INVx2_ASAP7_75t_L g6865 ( 
.A(n_6191),
.Y(n_6865)
);

INVx2_ASAP7_75t_L g6866 ( 
.A(n_6198),
.Y(n_6866)
);

AND2x4_ASAP7_75t_L g6867 ( 
.A(n_6188),
.B(n_5834),
.Y(n_6867)
);

BUFx3_ASAP7_75t_L g6868 ( 
.A(n_6116),
.Y(n_6868)
);

INVx2_ASAP7_75t_L g6869 ( 
.A(n_6198),
.Y(n_6869)
);

OR2x2_ASAP7_75t_L g6870 ( 
.A(n_6392),
.B(n_5732),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6264),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6267),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_6268),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6274),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6278),
.Y(n_6875)
);

INVx2_ASAP7_75t_L g6876 ( 
.A(n_6223),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6188),
.B(n_6200),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_6146),
.B(n_5636),
.Y(n_6878)
);

BUFx2_ASAP7_75t_L g6879 ( 
.A(n_6476),
.Y(n_6879)
);

INVx2_ASAP7_75t_L g6880 ( 
.A(n_6223),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_6165),
.B(n_6087),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6283),
.Y(n_6882)
);

INVxp67_ASAP7_75t_SL g6883 ( 
.A(n_6088),
.Y(n_6883)
);

AND2x4_ASAP7_75t_L g6884 ( 
.A(n_6200),
.B(n_5839),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6200),
.B(n_5738),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6211),
.B(n_5738),
.Y(n_6886)
);

OR2x2_ASAP7_75t_SL g6887 ( 
.A(n_6116),
.B(n_5905),
.Y(n_6887)
);

INVx2_ASAP7_75t_L g6888 ( 
.A(n_6262),
.Y(n_6888)
);

INVx2_ASAP7_75t_L g6889 ( 
.A(n_6262),
.Y(n_6889)
);

INVx3_ASAP7_75t_L g6890 ( 
.A(n_6426),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6294),
.Y(n_6891)
);

AND2x2_ASAP7_75t_L g6892 ( 
.A(n_6211),
.B(n_5738),
.Y(n_6892)
);

INVx2_ASAP7_75t_L g6893 ( 
.A(n_6088),
.Y(n_6893)
);

OR2x2_ASAP7_75t_L g6894 ( 
.A(n_6314),
.B(n_5732),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_L g6895 ( 
.A(n_6087),
.B(n_5638),
.Y(n_6895)
);

AND2x2_ASAP7_75t_L g6896 ( 
.A(n_6211),
.B(n_5838),
.Y(n_6896)
);

AND2x2_ASAP7_75t_L g6897 ( 
.A(n_6218),
.B(n_6069),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6299),
.Y(n_6898)
);

BUFx2_ASAP7_75t_L g6899 ( 
.A(n_6476),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_6092),
.Y(n_6900)
);

HB1xp67_ASAP7_75t_L g6901 ( 
.A(n_6548),
.Y(n_6901)
);

HB1xp67_ASAP7_75t_L g6902 ( 
.A(n_6559),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6304),
.Y(n_6903)
);

AND2x2_ASAP7_75t_L g6904 ( 
.A(n_6218),
.B(n_5839),
.Y(n_6904)
);

INVx2_ASAP7_75t_L g6905 ( 
.A(n_6092),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_6306),
.Y(n_6906)
);

BUFx2_ASAP7_75t_L g6907 ( 
.A(n_6487),
.Y(n_6907)
);

INVxp67_ASAP7_75t_SL g6908 ( 
.A(n_6099),
.Y(n_6908)
);

AND2x4_ASAP7_75t_L g6909 ( 
.A(n_6218),
.B(n_5839),
.Y(n_6909)
);

AND2x2_ASAP7_75t_L g6910 ( 
.A(n_6229),
.B(n_5839),
.Y(n_6910)
);

AND2x4_ASAP7_75t_L g6911 ( 
.A(n_6229),
.B(n_5884),
.Y(n_6911)
);

BUFx2_ASAP7_75t_L g6912 ( 
.A(n_6487),
.Y(n_6912)
);

BUFx2_ASAP7_75t_L g6913 ( 
.A(n_6488),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6313),
.Y(n_6914)
);

INVx2_ASAP7_75t_L g6915 ( 
.A(n_6099),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6322),
.Y(n_6916)
);

INVx3_ASAP7_75t_L g6917 ( 
.A(n_6510),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6344),
.Y(n_6918)
);

INVx2_ASAP7_75t_L g6919 ( 
.A(n_6101),
.Y(n_6919)
);

AND2x2_ASAP7_75t_L g6920 ( 
.A(n_6229),
.B(n_6325),
.Y(n_6920)
);

AND2x2_ASAP7_75t_L g6921 ( 
.A(n_6325),
.B(n_5884),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6347),
.Y(n_6922)
);

INVx2_ASAP7_75t_L g6923 ( 
.A(n_6101),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6354),
.Y(n_6924)
);

NAND2xp5_ASAP7_75t_L g6925 ( 
.A(n_6087),
.B(n_5638),
.Y(n_6925)
);

OAI21xp5_ASAP7_75t_SL g6926 ( 
.A1(n_6473),
.A2(n_5979),
.B(n_5905),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6325),
.B(n_6457),
.Y(n_6927)
);

BUFx2_ASAP7_75t_L g6928 ( 
.A(n_6160),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_L g6929 ( 
.A(n_6617),
.B(n_5587),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6355),
.Y(n_6930)
);

HB1xp67_ASAP7_75t_L g6931 ( 
.A(n_6573),
.Y(n_6931)
);

AND2x2_ASAP7_75t_L g6932 ( 
.A(n_6457),
.B(n_5884),
.Y(n_6932)
);

INVx2_ASAP7_75t_L g6933 ( 
.A(n_6112),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6360),
.Y(n_6934)
);

BUFx3_ASAP7_75t_L g6935 ( 
.A(n_6116),
.Y(n_6935)
);

OR2x6_ASAP7_75t_L g6936 ( 
.A(n_6326),
.B(n_5905),
.Y(n_6936)
);

INVx2_ASAP7_75t_L g6937 ( 
.A(n_6112),
.Y(n_6937)
);

AND2x2_ASAP7_75t_L g6938 ( 
.A(n_6457),
.B(n_5884),
.Y(n_6938)
);

INVx3_ASAP7_75t_L g6939 ( 
.A(n_6510),
.Y(n_6939)
);

NAND2xp5_ASAP7_75t_L g6940 ( 
.A(n_6113),
.B(n_5994),
.Y(n_6940)
);

AND2x2_ASAP7_75t_L g6941 ( 
.A(n_6457),
.B(n_5924),
.Y(n_6941)
);

AOI22xp33_ASAP7_75t_SL g6942 ( 
.A1(n_6588),
.A2(n_5868),
.B1(n_5663),
.B2(n_5574),
.Y(n_6942)
);

NAND2xp5_ASAP7_75t_SL g6943 ( 
.A(n_6492),
.B(n_5654),
.Y(n_6943)
);

INVx1_ASAP7_75t_SL g6944 ( 
.A(n_6370),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6396),
.B(n_5924),
.Y(n_6945)
);

BUFx6f_ASAP7_75t_L g6946 ( 
.A(n_6116),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6374),
.Y(n_6947)
);

INVx3_ASAP7_75t_L g6948 ( 
.A(n_6510),
.Y(n_6948)
);

AOI221xp5_ASAP7_75t_L g6949 ( 
.A1(n_6600),
.A2(n_5926),
.B1(n_5979),
.B2(n_6044),
.C(n_5905),
.Y(n_6949)
);

INVx3_ASAP7_75t_L g6950 ( 
.A(n_6357),
.Y(n_6950)
);

AOI22xp5_ASAP7_75t_L g6951 ( 
.A1(n_6128),
.A2(n_5868),
.B1(n_6046),
.B2(n_5574),
.Y(n_6951)
);

OAI221xp5_ASAP7_75t_L g6952 ( 
.A1(n_6551),
.A2(n_5977),
.B1(n_6062),
.B2(n_5921),
.C(n_5840),
.Y(n_6952)
);

AOI22xp33_ASAP7_75t_L g6953 ( 
.A1(n_6566),
.A2(n_5492),
.B1(n_5486),
.B2(n_5921),
.Y(n_6953)
);

OR2x2_ASAP7_75t_L g6954 ( 
.A(n_6130),
.B(n_5761),
.Y(n_6954)
);

INVx2_ASAP7_75t_L g6955 ( 
.A(n_6114),
.Y(n_6955)
);

INVx2_ASAP7_75t_L g6956 ( 
.A(n_6114),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6377),
.Y(n_6957)
);

NAND2x1_ASAP7_75t_L g6958 ( 
.A(n_6357),
.B(n_5924),
.Y(n_6958)
);

AND2x2_ASAP7_75t_L g6959 ( 
.A(n_6396),
.B(n_5924),
.Y(n_6959)
);

INVx3_ASAP7_75t_L g6960 ( 
.A(n_6357),
.Y(n_6960)
);

INVx2_ASAP7_75t_R g6961 ( 
.A(n_6526),
.Y(n_6961)
);

AND2x2_ASAP7_75t_L g6962 ( 
.A(n_6398),
.B(n_5650),
.Y(n_6962)
);

INVx2_ASAP7_75t_L g6963 ( 
.A(n_6550),
.Y(n_6963)
);

INVx2_ASAP7_75t_SL g6964 ( 
.A(n_6526),
.Y(n_6964)
);

AND2x2_ASAP7_75t_L g6965 ( 
.A(n_6398),
.B(n_5650),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6385),
.Y(n_6966)
);

INVxp67_ASAP7_75t_SL g6967 ( 
.A(n_6277),
.Y(n_6967)
);

OR2x2_ASAP7_75t_L g6968 ( 
.A(n_6130),
.B(n_5620),
.Y(n_6968)
);

AND2x2_ASAP7_75t_L g6969 ( 
.A(n_6582),
.B(n_5921),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6386),
.Y(n_6970)
);

AND2x2_ASAP7_75t_L g6971 ( 
.A(n_6187),
.B(n_5977),
.Y(n_6971)
);

AND2x2_ASAP7_75t_L g6972 ( 
.A(n_6187),
.B(n_5977),
.Y(n_6972)
);

AND2x2_ASAP7_75t_L g6973 ( 
.A(n_6187),
.B(n_6199),
.Y(n_6973)
);

INVxp67_ASAP7_75t_R g6974 ( 
.A(n_6561),
.Y(n_6974)
);

HB1xp67_ASAP7_75t_L g6975 ( 
.A(n_6592),
.Y(n_6975)
);

NAND2x1_ASAP7_75t_L g6976 ( 
.A(n_6378),
.B(n_5784),
.Y(n_6976)
);

INVx2_ASAP7_75t_L g6977 ( 
.A(n_6550),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6388),
.Y(n_6978)
);

BUFx3_ASAP7_75t_L g6979 ( 
.A(n_6134),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6550),
.Y(n_6980)
);

INVx2_ASAP7_75t_L g6981 ( 
.A(n_6131),
.Y(n_6981)
);

INVx2_ASAP7_75t_L g6982 ( 
.A(n_6131),
.Y(n_6982)
);

OR2x2_ASAP7_75t_L g6983 ( 
.A(n_6328),
.B(n_5620),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6131),
.Y(n_6984)
);

NAND2xp5_ASAP7_75t_L g6985 ( 
.A(n_6575),
.B(n_6024),
.Y(n_6985)
);

INVx2_ASAP7_75t_SL g6986 ( 
.A(n_6526),
.Y(n_6986)
);

INVx2_ASAP7_75t_L g6987 ( 
.A(n_6275),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6389),
.Y(n_6988)
);

INVx2_ASAP7_75t_L g6989 ( 
.A(n_6275),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6393),
.Y(n_6990)
);

AND2x2_ASAP7_75t_L g6991 ( 
.A(n_6187),
.B(n_6062),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6395),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_6399),
.Y(n_6993)
);

INVxp67_ASAP7_75t_L g6994 ( 
.A(n_6315),
.Y(n_6994)
);

BUFx2_ASAP7_75t_L g6995 ( 
.A(n_6366),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6400),
.Y(n_6996)
);

AND2x4_ASAP7_75t_L g6997 ( 
.A(n_6199),
.B(n_5654),
.Y(n_6997)
);

INVx2_ASAP7_75t_SL g6998 ( 
.A(n_6526),
.Y(n_6998)
);

INVx2_ASAP7_75t_L g6999 ( 
.A(n_6275),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6402),
.Y(n_7000)
);

AND2x2_ASAP7_75t_L g7001 ( 
.A(n_6199),
.B(n_6062),
.Y(n_7001)
);

HB1xp67_ASAP7_75t_L g7002 ( 
.A(n_6602),
.Y(n_7002)
);

INVx1_ASAP7_75t_L g7003 ( 
.A(n_6406),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6309),
.Y(n_7004)
);

INVx2_ASAP7_75t_L g7005 ( 
.A(n_6309),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6577),
.B(n_6619),
.Y(n_7006)
);

INVx1_ASAP7_75t_L g7007 ( 
.A(n_6409),
.Y(n_7007)
);

NAND2xp5_ASAP7_75t_L g7008 ( 
.A(n_6242),
.B(n_6024),
.Y(n_7008)
);

NAND2xp5_ASAP7_75t_L g7009 ( 
.A(n_6596),
.B(n_6026),
.Y(n_7009)
);

AND2x2_ASAP7_75t_L g7010 ( 
.A(n_6619),
.B(n_5790),
.Y(n_7010)
);

BUFx2_ASAP7_75t_L g7011 ( 
.A(n_6366),
.Y(n_7011)
);

AOI22xp33_ASAP7_75t_L g7012 ( 
.A1(n_6612),
.A2(n_5486),
.B1(n_6044),
.B2(n_5979),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6410),
.Y(n_7013)
);

AND2x2_ASAP7_75t_L g7014 ( 
.A(n_6199),
.B(n_6042),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6415),
.Y(n_7015)
);

HB1xp67_ASAP7_75t_L g7016 ( 
.A(n_6606),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6419),
.Y(n_7017)
);

AND2x2_ASAP7_75t_L g7018 ( 
.A(n_6512),
.B(n_6042),
.Y(n_7018)
);

CKINVDCx5p33_ASAP7_75t_R g7019 ( 
.A(n_6376),
.Y(n_7019)
);

INVx2_ASAP7_75t_L g7020 ( 
.A(n_6309),
.Y(n_7020)
);

NAND2xp5_ASAP7_75t_L g7021 ( 
.A(n_6587),
.B(n_6026),
.Y(n_7021)
);

INVx1_ASAP7_75t_L g7022 ( 
.A(n_6425),
.Y(n_7022)
);

OR2x2_ASAP7_75t_L g7023 ( 
.A(n_6328),
.B(n_5624),
.Y(n_7023)
);

AND2x2_ASAP7_75t_L g7024 ( 
.A(n_6512),
.B(n_6051),
.Y(n_7024)
);

INVx3_ASAP7_75t_L g7025 ( 
.A(n_6378),
.Y(n_7025)
);

INVx2_ASAP7_75t_L g7026 ( 
.A(n_6310),
.Y(n_7026)
);

INVx2_ASAP7_75t_L g7027 ( 
.A(n_6310),
.Y(n_7027)
);

NAND2xp5_ASAP7_75t_L g7028 ( 
.A(n_6558),
.B(n_5994),
.Y(n_7028)
);

INVx2_ASAP7_75t_L g7029 ( 
.A(n_6310),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6558),
.B(n_6051),
.Y(n_7030)
);

CKINVDCx20_ASAP7_75t_R g7031 ( 
.A(n_6370),
.Y(n_7031)
);

INVx1_ASAP7_75t_L g7032 ( 
.A(n_6430),
.Y(n_7032)
);

OAI21x1_ASAP7_75t_L g7033 ( 
.A1(n_6225),
.A2(n_5923),
.B(n_5852),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_6179),
.B(n_4835),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6435),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_6431),
.Y(n_7036)
);

AOI22xp33_ASAP7_75t_L g7037 ( 
.A1(n_6125),
.A2(n_5486),
.B1(n_6044),
.B2(n_5979),
.Y(n_7037)
);

INVxp67_ASAP7_75t_R g7038 ( 
.A(n_6561),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6179),
.B(n_6077),
.Y(n_7039)
);

INVxp67_ASAP7_75t_L g7040 ( 
.A(n_6315),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6438),
.Y(n_7041)
);

INVx3_ASAP7_75t_L g7042 ( 
.A(n_6378),
.Y(n_7042)
);

INVx1_ASAP7_75t_SL g7043 ( 
.A(n_6387),
.Y(n_7043)
);

INVx2_ASAP7_75t_L g7044 ( 
.A(n_6431),
.Y(n_7044)
);

INVx2_ASAP7_75t_L g7045 ( 
.A(n_6431),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6439),
.Y(n_7046)
);

INVx1_ASAP7_75t_L g7047 ( 
.A(n_6444),
.Y(n_7047)
);

CKINVDCx20_ASAP7_75t_R g7048 ( 
.A(n_6376),
.Y(n_7048)
);

NAND2xp5_ASAP7_75t_L g7049 ( 
.A(n_6315),
.B(n_5654),
.Y(n_7049)
);

AND2x4_ASAP7_75t_L g7050 ( 
.A(n_6366),
.B(n_5654),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6450),
.Y(n_7051)
);

OR2x2_ASAP7_75t_L g7052 ( 
.A(n_6158),
.B(n_5624),
.Y(n_7052)
);

INVx2_ASAP7_75t_SL g7053 ( 
.A(n_6526),
.Y(n_7053)
);

BUFx6f_ASAP7_75t_L g7054 ( 
.A(n_6134),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_6452),
.Y(n_7055)
);

AND2x4_ASAP7_75t_L g7056 ( 
.A(n_6366),
.B(n_5654),
.Y(n_7056)
);

AND2x2_ASAP7_75t_L g7057 ( 
.A(n_6185),
.B(n_6077),
.Y(n_7057)
);

INVx1_ASAP7_75t_L g7058 ( 
.A(n_6460),
.Y(n_7058)
);

NAND2xp5_ASAP7_75t_L g7059 ( 
.A(n_6315),
.B(n_5979),
.Y(n_7059)
);

OR2x2_ASAP7_75t_L g7060 ( 
.A(n_6158),
.B(n_5451),
.Y(n_7060)
);

BUFx2_ASAP7_75t_L g7061 ( 
.A(n_6394),
.Y(n_7061)
);

OR2x2_ASAP7_75t_L g7062 ( 
.A(n_6312),
.B(n_5506),
.Y(n_7062)
);

INVxp67_ASAP7_75t_SL g7063 ( 
.A(n_6081),
.Y(n_7063)
);

AND2x2_ASAP7_75t_L g7064 ( 
.A(n_6185),
.B(n_5980),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6461),
.Y(n_7065)
);

AOI22xp33_ASAP7_75t_SL g7066 ( 
.A1(n_6120),
.A2(n_6046),
.B1(n_5574),
.B2(n_5359),
.Y(n_7066)
);

AND2x2_ASAP7_75t_L g7067 ( 
.A(n_6206),
.B(n_5980),
.Y(n_7067)
);

INVx2_ASAP7_75t_SL g7068 ( 
.A(n_6217),
.Y(n_7068)
);

HB1xp67_ASAP7_75t_L g7069 ( 
.A(n_6620),
.Y(n_7069)
);

INVx2_ASAP7_75t_SL g7070 ( 
.A(n_6217),
.Y(n_7070)
);

INVx3_ASAP7_75t_L g7071 ( 
.A(n_6382),
.Y(n_7071)
);

INVx5_ASAP7_75t_L g7072 ( 
.A(n_6202),
.Y(n_7072)
);

AND2x2_ASAP7_75t_L g7073 ( 
.A(n_6418),
.B(n_6420),
.Y(n_7073)
);

HB1xp67_ASAP7_75t_L g7074 ( 
.A(n_6462),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6623),
.Y(n_7075)
);

AO21x2_ASAP7_75t_L g7076 ( 
.A1(n_6981),
.A2(n_6553),
.B(n_6320),
.Y(n_7076)
);

OR2x2_ASAP7_75t_L g7077 ( 
.A(n_6801),
.B(n_6286),
.Y(n_7077)
);

INVx2_ASAP7_75t_L g7078 ( 
.A(n_6721),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6623),
.Y(n_7079)
);

AND2x2_ASAP7_75t_SL g7080 ( 
.A(n_6668),
.B(n_6189),
.Y(n_7080)
);

BUFx6f_ASAP7_75t_L g7081 ( 
.A(n_6946),
.Y(n_7081)
);

INVx2_ASAP7_75t_L g7082 ( 
.A(n_6740),
.Y(n_7082)
);

INVxp67_ASAP7_75t_SL g7083 ( 
.A(n_6864),
.Y(n_7083)
);

AND2x2_ASAP7_75t_L g7084 ( 
.A(n_6633),
.B(n_6102),
.Y(n_7084)
);

AND2x2_ASAP7_75t_L g7085 ( 
.A(n_6636),
.B(n_6102),
.Y(n_7085)
);

INVx2_ASAP7_75t_L g7086 ( 
.A(n_6721),
.Y(n_7086)
);

AND2x2_ASAP7_75t_L g7087 ( 
.A(n_6928),
.B(n_6102),
.Y(n_7087)
);

OR2x2_ASAP7_75t_L g7088 ( 
.A(n_6674),
.B(n_6286),
.Y(n_7088)
);

NOR2x1_ASAP7_75t_L g7089 ( 
.A(n_6627),
.B(n_6326),
.Y(n_7089)
);

INVx3_ASAP7_75t_L g7090 ( 
.A(n_6721),
.Y(n_7090)
);

INVx2_ASAP7_75t_L g7091 ( 
.A(n_6917),
.Y(n_7091)
);

BUFx2_ASAP7_75t_L g7092 ( 
.A(n_6740),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6632),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6665),
.B(n_6102),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6917),
.Y(n_7095)
);

NAND2xp5_ASAP7_75t_L g7096 ( 
.A(n_6694),
.B(n_6464),
.Y(n_7096)
);

INVx2_ASAP7_75t_L g7097 ( 
.A(n_6917),
.Y(n_7097)
);

AND2x4_ASAP7_75t_L g7098 ( 
.A(n_6777),
.B(n_6383),
.Y(n_7098)
);

INVx2_ASAP7_75t_L g7099 ( 
.A(n_6939),
.Y(n_7099)
);

INVxp67_ASAP7_75t_SL g7100 ( 
.A(n_6864),
.Y(n_7100)
);

AND2x2_ASAP7_75t_L g7101 ( 
.A(n_6777),
.B(n_6201),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_6939),
.Y(n_7102)
);

OR2x2_ASAP7_75t_SL g7103 ( 
.A(n_6683),
.B(n_6134),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_6632),
.Y(n_7104)
);

AND2x2_ASAP7_75t_L g7105 ( 
.A(n_6860),
.B(n_6394),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_L g7106 ( 
.A(n_6694),
.B(n_6470),
.Y(n_7106)
);

OR2x2_ASAP7_75t_L g7107 ( 
.A(n_6752),
.B(n_6273),
.Y(n_7107)
);

AND2x2_ASAP7_75t_L g7108 ( 
.A(n_6856),
.B(n_6394),
.Y(n_7108)
);

INVx4_ASAP7_75t_L g7109 ( 
.A(n_7072),
.Y(n_7109)
);

NAND2xp5_ASAP7_75t_L g7110 ( 
.A(n_6737),
.B(n_6479),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6637),
.Y(n_7111)
);

INVx2_ASAP7_75t_L g7112 ( 
.A(n_6939),
.Y(n_7112)
);

BUFx6f_ASAP7_75t_L g7113 ( 
.A(n_6946),
.Y(n_7113)
);

INVx2_ASAP7_75t_L g7114 ( 
.A(n_6948),
.Y(n_7114)
);

HB1xp67_ASAP7_75t_L g7115 ( 
.A(n_6637),
.Y(n_7115)
);

AND2x2_ASAP7_75t_L g7116 ( 
.A(n_6630),
.B(n_6394),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_6737),
.B(n_6480),
.Y(n_7117)
);

AOI22xp33_ASAP7_75t_SL g7118 ( 
.A1(n_6952),
.A2(n_6320),
.B1(n_5574),
.B2(n_6046),
.Y(n_7118)
);

AND2x4_ASAP7_75t_L g7119 ( 
.A(n_6634),
.B(n_6383),
.Y(n_7119)
);

INVx2_ASAP7_75t_L g7120 ( 
.A(n_6868),
.Y(n_7120)
);

INVx2_ASAP7_75t_L g7121 ( 
.A(n_6948),
.Y(n_7121)
);

AND2x2_ASAP7_75t_L g7122 ( 
.A(n_6749),
.B(n_6134),
.Y(n_7122)
);

INVxp67_ASAP7_75t_SL g7123 ( 
.A(n_6864),
.Y(n_7123)
);

OR2x2_ASAP7_75t_L g7124 ( 
.A(n_6778),
.B(n_6273),
.Y(n_7124)
);

HB1xp67_ASAP7_75t_L g7125 ( 
.A(n_6662),
.Y(n_7125)
);

INVx2_ASAP7_75t_L g7126 ( 
.A(n_6948),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6974),
.B(n_6154),
.Y(n_7127)
);

AND2x2_ASAP7_75t_L g7128 ( 
.A(n_7038),
.B(n_6639),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6662),
.Y(n_7129)
);

INVx4_ASAP7_75t_L g7130 ( 
.A(n_7072),
.Y(n_7130)
);

HB1xp67_ASAP7_75t_L g7131 ( 
.A(n_6666),
.Y(n_7131)
);

AND2x2_ASAP7_75t_L g7132 ( 
.A(n_6678),
.B(n_6154),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6666),
.Y(n_7133)
);

INVx2_ASAP7_75t_L g7134 ( 
.A(n_6868),
.Y(n_7134)
);

BUFx3_ASAP7_75t_L g7135 ( 
.A(n_7031),
.Y(n_7135)
);

AND2x2_ASAP7_75t_L g7136 ( 
.A(n_6680),
.B(n_6154),
.Y(n_7136)
);

INVx2_ASAP7_75t_L g7137 ( 
.A(n_6935),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6935),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_6693),
.Y(n_7139)
);

INVx2_ASAP7_75t_SL g7140 ( 
.A(n_7072),
.Y(n_7140)
);

NAND2xp5_ASAP7_75t_L g7141 ( 
.A(n_6756),
.B(n_6594),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6979),
.Y(n_7142)
);

BUFx3_ASAP7_75t_L g7143 ( 
.A(n_7031),
.Y(n_7143)
);

INVx4_ASAP7_75t_SL g7144 ( 
.A(n_6946),
.Y(n_7144)
);

AND2x2_ASAP7_75t_L g7145 ( 
.A(n_6746),
.B(n_6154),
.Y(n_7145)
);

AND2x2_ASAP7_75t_L g7146 ( 
.A(n_6631),
.B(n_6326),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6693),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6697),
.Y(n_7148)
);

INVx2_ASAP7_75t_L g7149 ( 
.A(n_6979),
.Y(n_7149)
);

INVx2_ASAP7_75t_L g7150 ( 
.A(n_6775),
.Y(n_7150)
);

AND2x2_ASAP7_75t_L g7151 ( 
.A(n_6822),
.B(n_6326),
.Y(n_7151)
);

INVx1_ASAP7_75t_L g7152 ( 
.A(n_6697),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6728),
.Y(n_7153)
);

NAND2xp5_ASAP7_75t_L g7154 ( 
.A(n_6756),
.B(n_6656),
.Y(n_7154)
);

AND2x2_ASAP7_75t_L g7155 ( 
.A(n_6826),
.B(n_6834),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6728),
.Y(n_7156)
);

AND2x4_ASAP7_75t_L g7157 ( 
.A(n_6634),
.B(n_6383),
.Y(n_7157)
);

AND2x2_ASAP7_75t_L g7158 ( 
.A(n_6839),
.B(n_6331),
.Y(n_7158)
);

INVx1_ASAP7_75t_L g7159 ( 
.A(n_6780),
.Y(n_7159)
);

AND2x2_ASAP7_75t_L g7160 ( 
.A(n_6841),
.B(n_6331),
.Y(n_7160)
);

AND2x2_ASAP7_75t_L g7161 ( 
.A(n_6852),
.B(n_6331),
.Y(n_7161)
);

INVx3_ASAP7_75t_L g7162 ( 
.A(n_6775),
.Y(n_7162)
);

INVx2_ASAP7_75t_L g7163 ( 
.A(n_6725),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_6780),
.Y(n_7164)
);

AND2x2_ASAP7_75t_L g7165 ( 
.A(n_6855),
.B(n_6331),
.Y(n_7165)
);

INVx2_ASAP7_75t_L g7166 ( 
.A(n_6725),
.Y(n_7166)
);

OR2x2_ASAP7_75t_L g7167 ( 
.A(n_6792),
.B(n_6349),
.Y(n_7167)
);

HB1xp67_ASAP7_75t_L g7168 ( 
.A(n_6800),
.Y(n_7168)
);

AND2x4_ASAP7_75t_L g7169 ( 
.A(n_6635),
.B(n_6383),
.Y(n_7169)
);

AND2x2_ASAP7_75t_L g7170 ( 
.A(n_6858),
.B(n_6349),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_6800),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_6901),
.Y(n_7172)
);

NAND2xp5_ASAP7_75t_L g7173 ( 
.A(n_6679),
.B(n_6605),
.Y(n_7173)
);

AND2x2_ASAP7_75t_L g7174 ( 
.A(n_6815),
.B(n_6349),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6901),
.Y(n_7175)
);

AND2x2_ASAP7_75t_L g7176 ( 
.A(n_6816),
.B(n_6349),
.Y(n_7176)
);

HB1xp67_ASAP7_75t_L g7177 ( 
.A(n_6902),
.Y(n_7177)
);

NOR2x1_ASAP7_75t_SL g7178 ( 
.A(n_6936),
.B(n_6358),
.Y(n_7178)
);

AND2x2_ASAP7_75t_L g7179 ( 
.A(n_6817),
.B(n_6358),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6902),
.Y(n_7180)
);

HB1xp67_ASAP7_75t_L g7181 ( 
.A(n_6931),
.Y(n_7181)
);

INVx3_ASAP7_75t_L g7182 ( 
.A(n_6782),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_6679),
.B(n_6609),
.Y(n_7183)
);

INVx2_ASAP7_75t_L g7184 ( 
.A(n_6725),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_6931),
.Y(n_7185)
);

NAND2xp5_ASAP7_75t_L g7186 ( 
.A(n_6975),
.B(n_6485),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_6975),
.Y(n_7187)
);

INVx2_ASAP7_75t_L g7188 ( 
.A(n_6786),
.Y(n_7188)
);

AND2x2_ASAP7_75t_L g7189 ( 
.A(n_6791),
.B(n_6358),
.Y(n_7189)
);

INVx2_ASAP7_75t_L g7190 ( 
.A(n_6786),
.Y(n_7190)
);

BUFx6f_ASAP7_75t_L g7191 ( 
.A(n_6946),
.Y(n_7191)
);

NOR2x1_ASAP7_75t_SL g7192 ( 
.A(n_6936),
.B(n_6358),
.Y(n_7192)
);

INVxp67_ASAP7_75t_SL g7193 ( 
.A(n_7063),
.Y(n_7193)
);

OR2x2_ASAP7_75t_L g7194 ( 
.A(n_6771),
.B(n_6312),
.Y(n_7194)
);

NAND2xp5_ASAP7_75t_L g7195 ( 
.A(n_7002),
.B(n_6490),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_7002),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_7016),
.Y(n_7197)
);

AND2x4_ASAP7_75t_L g7198 ( 
.A(n_6635),
.B(n_6428),
.Y(n_7198)
);

INVx3_ASAP7_75t_L g7199 ( 
.A(n_6782),
.Y(n_7199)
);

AND2x2_ASAP7_75t_L g7200 ( 
.A(n_7034),
.B(n_6202),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_L g7201 ( 
.A(n_7016),
.B(n_6491),
.Y(n_7201)
);

AND2x2_ASAP7_75t_L g7202 ( 
.A(n_6710),
.B(n_6428),
.Y(n_7202)
);

AND2x2_ASAP7_75t_L g7203 ( 
.A(n_6809),
.B(n_6428),
.Y(n_7203)
);

HB1xp67_ASAP7_75t_L g7204 ( 
.A(n_7069),
.Y(n_7204)
);

INVx2_ASAP7_75t_L g7205 ( 
.A(n_6786),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_7069),
.Y(n_7206)
);

INVx2_ASAP7_75t_L g7207 ( 
.A(n_6830),
.Y(n_7207)
);

INVx2_ASAP7_75t_L g7208 ( 
.A(n_6830),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_7074),
.Y(n_7209)
);

AND2x2_ASAP7_75t_L g7210 ( 
.A(n_6969),
.B(n_6428),
.Y(n_7210)
);

INVxp67_ASAP7_75t_L g7211 ( 
.A(n_6648),
.Y(n_7211)
);

AOI22xp33_ASAP7_75t_L g7212 ( 
.A1(n_6668),
.A2(n_6320),
.B1(n_6532),
.B2(n_6348),
.Y(n_7212)
);

INVx5_ASAP7_75t_L g7213 ( 
.A(n_7054),
.Y(n_7213)
);

NOR2xp33_ASAP7_75t_L g7214 ( 
.A(n_6688),
.B(n_6387),
.Y(n_7214)
);

AND2x2_ASAP7_75t_L g7215 ( 
.A(n_6750),
.B(n_6544),
.Y(n_7215)
);

AND2x2_ASAP7_75t_L g7216 ( 
.A(n_6751),
.B(n_6544),
.Y(n_7216)
);

INVx2_ASAP7_75t_L g7217 ( 
.A(n_6830),
.Y(n_7217)
);

INVxp67_ASAP7_75t_SL g7218 ( 
.A(n_7063),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_L g7219 ( 
.A(n_6626),
.B(n_6591),
.Y(n_7219)
);

HB1xp67_ASAP7_75t_L g7220 ( 
.A(n_6626),
.Y(n_7220)
);

NAND2xp5_ASAP7_75t_L g7221 ( 
.A(n_6640),
.B(n_6498),
.Y(n_7221)
);

BUFx3_ASAP7_75t_L g7222 ( 
.A(n_7048),
.Y(n_7222)
);

OR2x2_ASAP7_75t_L g7223 ( 
.A(n_6784),
.B(n_6323),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_6754),
.B(n_6544),
.Y(n_7224)
);

OR2x2_ASAP7_75t_L g7225 ( 
.A(n_6714),
.B(n_6323),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_7074),
.Y(n_7226)
);

AND2x2_ASAP7_75t_L g7227 ( 
.A(n_6790),
.B(n_6544),
.Y(n_7227)
);

INVx2_ASAP7_75t_L g7228 ( 
.A(n_6846),
.Y(n_7228)
);

BUFx6f_ASAP7_75t_L g7229 ( 
.A(n_7054),
.Y(n_7229)
);

AND2x2_ASAP7_75t_L g7230 ( 
.A(n_6790),
.B(n_6555),
.Y(n_7230)
);

OR2x2_ASAP7_75t_L g7231 ( 
.A(n_6847),
.B(n_6474),
.Y(n_7231)
);

AND2x2_ASAP7_75t_L g7232 ( 
.A(n_6739),
.B(n_6555),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_6640),
.Y(n_7233)
);

INVx2_ASAP7_75t_SL g7234 ( 
.A(n_7072),
.Y(n_7234)
);

INVx1_ASAP7_75t_L g7235 ( 
.A(n_6649),
.Y(n_7235)
);

BUFx12f_ASAP7_75t_L g7236 ( 
.A(n_7019),
.Y(n_7236)
);

INVx2_ASAP7_75t_L g7237 ( 
.A(n_7054),
.Y(n_7237)
);

AND2x2_ASAP7_75t_L g7238 ( 
.A(n_6739),
.B(n_6555),
.Y(n_7238)
);

HB1xp67_ASAP7_75t_L g7239 ( 
.A(n_6649),
.Y(n_7239)
);

NOR2x1_ASAP7_75t_L g7240 ( 
.A(n_6926),
.B(n_6555),
.Y(n_7240)
);

INVx4_ASAP7_75t_L g7241 ( 
.A(n_7054),
.Y(n_7241)
);

INVx2_ASAP7_75t_L g7242 ( 
.A(n_6776),
.Y(n_7242)
);

AND2x2_ASAP7_75t_L g7243 ( 
.A(n_6685),
.B(n_6044),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_6651),
.Y(n_7244)
);

INVx1_ASAP7_75t_SL g7245 ( 
.A(n_7048),
.Y(n_7245)
);

AND2x2_ASAP7_75t_L g7246 ( 
.A(n_6689),
.B(n_6044),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_SL g7247 ( 
.A(n_6942),
.B(n_6364),
.Y(n_7247)
);

INVxp67_ASAP7_75t_L g7248 ( 
.A(n_6729),
.Y(n_7248)
);

INVx2_ASAP7_75t_L g7249 ( 
.A(n_6776),
.Y(n_7249)
);

INVx2_ASAP7_75t_L g7250 ( 
.A(n_6776),
.Y(n_7250)
);

AND2x2_ASAP7_75t_L g7251 ( 
.A(n_6628),
.B(n_6863),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6651),
.Y(n_7252)
);

HB1xp67_ASAP7_75t_L g7253 ( 
.A(n_6653),
.Y(n_7253)
);

AOI22xp33_ASAP7_75t_L g7254 ( 
.A1(n_6807),
.A2(n_6543),
.B1(n_6348),
.B2(n_6601),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_L g7255 ( 
.A(n_6653),
.B(n_6499),
.Y(n_7255)
);

INVx1_ASAP7_75t_L g7256 ( 
.A(n_6657),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_6657),
.Y(n_7257)
);

HB1xp67_ASAP7_75t_L g7258 ( 
.A(n_6621),
.Y(n_7258)
);

INVx1_ASAP7_75t_L g7259 ( 
.A(n_6654),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_6885),
.B(n_6886),
.Y(n_7260)
);

AND2x2_ASAP7_75t_L g7261 ( 
.A(n_6892),
.B(n_6209),
.Y(n_7261)
);

AND2x2_ASAP7_75t_L g7262 ( 
.A(n_6701),
.B(n_6301),
.Y(n_7262)
);

HB1xp67_ASAP7_75t_L g7263 ( 
.A(n_6625),
.Y(n_7263)
);

INVx1_ASAP7_75t_L g7264 ( 
.A(n_6658),
.Y(n_7264)
);

BUFx2_ASAP7_75t_L g7265 ( 
.A(n_6840),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_6663),
.Y(n_7266)
);

BUFx3_ASAP7_75t_L g7267 ( 
.A(n_6887),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_6669),
.Y(n_7268)
);

INVxp67_ASAP7_75t_SL g7269 ( 
.A(n_6981),
.Y(n_7269)
);

AND2x2_ASAP7_75t_L g7270 ( 
.A(n_6703),
.B(n_6302),
.Y(n_7270)
);

BUFx2_ASAP7_75t_L g7271 ( 
.A(n_6840),
.Y(n_7271)
);

INVx2_ASAP7_75t_L g7272 ( 
.A(n_6846),
.Y(n_7272)
);

HB1xp67_ASAP7_75t_L g7273 ( 
.A(n_6629),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_L g7274 ( 
.A(n_6638),
.B(n_6503),
.Y(n_7274)
);

INVx1_ASAP7_75t_L g7275 ( 
.A(n_6672),
.Y(n_7275)
);

AND2x2_ASAP7_75t_L g7276 ( 
.A(n_6704),
.B(n_6206),
.Y(n_7276)
);

OR2x2_ASAP7_75t_L g7277 ( 
.A(n_6823),
.B(n_6445),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_6677),
.Y(n_7278)
);

AND2x2_ASAP7_75t_L g7279 ( 
.A(n_6706),
.B(n_6207),
.Y(n_7279)
);

AND2x2_ASAP7_75t_L g7280 ( 
.A(n_6708),
.B(n_6207),
.Y(n_7280)
);

INVx2_ASAP7_75t_L g7281 ( 
.A(n_6846),
.Y(n_7281)
);

INVx2_ASAP7_75t_L g7282 ( 
.A(n_6736),
.Y(n_7282)
);

INVx2_ASAP7_75t_L g7283 ( 
.A(n_6736),
.Y(n_7283)
);

AND2x2_ASAP7_75t_L g7284 ( 
.A(n_6711),
.B(n_6208),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_6682),
.Y(n_7285)
);

INVx2_ASAP7_75t_L g7286 ( 
.A(n_6736),
.Y(n_7286)
);

NAND2xp5_ASAP7_75t_L g7287 ( 
.A(n_6643),
.B(n_6589),
.Y(n_7287)
);

INVx2_ASAP7_75t_SL g7288 ( 
.A(n_6675),
.Y(n_7288)
);

OR2x2_ASAP7_75t_L g7289 ( 
.A(n_6690),
.B(n_6454),
.Y(n_7289)
);

AND2x2_ASAP7_75t_L g7290 ( 
.A(n_6726),
.B(n_6208),
.Y(n_7290)
);

INVx3_ASAP7_75t_L g7291 ( 
.A(n_6797),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_6687),
.Y(n_7292)
);

HB1xp67_ASAP7_75t_L g7293 ( 
.A(n_6645),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_6692),
.Y(n_7294)
);

BUFx3_ASAP7_75t_L g7295 ( 
.A(n_6797),
.Y(n_7295)
);

INVx3_ASAP7_75t_L g7296 ( 
.A(n_6890),
.Y(n_7296)
);

AND2x2_ASAP7_75t_L g7297 ( 
.A(n_6732),
.B(n_6224),
.Y(n_7297)
);

OR2x2_ASAP7_75t_L g7298 ( 
.A(n_6681),
.B(n_6280),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6696),
.Y(n_7299)
);

AND2x4_ASAP7_75t_L g7300 ( 
.A(n_6670),
.B(n_6705),
.Y(n_7300)
);

AND2x2_ASAP7_75t_L g7301 ( 
.A(n_6745),
.B(n_6224),
.Y(n_7301)
);

AND2x2_ASAP7_75t_L g7302 ( 
.A(n_6747),
.B(n_7073),
.Y(n_7302)
);

INVx4_ASAP7_75t_L g7303 ( 
.A(n_6675),
.Y(n_7303)
);

AND2x2_ASAP7_75t_L g7304 ( 
.A(n_7073),
.B(n_6246),
.Y(n_7304)
);

AND2x2_ASAP7_75t_L g7305 ( 
.A(n_6733),
.B(n_6246),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_6787),
.B(n_6260),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_6700),
.Y(n_7307)
);

BUFx6f_ASAP7_75t_L g7308 ( 
.A(n_6707),
.Y(n_7308)
);

AND2x2_ASAP7_75t_L g7309 ( 
.A(n_6879),
.B(n_6260),
.Y(n_7309)
);

OR2x2_ASAP7_75t_L g7310 ( 
.A(n_6837),
.B(n_6713),
.Y(n_7310)
);

NOR2x1p5_ASAP7_75t_L g7311 ( 
.A(n_6707),
.B(n_7019),
.Y(n_7311)
);

INVx1_ASAP7_75t_L g7312 ( 
.A(n_6702),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_6716),
.Y(n_7313)
);

OR2x2_ASAP7_75t_L g7314 ( 
.A(n_6713),
.B(n_6280),
.Y(n_7314)
);

OR2x2_ASAP7_75t_L g7315 ( 
.A(n_6715),
.B(n_6250),
.Y(n_7315)
);

AND2x4_ASAP7_75t_L g7316 ( 
.A(n_6670),
.B(n_6705),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_6720),
.Y(n_7317)
);

HB1xp67_ASAP7_75t_L g7318 ( 
.A(n_6646),
.Y(n_7318)
);

NOR2x1_ASAP7_75t_L g7319 ( 
.A(n_6748),
.B(n_6601),
.Y(n_7319)
);

AND2x2_ASAP7_75t_L g7320 ( 
.A(n_6899),
.B(n_6271),
.Y(n_7320)
);

INVx2_ASAP7_75t_L g7321 ( 
.A(n_6811),
.Y(n_7321)
);

NAND2xp5_ASAP7_75t_L g7322 ( 
.A(n_6647),
.B(n_6508),
.Y(n_7322)
);

INVx2_ASAP7_75t_L g7323 ( 
.A(n_6811),
.Y(n_7323)
);

NOR2xp33_ASAP7_75t_L g7324 ( 
.A(n_6688),
.B(n_4884),
.Y(n_7324)
);

AND2x4_ASAP7_75t_L g7325 ( 
.A(n_6748),
.B(n_6583),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_6772),
.Y(n_7326)
);

INVxp67_ASAP7_75t_L g7327 ( 
.A(n_6650),
.Y(n_7327)
);

NAND2xp5_ASAP7_75t_L g7328 ( 
.A(n_6808),
.B(n_6513),
.Y(n_7328)
);

OR2x2_ASAP7_75t_L g7329 ( 
.A(n_6715),
.B(n_6250),
.Y(n_7329)
);

AND2x2_ASAP7_75t_L g7330 ( 
.A(n_6907),
.B(n_6271),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_6727),
.Y(n_7331)
);

AND2x2_ASAP7_75t_L g7332 ( 
.A(n_6912),
.B(n_6287),
.Y(n_7332)
);

AND2x2_ASAP7_75t_L g7333 ( 
.A(n_6897),
.B(n_6287),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_6731),
.Y(n_7334)
);

BUFx6f_ASAP7_75t_L g7335 ( 
.A(n_6707),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_6738),
.Y(n_7336)
);

INVx2_ASAP7_75t_L g7337 ( 
.A(n_6772),
.Y(n_7337)
);

NAND2xp5_ASAP7_75t_L g7338 ( 
.A(n_6808),
.B(n_6743),
.Y(n_7338)
);

AOI22xp33_ASAP7_75t_L g7339 ( 
.A1(n_6949),
.A2(n_6543),
.B1(n_6348),
.B2(n_6601),
.Y(n_7339)
);

AND2x2_ASAP7_75t_L g7340 ( 
.A(n_7014),
.B(n_6293),
.Y(n_7340)
);

HB1xp67_ASAP7_75t_L g7341 ( 
.A(n_6982),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_6744),
.Y(n_7342)
);

BUFx2_ASAP7_75t_L g7343 ( 
.A(n_6774),
.Y(n_7343)
);

AND2x2_ASAP7_75t_L g7344 ( 
.A(n_7006),
.B(n_6293),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7006),
.B(n_6295),
.Y(n_7345)
);

HB1xp67_ASAP7_75t_L g7346 ( 
.A(n_6982),
.Y(n_7346)
);

AND2x4_ASAP7_75t_L g7347 ( 
.A(n_6774),
.B(n_6583),
.Y(n_7347)
);

AND2x2_ASAP7_75t_L g7348 ( 
.A(n_6764),
.B(n_6295),
.Y(n_7348)
);

BUFx2_ASAP7_75t_SL g7349 ( 
.A(n_6944),
.Y(n_7349)
);

AND2x2_ASAP7_75t_L g7350 ( 
.A(n_6813),
.B(n_6317),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_6759),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6760),
.Y(n_7352)
);

AND2x2_ASAP7_75t_L g7353 ( 
.A(n_7018),
.B(n_6317),
.Y(n_7353)
);

AND2x2_ASAP7_75t_L g7354 ( 
.A(n_7024),
.B(n_6319),
.Y(n_7354)
);

AND2x4_ASAP7_75t_L g7355 ( 
.A(n_6772),
.B(n_6607),
.Y(n_7355)
);

INVx5_ASAP7_75t_L g7356 ( 
.A(n_6936),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_6761),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_6811),
.Y(n_7358)
);

AND2x4_ASAP7_75t_SL g7359 ( 
.A(n_7050),
.B(n_4906),
.Y(n_7359)
);

INVx1_ASAP7_75t_L g7360 ( 
.A(n_6765),
.Y(n_7360)
);

BUFx2_ASAP7_75t_L g7361 ( 
.A(n_6913),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_6781),
.Y(n_7362)
);

HB1xp67_ASAP7_75t_L g7363 ( 
.A(n_6984),
.Y(n_7363)
);

INVx2_ASAP7_75t_L g7364 ( 
.A(n_6964),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_L g7365 ( 
.A(n_6783),
.B(n_6514),
.Y(n_7365)
);

AND2x2_ASAP7_75t_L g7366 ( 
.A(n_7030),
.B(n_6319),
.Y(n_7366)
);

INVx2_ASAP7_75t_L g7367 ( 
.A(n_6964),
.Y(n_7367)
);

INVx2_ASAP7_75t_L g7368 ( 
.A(n_6986),
.Y(n_7368)
);

NAND2xp5_ASAP7_75t_L g7369 ( 
.A(n_6785),
.B(n_6515),
.Y(n_7369)
);

OR2x2_ASAP7_75t_L g7370 ( 
.A(n_6718),
.B(n_6257),
.Y(n_7370)
);

AND2x2_ASAP7_75t_L g7371 ( 
.A(n_6971),
.B(n_6418),
.Y(n_7371)
);

INVx2_ASAP7_75t_SL g7372 ( 
.A(n_6641),
.Y(n_7372)
);

INVx1_ASAP7_75t_L g7373 ( 
.A(n_6789),
.Y(n_7373)
);

AND2x2_ASAP7_75t_L g7374 ( 
.A(n_6972),
.B(n_6991),
.Y(n_7374)
);

AND2x2_ASAP7_75t_L g7375 ( 
.A(n_7001),
.B(n_6420),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6803),
.Y(n_7376)
);

AND2x2_ASAP7_75t_L g7377 ( 
.A(n_6718),
.B(n_6429),
.Y(n_7377)
);

HB1xp67_ASAP7_75t_L g7378 ( 
.A(n_6984),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_6812),
.Y(n_7379)
);

AND2x2_ASAP7_75t_L g7380 ( 
.A(n_6723),
.B(n_6429),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_6820),
.Y(n_7381)
);

INVxp67_ASAP7_75t_SL g7382 ( 
.A(n_6659),
.Y(n_7382)
);

BUFx3_ASAP7_75t_L g7383 ( 
.A(n_6995),
.Y(n_7383)
);

NAND2x1p5_ASAP7_75t_L g7384 ( 
.A(n_6997),
.B(n_5197),
.Y(n_7384)
);

HB1xp67_ASAP7_75t_L g7385 ( 
.A(n_6659),
.Y(n_7385)
);

INVx2_ASAP7_75t_L g7386 ( 
.A(n_6986),
.Y(n_7386)
);

INVx2_ASAP7_75t_L g7387 ( 
.A(n_6998),
.Y(n_7387)
);

INVx2_ASAP7_75t_L g7388 ( 
.A(n_6998),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_6821),
.B(n_6518),
.Y(n_7389)
);

NOR2xp33_ASAP7_75t_L g7390 ( 
.A(n_6831),
.B(n_7043),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_6832),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_7053),
.Y(n_7392)
);

AND2x2_ASAP7_75t_L g7393 ( 
.A(n_6723),
.B(n_6437),
.Y(n_7393)
);

NOR2xp33_ASAP7_75t_L g7394 ( 
.A(n_6624),
.B(n_4948),
.Y(n_7394)
);

NAND2x1_ASAP7_75t_L g7395 ( 
.A(n_6890),
.B(n_6382),
.Y(n_7395)
);

AND2x2_ASAP7_75t_L g7396 ( 
.A(n_6734),
.B(n_6437),
.Y(n_7396)
);

AND2x2_ASAP7_75t_L g7397 ( 
.A(n_6734),
.B(n_6455),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6833),
.Y(n_7398)
);

NOR2xp33_ASAP7_75t_L g7399 ( 
.A(n_7011),
.B(n_4948),
.Y(n_7399)
);

AND2x2_ASAP7_75t_L g7400 ( 
.A(n_6735),
.B(n_6455),
.Y(n_7400)
);

INVx2_ASAP7_75t_L g7401 ( 
.A(n_7053),
.Y(n_7401)
);

BUFx3_ASAP7_75t_L g7402 ( 
.A(n_7061),
.Y(n_7402)
);

INVx1_ASAP7_75t_SL g7403 ( 
.A(n_6943),
.Y(n_7403)
);

BUFx6f_ASAP7_75t_L g7404 ( 
.A(n_7050),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_6842),
.Y(n_7405)
);

NAND2xp5_ASAP7_75t_L g7406 ( 
.A(n_6859),
.B(n_6524),
.Y(n_7406)
);

INVx2_ASAP7_75t_L g7407 ( 
.A(n_6890),
.Y(n_7407)
);

OR2x2_ASAP7_75t_L g7408 ( 
.A(n_6735),
.B(n_6257),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_6877),
.Y(n_7409)
);

NOR2xp67_ASAP7_75t_L g7410 ( 
.A(n_6943),
.B(n_6382),
.Y(n_7410)
);

BUFx3_ASAP7_75t_L g7411 ( 
.A(n_6861),
.Y(n_7411)
);

INVx2_ASAP7_75t_L g7412 ( 
.A(n_6920),
.Y(n_7412)
);

BUFx2_ASAP7_75t_L g7413 ( 
.A(n_6967),
.Y(n_7413)
);

INVx2_ASAP7_75t_L g7414 ( 
.A(n_7010),
.Y(n_7414)
);

INVx2_ASAP7_75t_L g7415 ( 
.A(n_7010),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_6871),
.B(n_6586),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_6872),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6873),
.Y(n_7418)
);

AND2x2_ASAP7_75t_L g7419 ( 
.A(n_6741),
.B(n_6456),
.Y(n_7419)
);

OR2x2_ASAP7_75t_L g7420 ( 
.A(n_6741),
.B(n_6269),
.Y(n_7420)
);

INVx3_ASAP7_75t_L g7421 ( 
.A(n_6867),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_6874),
.B(n_6590),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6875),
.Y(n_7423)
);

HB1xp67_ASAP7_75t_L g7424 ( 
.A(n_6661),
.Y(n_7424)
);

AND2x2_ASAP7_75t_L g7425 ( 
.A(n_6753),
.B(n_6456),
.Y(n_7425)
);

AND2x2_ASAP7_75t_L g7426 ( 
.A(n_6753),
.B(n_6458),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_6882),
.Y(n_7427)
);

INVx1_ASAP7_75t_L g7428 ( 
.A(n_6891),
.Y(n_7428)
);

NAND2xp5_ASAP7_75t_L g7429 ( 
.A(n_6898),
.B(n_6527),
.Y(n_7429)
);

AND2x4_ASAP7_75t_L g7430 ( 
.A(n_6896),
.B(n_6607),
.Y(n_7430)
);

INVx1_ASAP7_75t_SL g7431 ( 
.A(n_6973),
.Y(n_7431)
);

INVx2_ASAP7_75t_L g7432 ( 
.A(n_7068),
.Y(n_7432)
);

NAND2xp5_ASAP7_75t_L g7433 ( 
.A(n_6903),
.B(n_6533),
.Y(n_7433)
);

AND2x2_ASAP7_75t_L g7434 ( 
.A(n_6762),
.B(n_6458),
.Y(n_7434)
);

AND2x4_ASAP7_75t_L g7435 ( 
.A(n_7050),
.B(n_6611),
.Y(n_7435)
);

OR2x2_ASAP7_75t_L g7436 ( 
.A(n_6762),
.B(n_6269),
.Y(n_7436)
);

INVx2_ASAP7_75t_SL g7437 ( 
.A(n_6641),
.Y(n_7437)
);

INVx3_ASAP7_75t_L g7438 ( 
.A(n_6867),
.Y(n_7438)
);

INVxp67_ASAP7_75t_L g7439 ( 
.A(n_6722),
.Y(n_7439)
);

INVx2_ASAP7_75t_L g7440 ( 
.A(n_7068),
.Y(n_7440)
);

OR2x2_ASAP7_75t_L g7441 ( 
.A(n_6763),
.B(n_6601),
.Y(n_7441)
);

AND2x2_ASAP7_75t_L g7442 ( 
.A(n_6763),
.B(n_6465),
.Y(n_7442)
);

AOI22xp33_ASAP7_75t_L g7443 ( 
.A1(n_6719),
.A2(n_7012),
.B1(n_6849),
.B2(n_6942),
.Y(n_7443)
);

AND2x4_ASAP7_75t_L g7444 ( 
.A(n_7056),
.B(n_6611),
.Y(n_7444)
);

AND2x2_ASAP7_75t_L g7445 ( 
.A(n_6755),
.B(n_6465),
.Y(n_7445)
);

INVxp67_ASAP7_75t_L g7446 ( 
.A(n_6742),
.Y(n_7446)
);

INVx2_ASAP7_75t_L g7447 ( 
.A(n_6867),
.Y(n_7447)
);

AND2x2_ASAP7_75t_L g7448 ( 
.A(n_6766),
.B(n_6468),
.Y(n_7448)
);

NAND2xp5_ASAP7_75t_L g7449 ( 
.A(n_6906),
.B(n_6541),
.Y(n_7449)
);

INVx2_ASAP7_75t_L g7450 ( 
.A(n_6884),
.Y(n_7450)
);

INVx1_ASAP7_75t_L g7451 ( 
.A(n_6914),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_6916),
.Y(n_7452)
);

AND2x2_ASAP7_75t_L g7453 ( 
.A(n_6769),
.B(n_6468),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_6918),
.Y(n_7454)
);

AND2x2_ASAP7_75t_L g7455 ( 
.A(n_6770),
.B(n_6530),
.Y(n_7455)
);

INVx2_ASAP7_75t_SL g7456 ( 
.A(n_6641),
.Y(n_7456)
);

BUFx3_ASAP7_75t_L g7457 ( 
.A(n_7056),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_6922),
.Y(n_7458)
);

AND2x2_ASAP7_75t_L g7459 ( 
.A(n_6773),
.B(n_6798),
.Y(n_7459)
);

AND2x2_ASAP7_75t_L g7460 ( 
.A(n_6798),
.B(n_6530),
.Y(n_7460)
);

NAND2xp5_ASAP7_75t_L g7461 ( 
.A(n_6924),
.B(n_6546),
.Y(n_7461)
);

AND2x4_ASAP7_75t_L g7462 ( 
.A(n_7056),
.B(n_6616),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_6930),
.Y(n_7463)
);

INVx1_ASAP7_75t_L g7464 ( 
.A(n_6934),
.Y(n_7464)
);

INVx2_ASAP7_75t_L g7465 ( 
.A(n_7070),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_6947),
.B(n_6572),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_6957),
.Y(n_7467)
);

NAND2xp5_ASAP7_75t_L g7468 ( 
.A(n_6966),
.B(n_6574),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_6970),
.Y(n_7469)
);

AND2x2_ASAP7_75t_L g7470 ( 
.A(n_6652),
.B(n_6536),
.Y(n_7470)
);

AND2x2_ASAP7_75t_L g7471 ( 
.A(n_6652),
.B(n_6536),
.Y(n_7471)
);

AND2x2_ASAP7_75t_L g7472 ( 
.A(n_6795),
.B(n_6538),
.Y(n_7472)
);

AND2x2_ASAP7_75t_L g7473 ( 
.A(n_6795),
.B(n_6538),
.Y(n_7473)
);

AND2x2_ASAP7_75t_L g7474 ( 
.A(n_6967),
.B(n_6539),
.Y(n_7474)
);

HB1xp67_ASAP7_75t_L g7475 ( 
.A(n_6661),
.Y(n_7475)
);

BUFx4f_ASAP7_75t_SL g7476 ( 
.A(n_6997),
.Y(n_7476)
);

AND2x4_ASAP7_75t_L g7477 ( 
.A(n_6994),
.B(n_6616),
.Y(n_7477)
);

AOI22xp33_ASAP7_75t_L g7478 ( 
.A1(n_7012),
.A2(n_6543),
.B1(n_6348),
.B2(n_6604),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_6978),
.Y(n_7479)
);

AND2x4_ASAP7_75t_L g7480 ( 
.A(n_6994),
.B(n_6364),
.Y(n_7480)
);

BUFx2_ASAP7_75t_L g7481 ( 
.A(n_6642),
.Y(n_7481)
);

NOR2xp33_ASAP7_75t_L g7482 ( 
.A(n_7059),
.B(n_4948),
.Y(n_7482)
);

INVxp67_ASAP7_75t_SL g7483 ( 
.A(n_6667),
.Y(n_7483)
);

NAND2xp5_ASAP7_75t_L g7484 ( 
.A(n_6988),
.B(n_6547),
.Y(n_7484)
);

HB1xp67_ASAP7_75t_L g7485 ( 
.A(n_6667),
.Y(n_7485)
);

AND2x2_ASAP7_75t_L g7486 ( 
.A(n_6927),
.B(n_6539),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_L g7487 ( 
.A(n_6990),
.B(n_6556),
.Y(n_7487)
);

BUFx2_ASAP7_75t_L g7488 ( 
.A(n_6642),
.Y(n_7488)
);

NOR2xp33_ASAP7_75t_L g7489 ( 
.A(n_6767),
.B(n_6421),
.Y(n_7489)
);

INVx3_ASAP7_75t_L g7490 ( 
.A(n_6884),
.Y(n_7490)
);

AND2x4_ASAP7_75t_L g7491 ( 
.A(n_7040),
.B(n_6364),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_6992),
.Y(n_7492)
);

INVx2_ASAP7_75t_L g7493 ( 
.A(n_7070),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_6993),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_6996),
.Y(n_7495)
);

BUFx2_ASAP7_75t_L g7496 ( 
.A(n_6642),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7000),
.Y(n_7497)
);

AND2x4_ASAP7_75t_L g7498 ( 
.A(n_7040),
.B(n_6604),
.Y(n_7498)
);

AND2x2_ASAP7_75t_SL g7499 ( 
.A(n_6757),
.B(n_5555),
.Y(n_7499)
);

INVx2_ASAP7_75t_L g7500 ( 
.A(n_6884),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_7003),
.Y(n_7501)
);

AND2x2_ASAP7_75t_L g7502 ( 
.A(n_6932),
.B(n_6390),
.Y(n_7502)
);

AND2x4_ASAP7_75t_L g7503 ( 
.A(n_6691),
.B(n_6938),
.Y(n_7503)
);

HB1xp67_ASAP7_75t_L g7504 ( 
.A(n_6802),
.Y(n_7504)
);

BUFx2_ASAP7_75t_L g7505 ( 
.A(n_6691),
.Y(n_7505)
);

NOR2x1_ASAP7_75t_L g7506 ( 
.A(n_6997),
.B(n_6604),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_6909),
.Y(n_7507)
);

BUFx2_ASAP7_75t_L g7508 ( 
.A(n_6691),
.Y(n_7508)
);

INVx2_ASAP7_75t_L g7509 ( 
.A(n_6909),
.Y(n_7509)
);

INVx1_ASAP7_75t_L g7510 ( 
.A(n_7007),
.Y(n_7510)
);

HB1xp67_ASAP7_75t_L g7511 ( 
.A(n_6802),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_7115),
.Y(n_7512)
);

BUFx2_ASAP7_75t_L g7513 ( 
.A(n_7135),
.Y(n_7513)
);

INVx2_ASAP7_75t_L g7514 ( 
.A(n_7135),
.Y(n_7514)
);

OR2x6_ASAP7_75t_L g7515 ( 
.A(n_7349),
.B(n_6543),
.Y(n_7515)
);

NAND2xp5_ASAP7_75t_L g7516 ( 
.A(n_7143),
.B(n_6757),
.Y(n_7516)
);

AOI21xp33_ASAP7_75t_L g7517 ( 
.A1(n_7154),
.A2(n_7037),
.B(n_6953),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7115),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_7143),
.B(n_6758),
.Y(n_7519)
);

INVx2_ASAP7_75t_L g7520 ( 
.A(n_7222),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7125),
.Y(n_7521)
);

OR2x2_ASAP7_75t_L g7522 ( 
.A(n_7088),
.B(n_6660),
.Y(n_7522)
);

BUFx3_ASAP7_75t_L g7523 ( 
.A(n_7236),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_7125),
.Y(n_7524)
);

OR2x6_ASAP7_75t_L g7525 ( 
.A(n_7222),
.B(n_4790),
.Y(n_7525)
);

AND2x2_ASAP7_75t_L g7526 ( 
.A(n_7132),
.B(n_6941),
.Y(n_7526)
);

INVxp67_ASAP7_75t_SL g7527 ( 
.A(n_7131),
.Y(n_7527)
);

AOI21xp5_ASAP7_75t_L g7528 ( 
.A1(n_7154),
.A2(n_7080),
.B(n_7499),
.Y(n_7528)
);

INVxp67_ASAP7_75t_SL g7529 ( 
.A(n_7131),
.Y(n_7529)
);

AND2x2_ASAP7_75t_L g7530 ( 
.A(n_7136),
.B(n_6851),
.Y(n_7530)
);

OR2x2_ASAP7_75t_L g7531 ( 
.A(n_7077),
.B(n_6695),
.Y(n_7531)
);

NAND2xp5_ASAP7_75t_SL g7532 ( 
.A(n_7356),
.B(n_7066),
.Y(n_7532)
);

NOR2xp67_ASAP7_75t_L g7533 ( 
.A(n_7356),
.B(n_6411),
.Y(n_7533)
);

NAND4xp25_ASAP7_75t_L g7534 ( 
.A(n_7443),
.B(n_7037),
.C(n_6838),
.D(n_6953),
.Y(n_7534)
);

INVx4_ASAP7_75t_L g7535 ( 
.A(n_7308),
.Y(n_7535)
);

INVx2_ASAP7_75t_L g7536 ( 
.A(n_7109),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7168),
.Y(n_7537)
);

INVx1_ASAP7_75t_L g7538 ( 
.A(n_7168),
.Y(n_7538)
);

OAI21x1_ASAP7_75t_L g7539 ( 
.A1(n_7395),
.A2(n_6664),
.B(n_6958),
.Y(n_7539)
);

BUFx3_ASAP7_75t_L g7540 ( 
.A(n_7295),
.Y(n_7540)
);

A2O1A1Ixp33_ASAP7_75t_L g7541 ( 
.A1(n_7443),
.A2(n_7089),
.B(n_7212),
.C(n_7394),
.Y(n_7541)
);

OAI21x1_ASAP7_75t_L g7542 ( 
.A1(n_7090),
.A2(n_6976),
.B(n_6819),
.Y(n_7542)
);

INVx2_ASAP7_75t_SL g7543 ( 
.A(n_7213),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7177),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7177),
.Y(n_7545)
);

AOI21xp5_ASAP7_75t_L g7546 ( 
.A1(n_7080),
.A2(n_6644),
.B(n_6881),
.Y(n_7546)
);

NAND2xp5_ASAP7_75t_L g7547 ( 
.A(n_7361),
.B(n_6768),
.Y(n_7547)
);

AND2x2_ASAP7_75t_L g7548 ( 
.A(n_7251),
.B(n_7245),
.Y(n_7548)
);

OAI21x1_ASAP7_75t_L g7549 ( 
.A1(n_7090),
.A2(n_7296),
.B(n_7506),
.Y(n_7549)
);

INVx2_ASAP7_75t_SL g7550 ( 
.A(n_7213),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7181),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7181),
.Y(n_7552)
);

BUFx3_ASAP7_75t_L g7553 ( 
.A(n_7295),
.Y(n_7553)
);

OAI21x1_ASAP7_75t_L g7554 ( 
.A1(n_7296),
.A2(n_7033),
.B(n_6819),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_L g7555 ( 
.A(n_7211),
.B(n_6698),
.Y(n_7555)
);

INVxp67_ASAP7_75t_L g7556 ( 
.A(n_7413),
.Y(n_7556)
);

AND2x2_ASAP7_75t_L g7557 ( 
.A(n_7145),
.B(n_6945),
.Y(n_7557)
);

INVxp67_ASAP7_75t_L g7558 ( 
.A(n_7092),
.Y(n_7558)
);

AND2x2_ASAP7_75t_L g7559 ( 
.A(n_7122),
.B(n_6959),
.Y(n_7559)
);

OAI21xp5_ASAP7_75t_L g7560 ( 
.A1(n_7499),
.A2(n_6717),
.B(n_6712),
.Y(n_7560)
);

INVx2_ASAP7_75t_L g7561 ( 
.A(n_7109),
.Y(n_7561)
);

AND2x2_ASAP7_75t_L g7562 ( 
.A(n_7101),
.B(n_6862),
.Y(n_7562)
);

INVx2_ASAP7_75t_L g7563 ( 
.A(n_7130),
.Y(n_7563)
);

AND2x2_ASAP7_75t_L g7564 ( 
.A(n_7127),
.B(n_7039),
.Y(n_7564)
);

A2O1A1Ixp33_ASAP7_75t_L g7565 ( 
.A1(n_7212),
.A2(n_7394),
.B(n_7410),
.C(n_7267),
.Y(n_7565)
);

NAND2xp5_ASAP7_75t_L g7566 ( 
.A(n_7211),
.B(n_6805),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_7204),
.Y(n_7567)
);

INVxp67_ASAP7_75t_L g7568 ( 
.A(n_7343),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_7204),
.Y(n_7569)
);

AND2x2_ASAP7_75t_L g7570 ( 
.A(n_7128),
.B(n_7057),
.Y(n_7570)
);

O2A1O1Ixp5_ASAP7_75t_L g7571 ( 
.A1(n_7247),
.A2(n_6622),
.B(n_6730),
.C(n_6724),
.Y(n_7571)
);

OR2x2_ASAP7_75t_L g7572 ( 
.A(n_7107),
.B(n_7248),
.Y(n_7572)
);

AND2x2_ASAP7_75t_L g7573 ( 
.A(n_7265),
.B(n_6962),
.Y(n_7573)
);

O2A1O1Ixp5_ASAP7_75t_L g7574 ( 
.A1(n_7247),
.A2(n_7218),
.B(n_7193),
.C(n_7182),
.Y(n_7574)
);

AND2x2_ASAP7_75t_L g7575 ( 
.A(n_7271),
.B(n_6965),
.Y(n_7575)
);

HB1xp67_ASAP7_75t_L g7576 ( 
.A(n_7220),
.Y(n_7576)
);

OR2x2_ASAP7_75t_L g7577 ( 
.A(n_7248),
.B(n_6929),
.Y(n_7577)
);

NOR2xp33_ASAP7_75t_R g7578 ( 
.A(n_7291),
.B(n_4790),
.Y(n_7578)
);

INVx2_ASAP7_75t_L g7579 ( 
.A(n_7130),
.Y(n_7579)
);

AOI21xp5_ASAP7_75t_L g7580 ( 
.A1(n_7214),
.A2(n_6717),
.B(n_6712),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7220),
.Y(n_7581)
);

BUFx3_ASAP7_75t_L g7582 ( 
.A(n_7098),
.Y(n_7582)
);

A2O1A1Ixp33_ASAP7_75t_L g7583 ( 
.A1(n_7267),
.A2(n_7066),
.B(n_6951),
.C(n_6835),
.Y(n_7583)
);

OAI21xp33_ASAP7_75t_L g7584 ( 
.A1(n_7254),
.A2(n_6671),
.B(n_6655),
.Y(n_7584)
);

INVx1_ASAP7_75t_SL g7585 ( 
.A(n_7103),
.Y(n_7585)
);

INVx3_ASAP7_75t_L g7586 ( 
.A(n_7308),
.Y(n_7586)
);

OAI21xp5_ASAP7_75t_L g7587 ( 
.A1(n_7254),
.A2(n_7049),
.B(n_6730),
.Y(n_7587)
);

NOR2xp33_ASAP7_75t_L g7588 ( 
.A(n_7303),
.B(n_5753),
.Y(n_7588)
);

INVxp67_ASAP7_75t_L g7589 ( 
.A(n_7390),
.Y(n_7589)
);

AOI21xp5_ASAP7_75t_L g7590 ( 
.A1(n_7214),
.A2(n_6724),
.B(n_6895),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7239),
.Y(n_7591)
);

CKINVDCx5p33_ASAP7_75t_R g7592 ( 
.A(n_7324),
.Y(n_7592)
);

OA21x2_ASAP7_75t_L g7593 ( 
.A1(n_7193),
.A2(n_6699),
.B(n_6686),
.Y(n_7593)
);

NAND2xp5_ASAP7_75t_L g7594 ( 
.A(n_7383),
.B(n_6806),
.Y(n_7594)
);

AOI21xp5_ASAP7_75t_L g7595 ( 
.A1(n_7218),
.A2(n_6925),
.B(n_6604),
.Y(n_7595)
);

NAND3xp33_ASAP7_75t_L g7596 ( 
.A(n_7356),
.B(n_6804),
.C(n_6814),
.Y(n_7596)
);

NAND2xp5_ASAP7_75t_L g7597 ( 
.A(n_7383),
.B(n_6836),
.Y(n_7597)
);

AOI221xp5_ASAP7_75t_L g7598 ( 
.A1(n_7403),
.A2(n_6829),
.B1(n_6854),
.B2(n_6824),
.C(n_6818),
.Y(n_7598)
);

NAND4xp25_ASAP7_75t_L g7599 ( 
.A(n_7339),
.B(n_5835),
.C(n_5902),
.D(n_5851),
.Y(n_7599)
);

INVxp67_ASAP7_75t_L g7600 ( 
.A(n_7390),
.Y(n_7600)
);

AND2x2_ASAP7_75t_L g7601 ( 
.A(n_7291),
.B(n_7064),
.Y(n_7601)
);

HB1xp67_ASAP7_75t_L g7602 ( 
.A(n_7239),
.Y(n_7602)
);

INVx2_ASAP7_75t_L g7603 ( 
.A(n_7144),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_7253),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_L g7605 ( 
.A(n_7402),
.B(n_6843),
.Y(n_7605)
);

INVx2_ASAP7_75t_L g7606 ( 
.A(n_7144),
.Y(n_7606)
);

INVx2_ASAP7_75t_L g7607 ( 
.A(n_7144),
.Y(n_7607)
);

INVx1_ASAP7_75t_SL g7608 ( 
.A(n_7098),
.Y(n_7608)
);

OA21x2_ASAP7_75t_L g7609 ( 
.A1(n_7083),
.A2(n_6699),
.B(n_6686),
.Y(n_7609)
);

AND2x2_ASAP7_75t_L g7610 ( 
.A(n_7155),
.B(n_7459),
.Y(n_7610)
);

OR2x6_ASAP7_75t_L g7611 ( 
.A(n_7303),
.B(n_4861),
.Y(n_7611)
);

AO21x2_ASAP7_75t_L g7612 ( 
.A1(n_7083),
.A2(n_6788),
.B(n_6779),
.Y(n_7612)
);

AND2x2_ASAP7_75t_L g7613 ( 
.A(n_7470),
.B(n_7067),
.Y(n_7613)
);

INVx2_ASAP7_75t_L g7614 ( 
.A(n_7213),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7253),
.Y(n_7615)
);

NAND2x1_ASAP7_75t_L g7616 ( 
.A(n_7319),
.B(n_6909),
.Y(n_7616)
);

INVx2_ASAP7_75t_L g7617 ( 
.A(n_7213),
.Y(n_7617)
);

AOI21x1_ASAP7_75t_L g7618 ( 
.A1(n_7341),
.A2(n_6788),
.B(n_6779),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7258),
.Y(n_7619)
);

INVx1_ASAP7_75t_L g7620 ( 
.A(n_7258),
.Y(n_7620)
);

NAND2xp5_ASAP7_75t_L g7621 ( 
.A(n_7402),
.B(n_7021),
.Y(n_7621)
);

OR2x2_ASAP7_75t_L g7622 ( 
.A(n_7124),
.B(n_6985),
.Y(n_7622)
);

INVx1_ASAP7_75t_L g7623 ( 
.A(n_7263),
.Y(n_7623)
);

AOI21x1_ASAP7_75t_L g7624 ( 
.A1(n_7341),
.A2(n_6793),
.B(n_6794),
.Y(n_7624)
);

AND2x2_ASAP7_75t_L g7625 ( 
.A(n_7471),
.B(n_7028),
.Y(n_7625)
);

INVx2_ASAP7_75t_L g7626 ( 
.A(n_7421),
.Y(n_7626)
);

OAI21xp5_ASAP7_75t_L g7627 ( 
.A1(n_7118),
.A2(n_6145),
.B(n_6093),
.Y(n_7627)
);

INVx4_ASAP7_75t_L g7628 ( 
.A(n_7308),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7263),
.Y(n_7629)
);

NAND2xp5_ASAP7_75t_L g7630 ( 
.A(n_7300),
.B(n_7009),
.Y(n_7630)
);

NAND2x1_ASAP7_75t_L g7631 ( 
.A(n_7240),
.B(n_6911),
.Y(n_7631)
);

INVx3_ASAP7_75t_L g7632 ( 
.A(n_7308),
.Y(n_7632)
);

AOI21xp5_ASAP7_75t_L g7633 ( 
.A1(n_7324),
.A2(n_6908),
.B(n_6883),
.Y(n_7633)
);

OR2x6_ASAP7_75t_L g7634 ( 
.A(n_7288),
.B(n_4861),
.Y(n_7634)
);

INVx2_ASAP7_75t_L g7635 ( 
.A(n_7421),
.Y(n_7635)
);

NAND2xp5_ASAP7_75t_L g7636 ( 
.A(n_7300),
.B(n_6940),
.Y(n_7636)
);

AO21x1_ASAP7_75t_L g7637 ( 
.A1(n_7100),
.A2(n_6908),
.B(n_6883),
.Y(n_7637)
);

AND2x2_ASAP7_75t_L g7638 ( 
.A(n_7474),
.B(n_6904),
.Y(n_7638)
);

AND2x4_ASAP7_75t_L g7639 ( 
.A(n_7316),
.B(n_6911),
.Y(n_7639)
);

AND2x2_ASAP7_75t_L g7640 ( 
.A(n_7260),
.B(n_6910),
.Y(n_7640)
);

HB1xp67_ASAP7_75t_L g7641 ( 
.A(n_7504),
.Y(n_7641)
);

AND2x2_ASAP7_75t_L g7642 ( 
.A(n_7302),
.B(n_6921),
.Y(n_7642)
);

INVx2_ASAP7_75t_L g7643 ( 
.A(n_7438),
.Y(n_7643)
);

INVx1_ASAP7_75t_SL g7644 ( 
.A(n_7316),
.Y(n_7644)
);

AOI21xp5_ASAP7_75t_L g7645 ( 
.A1(n_7178),
.A2(n_6014),
.B(n_6093),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7273),
.Y(n_7646)
);

BUFx3_ASAP7_75t_L g7647 ( 
.A(n_7162),
.Y(n_7647)
);

BUFx3_ASAP7_75t_L g7648 ( 
.A(n_7162),
.Y(n_7648)
);

INVx1_ASAP7_75t_SL g7649 ( 
.A(n_7476),
.Y(n_7649)
);

OAI21xp33_ASAP7_75t_L g7650 ( 
.A1(n_7309),
.A2(n_6954),
.B(n_6894),
.Y(n_7650)
);

O2A1O1Ixp33_ASAP7_75t_L g7651 ( 
.A1(n_7327),
.A2(n_6900),
.B(n_6905),
.C(n_6893),
.Y(n_7651)
);

BUFx3_ASAP7_75t_L g7652 ( 
.A(n_7182),
.Y(n_7652)
);

BUFx2_ASAP7_75t_L g7653 ( 
.A(n_7438),
.Y(n_7653)
);

INVx1_ASAP7_75t_L g7654 ( 
.A(n_7273),
.Y(n_7654)
);

NAND2xp5_ASAP7_75t_L g7655 ( 
.A(n_7120),
.B(n_7013),
.Y(n_7655)
);

AND2x4_ASAP7_75t_L g7656 ( 
.A(n_7356),
.B(n_6911),
.Y(n_7656)
);

INVx2_ASAP7_75t_SL g7657 ( 
.A(n_7311),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7293),
.Y(n_7658)
);

INVx2_ASAP7_75t_L g7659 ( 
.A(n_7490),
.Y(n_7659)
);

NAND3xp33_ASAP7_75t_L g7660 ( 
.A(n_7478),
.B(n_7150),
.C(n_7199),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_7293),
.Y(n_7661)
);

AND2x2_ASAP7_75t_L g7662 ( 
.A(n_7084),
.B(n_6961),
.Y(n_7662)
);

OAI21xp33_ASAP7_75t_L g7663 ( 
.A1(n_7320),
.A2(n_7017),
.B(n_7015),
.Y(n_7663)
);

INVx2_ASAP7_75t_L g7664 ( 
.A(n_7490),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7318),
.Y(n_7665)
);

HB1xp67_ASAP7_75t_L g7666 ( 
.A(n_7504),
.Y(n_7666)
);

BUFx2_ASAP7_75t_L g7667 ( 
.A(n_7241),
.Y(n_7667)
);

HB1xp67_ASAP7_75t_L g7668 ( 
.A(n_7511),
.Y(n_7668)
);

NAND2x1_ASAP7_75t_L g7669 ( 
.A(n_7355),
.B(n_6950),
.Y(n_7669)
);

INVx2_ASAP7_75t_L g7670 ( 
.A(n_7335),
.Y(n_7670)
);

OR2x6_ASAP7_75t_L g7671 ( 
.A(n_7199),
.B(n_4861),
.Y(n_7671)
);

INVx2_ASAP7_75t_L g7672 ( 
.A(n_7335),
.Y(n_7672)
);

INVx1_ASAP7_75t_SL g7673 ( 
.A(n_7476),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_7318),
.Y(n_7674)
);

OA21x2_ASAP7_75t_L g7675 ( 
.A1(n_7100),
.A2(n_6709),
.B(n_6793),
.Y(n_7675)
);

INVx2_ASAP7_75t_L g7676 ( 
.A(n_7335),
.Y(n_7676)
);

BUFx6f_ASAP7_75t_L g7677 ( 
.A(n_7335),
.Y(n_7677)
);

AOI21xp33_ASAP7_75t_L g7678 ( 
.A1(n_7399),
.A2(n_6825),
.B(n_6810),
.Y(n_7678)
);

AND2x2_ASAP7_75t_L g7679 ( 
.A(n_7085),
.B(n_7305),
.Y(n_7679)
);

AND2x4_ASAP7_75t_L g7680 ( 
.A(n_7241),
.B(n_6810),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_7511),
.Y(n_7681)
);

AOI21xp5_ASAP7_75t_L g7682 ( 
.A1(n_7192),
.A2(n_6145),
.B(n_4772),
.Y(n_7682)
);

BUFx3_ASAP7_75t_L g7683 ( 
.A(n_7200),
.Y(n_7683)
);

INVx2_ASAP7_75t_L g7684 ( 
.A(n_7081),
.Y(n_7684)
);

A2O1A1Ixp33_ASAP7_75t_L g7685 ( 
.A1(n_7118),
.A2(n_7033),
.B(n_6226),
.C(n_6228),
.Y(n_7685)
);

AOI21xp5_ASAP7_75t_L g7686 ( 
.A1(n_7399),
.A2(n_7489),
.B(n_7478),
.Y(n_7686)
);

NOR2x1p5_ASAP7_75t_L g7687 ( 
.A(n_7411),
.B(n_5114),
.Y(n_7687)
);

NAND2xp5_ASAP7_75t_L g7688 ( 
.A(n_7134),
.B(n_7022),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_7075),
.Y(n_7689)
);

BUFx6f_ASAP7_75t_L g7690 ( 
.A(n_7081),
.Y(n_7690)
);

HB1xp67_ASAP7_75t_L g7691 ( 
.A(n_7081),
.Y(n_7691)
);

OAI21xp5_ASAP7_75t_L g7692 ( 
.A1(n_7339),
.A2(n_6449),
.B(n_6411),
.Y(n_7692)
);

OAI21x1_ASAP7_75t_L g7693 ( 
.A1(n_7384),
.A2(n_7025),
.B(n_6960),
.Y(n_7693)
);

BUFx3_ASAP7_75t_L g7694 ( 
.A(n_7210),
.Y(n_7694)
);

OR2x2_ASAP7_75t_L g7695 ( 
.A(n_7310),
.B(n_7225),
.Y(n_7695)
);

AND2x2_ASAP7_75t_L g7696 ( 
.A(n_7306),
.B(n_6961),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7079),
.Y(n_7697)
);

INVxp33_ASAP7_75t_L g7698 ( 
.A(n_7482),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7093),
.Y(n_7699)
);

INVx2_ASAP7_75t_L g7700 ( 
.A(n_7081),
.Y(n_7700)
);

INVx2_ASAP7_75t_L g7701 ( 
.A(n_7113),
.Y(n_7701)
);

AND2x2_ASAP7_75t_L g7702 ( 
.A(n_7472),
.B(n_6330),
.Y(n_7702)
);

AOI21xp33_ASAP7_75t_L g7703 ( 
.A1(n_7489),
.A2(n_6827),
.B(n_6825),
.Y(n_7703)
);

OAI21x1_ASAP7_75t_L g7704 ( 
.A1(n_7384),
.A2(n_6960),
.B(n_6950),
.Y(n_7704)
);

OAI21xp5_ASAP7_75t_SL g7705 ( 
.A1(n_7359),
.A2(n_5164),
.B(n_5382),
.Y(n_7705)
);

INVx1_ASAP7_75t_L g7706 ( 
.A(n_7104),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7111),
.Y(n_7707)
);

AOI21xp5_ASAP7_75t_L g7708 ( 
.A1(n_7482),
.A2(n_7035),
.B(n_7032),
.Y(n_7708)
);

AND2x2_ASAP7_75t_L g7709 ( 
.A(n_7473),
.B(n_7330),
.Y(n_7709)
);

INVx2_ASAP7_75t_L g7710 ( 
.A(n_7113),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7129),
.Y(n_7711)
);

HB1xp67_ASAP7_75t_L g7712 ( 
.A(n_7113),
.Y(n_7712)
);

NAND2xp5_ASAP7_75t_L g7713 ( 
.A(n_7137),
.B(n_7041),
.Y(n_7713)
);

INVx1_ASAP7_75t_SL g7714 ( 
.A(n_7481),
.Y(n_7714)
);

INVx2_ASAP7_75t_SL g7715 ( 
.A(n_7113),
.Y(n_7715)
);

AO21x2_ASAP7_75t_L g7716 ( 
.A1(n_7123),
.A2(n_6796),
.B(n_6794),
.Y(n_7716)
);

NAND2xp5_ASAP7_75t_L g7717 ( 
.A(n_7138),
.B(n_7046),
.Y(n_7717)
);

INVx1_ASAP7_75t_L g7718 ( 
.A(n_7123),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_7346),
.Y(n_7719)
);

NAND2xp5_ASAP7_75t_L g7720 ( 
.A(n_7142),
.B(n_7047),
.Y(n_7720)
);

INVxp67_ASAP7_75t_SL g7721 ( 
.A(n_7191),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_7346),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_7363),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7363),
.Y(n_7724)
);

INVx2_ASAP7_75t_L g7725 ( 
.A(n_7191),
.Y(n_7725)
);

INVx2_ASAP7_75t_L g7726 ( 
.A(n_7191),
.Y(n_7726)
);

NAND2xp33_ASAP7_75t_L g7727 ( 
.A(n_7404),
.B(n_5574),
.Y(n_7727)
);

AND2x2_ASAP7_75t_L g7728 ( 
.A(n_7332),
.B(n_6362),
.Y(n_7728)
);

INVx1_ASAP7_75t_SL g7729 ( 
.A(n_7488),
.Y(n_7729)
);

AOI21xp5_ASAP7_75t_L g7730 ( 
.A1(n_7096),
.A2(n_7055),
.B(n_7051),
.Y(n_7730)
);

HB1xp67_ASAP7_75t_L g7731 ( 
.A(n_7191),
.Y(n_7731)
);

INVx2_ASAP7_75t_L g7732 ( 
.A(n_7229),
.Y(n_7732)
);

INVx1_ASAP7_75t_L g7733 ( 
.A(n_7378),
.Y(n_7733)
);

OA21x2_ASAP7_75t_L g7734 ( 
.A1(n_7269),
.A2(n_6709),
.B(n_6676),
.Y(n_7734)
);

AO22x2_ASAP7_75t_L g7735 ( 
.A1(n_7133),
.A2(n_6676),
.B1(n_6684),
.B2(n_6673),
.Y(n_7735)
);

INVx2_ASAP7_75t_L g7736 ( 
.A(n_7229),
.Y(n_7736)
);

AOI21xp5_ASAP7_75t_L g7737 ( 
.A1(n_7096),
.A2(n_7065),
.B(n_7058),
.Y(n_7737)
);

INVx1_ASAP7_75t_SL g7738 ( 
.A(n_7496),
.Y(n_7738)
);

OR2x2_ASAP7_75t_L g7739 ( 
.A(n_7223),
.B(n_6968),
.Y(n_7739)
);

AND2x2_ASAP7_75t_L g7740 ( 
.A(n_7243),
.B(n_6362),
.Y(n_7740)
);

AOI21x1_ASAP7_75t_L g7741 ( 
.A1(n_7378),
.A2(n_6799),
.B(n_6796),
.Y(n_7741)
);

INVx2_ASAP7_75t_L g7742 ( 
.A(n_7229),
.Y(n_7742)
);

AND2x4_ASAP7_75t_SL g7743 ( 
.A(n_7087),
.B(n_4879),
.Y(n_7743)
);

NOR2xp33_ASAP7_75t_R g7744 ( 
.A(n_7140),
.B(n_5096),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7139),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_7147),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_7148),
.Y(n_7747)
);

A2O1A1Ixp33_ASAP7_75t_L g7748 ( 
.A1(n_7359),
.A2(n_6226),
.B(n_6228),
.C(n_6411),
.Y(n_7748)
);

INVx1_ASAP7_75t_SL g7749 ( 
.A(n_7505),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7152),
.Y(n_7750)
);

OR2x6_ASAP7_75t_L g7751 ( 
.A(n_7082),
.B(n_3736),
.Y(n_7751)
);

NAND2xp5_ASAP7_75t_SL g7752 ( 
.A(n_7404),
.B(n_6449),
.Y(n_7752)
);

AO21x2_ASAP7_75t_L g7753 ( 
.A1(n_7269),
.A2(n_6799),
.B(n_6684),
.Y(n_7753)
);

OR2x2_ASAP7_75t_L g7754 ( 
.A(n_7194),
.B(n_7008),
.Y(n_7754)
);

AND2x2_ASAP7_75t_L g7755 ( 
.A(n_7246),
.B(n_6339),
.Y(n_7755)
);

INVx1_ASAP7_75t_L g7756 ( 
.A(n_7153),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_L g7757 ( 
.A(n_7149),
.B(n_7237),
.Y(n_7757)
);

AOI21xp5_ASAP7_75t_L g7758 ( 
.A1(n_7106),
.A2(n_6828),
.B(n_6827),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7156),
.Y(n_7759)
);

INVx2_ASAP7_75t_SL g7760 ( 
.A(n_7229),
.Y(n_7760)
);

INVx2_ASAP7_75t_L g7761 ( 
.A(n_7404),
.Y(n_7761)
);

OAI21x1_ASAP7_75t_L g7762 ( 
.A1(n_7078),
.A2(n_6960),
.B(n_6950),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_7159),
.Y(n_7763)
);

NAND2xp5_ASAP7_75t_L g7764 ( 
.A(n_7078),
.B(n_6878),
.Y(n_7764)
);

HB1xp67_ASAP7_75t_L g7765 ( 
.A(n_7508),
.Y(n_7765)
);

INVx2_ASAP7_75t_L g7766 ( 
.A(n_7404),
.Y(n_7766)
);

CKINVDCx14_ASAP7_75t_R g7767 ( 
.A(n_7146),
.Y(n_7767)
);

INVx2_ASAP7_75t_L g7768 ( 
.A(n_7086),
.Y(n_7768)
);

OAI21xp5_ASAP7_75t_L g7769 ( 
.A1(n_7439),
.A2(n_6481),
.B(n_6449),
.Y(n_7769)
);

OAI21xp33_ASAP7_75t_L g7770 ( 
.A1(n_7431),
.A2(n_6870),
.B(n_7052),
.Y(n_7770)
);

INVx2_ASAP7_75t_L g7771 ( 
.A(n_7086),
.Y(n_7771)
);

AND2x2_ASAP7_75t_L g7772 ( 
.A(n_7445),
.B(n_6339),
.Y(n_7772)
);

AND2x4_ASAP7_75t_L g7773 ( 
.A(n_7234),
.B(n_6828),
.Y(n_7773)
);

INVx2_ASAP7_75t_SL g7774 ( 
.A(n_7169),
.Y(n_7774)
);

NAND2x1_ASAP7_75t_L g7775 ( 
.A(n_7355),
.B(n_7025),
.Y(n_7775)
);

OAI21xp5_ASAP7_75t_L g7776 ( 
.A1(n_7439),
.A2(n_6496),
.B(n_6481),
.Y(n_7776)
);

NAND3xp33_ASAP7_75t_SL g7777 ( 
.A(n_7167),
.B(n_5793),
.C(n_5124),
.Y(n_7777)
);

OA21x2_ASAP7_75t_L g7778 ( 
.A1(n_7382),
.A2(n_6673),
.B(n_7036),
.Y(n_7778)
);

INVx2_ASAP7_75t_L g7779 ( 
.A(n_7457),
.Y(n_7779)
);

CKINVDCx5p33_ASAP7_75t_R g7780 ( 
.A(n_7457),
.Y(n_7780)
);

INVx1_ASAP7_75t_L g7781 ( 
.A(n_7164),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7171),
.Y(n_7782)
);

INVx1_ASAP7_75t_L g7783 ( 
.A(n_7172),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_7175),
.Y(n_7784)
);

INVx4_ASAP7_75t_SL g7785 ( 
.A(n_7119),
.Y(n_7785)
);

INVx2_ASAP7_75t_L g7786 ( 
.A(n_7163),
.Y(n_7786)
);

INVx2_ASAP7_75t_L g7787 ( 
.A(n_7163),
.Y(n_7787)
);

OAI21x1_ASAP7_75t_L g7788 ( 
.A1(n_7407),
.A2(n_7042),
.B(n_7025),
.Y(n_7788)
);

INVx5_ASAP7_75t_L g7789 ( 
.A(n_7119),
.Y(n_7789)
);

HB1xp67_ASAP7_75t_L g7790 ( 
.A(n_7364),
.Y(n_7790)
);

OA21x2_ASAP7_75t_L g7791 ( 
.A1(n_7382),
.A2(n_7044),
.B(n_7036),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_7385),
.Y(n_7792)
);

INVx2_ASAP7_75t_L g7793 ( 
.A(n_7166),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_7385),
.Y(n_7794)
);

NOR2xp33_ASAP7_75t_L g7795 ( 
.A(n_7446),
.B(n_5180),
.Y(n_7795)
);

BUFx2_ASAP7_75t_L g7796 ( 
.A(n_7169),
.Y(n_7796)
);

NAND2xp5_ASAP7_75t_L g7797 ( 
.A(n_7227),
.B(n_6844),
.Y(n_7797)
);

AO21x2_ASAP7_75t_L g7798 ( 
.A1(n_7483),
.A2(n_7045),
.B(n_7044),
.Y(n_7798)
);

INVx2_ASAP7_75t_L g7799 ( 
.A(n_7166),
.Y(n_7799)
);

NAND4xp25_ASAP7_75t_L g7800 ( 
.A(n_7411),
.B(n_7071),
.C(n_7042),
.D(n_6845),
.Y(n_7800)
);

BUFx3_ASAP7_75t_L g7801 ( 
.A(n_7157),
.Y(n_7801)
);

A2O1A1Ixp33_ASAP7_75t_L g7802 ( 
.A1(n_7446),
.A2(n_6496),
.B(n_6481),
.C(n_6466),
.Y(n_7802)
);

BUFx2_ASAP7_75t_L g7803 ( 
.A(n_7198),
.Y(n_7803)
);

INVx2_ASAP7_75t_L g7804 ( 
.A(n_7184),
.Y(n_7804)
);

INVx2_ASAP7_75t_L g7805 ( 
.A(n_7184),
.Y(n_7805)
);

A2O1A1Ixp33_ASAP7_75t_L g7806 ( 
.A1(n_7180),
.A2(n_7187),
.B(n_7196),
.C(n_7185),
.Y(n_7806)
);

AOI21xp5_ASAP7_75t_L g7807 ( 
.A1(n_7106),
.A2(n_6845),
.B(n_6844),
.Y(n_7807)
);

INVx1_ASAP7_75t_L g7808 ( 
.A(n_7424),
.Y(n_7808)
);

AOI21xp5_ASAP7_75t_L g7809 ( 
.A1(n_7110),
.A2(n_6850),
.B(n_6848),
.Y(n_7809)
);

NAND2xp5_ASAP7_75t_L g7810 ( 
.A(n_7230),
.B(n_6850),
.Y(n_7810)
);

INVx1_ASAP7_75t_L g7811 ( 
.A(n_7424),
.Y(n_7811)
);

INVx4_ASAP7_75t_SL g7812 ( 
.A(n_7157),
.Y(n_7812)
);

INVx1_ASAP7_75t_L g7813 ( 
.A(n_7475),
.Y(n_7813)
);

INVx2_ASAP7_75t_SL g7814 ( 
.A(n_7198),
.Y(n_7814)
);

AOI21xp5_ASAP7_75t_L g7815 ( 
.A1(n_7110),
.A2(n_6853),
.B(n_6848),
.Y(n_7815)
);

INVx3_ASAP7_75t_L g7816 ( 
.A(n_7325),
.Y(n_7816)
);

O2A1O1Ixp33_ASAP7_75t_L g7817 ( 
.A1(n_7327),
.A2(n_6900),
.B(n_6905),
.C(n_6893),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7475),
.Y(n_7818)
);

HB1xp67_ASAP7_75t_L g7819 ( 
.A(n_7364),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_7485),
.Y(n_7820)
);

INVx1_ASAP7_75t_L g7821 ( 
.A(n_7485),
.Y(n_7821)
);

INVx4_ASAP7_75t_L g7822 ( 
.A(n_7367),
.Y(n_7822)
);

HB1xp67_ASAP7_75t_L g7823 ( 
.A(n_7367),
.Y(n_7823)
);

HB1xp67_ASAP7_75t_L g7824 ( 
.A(n_7368),
.Y(n_7824)
);

INVx2_ASAP7_75t_L g7825 ( 
.A(n_7188),
.Y(n_7825)
);

NOR2xp33_ASAP7_75t_L g7826 ( 
.A(n_7105),
.B(n_4879),
.Y(n_7826)
);

INVx2_ASAP7_75t_L g7827 ( 
.A(n_7188),
.Y(n_7827)
);

NOR2xp33_ASAP7_75t_L g7828 ( 
.A(n_7374),
.B(n_4879),
.Y(n_7828)
);

BUFx6f_ASAP7_75t_SL g7829 ( 
.A(n_7197),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7206),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_7209),
.Y(n_7831)
);

INVx2_ASAP7_75t_L g7832 ( 
.A(n_7190),
.Y(n_7832)
);

OR2x2_ASAP7_75t_L g7833 ( 
.A(n_7414),
.B(n_6983),
.Y(n_7833)
);

AND2x4_ASAP7_75t_L g7834 ( 
.A(n_7372),
.B(n_6853),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_7226),
.Y(n_7835)
);

INVx1_ASAP7_75t_L g7836 ( 
.A(n_7483),
.Y(n_7836)
);

AND2x2_ASAP7_75t_L g7837 ( 
.A(n_7448),
.B(n_6330),
.Y(n_7837)
);

INVx1_ASAP7_75t_L g7838 ( 
.A(n_7117),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7117),
.Y(n_7839)
);

OA21x2_ASAP7_75t_L g7840 ( 
.A1(n_7091),
.A2(n_7045),
.B(n_6977),
.Y(n_7840)
);

INVx1_ASAP7_75t_SL g7841 ( 
.A(n_7203),
.Y(n_7841)
);

NAND2xp5_ASAP7_75t_L g7842 ( 
.A(n_7368),
.B(n_6866),
.Y(n_7842)
);

INVx1_ASAP7_75t_L g7843 ( 
.A(n_7141),
.Y(n_7843)
);

INVx2_ASAP7_75t_L g7844 ( 
.A(n_7190),
.Y(n_7844)
);

OAI21xp5_ASAP7_75t_SL g7845 ( 
.A1(n_7108),
.A2(n_6496),
.B(n_5363),
.Y(n_7845)
);

AOI21xp5_ASAP7_75t_L g7846 ( 
.A1(n_7141),
.A2(n_6865),
.B(n_6857),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_7233),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_7235),
.Y(n_7848)
);

INVx4_ASAP7_75t_L g7849 ( 
.A(n_7386),
.Y(n_7849)
);

INVx2_ASAP7_75t_L g7850 ( 
.A(n_7205),
.Y(n_7850)
);

INVx1_ASAP7_75t_L g7851 ( 
.A(n_7244),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7252),
.Y(n_7852)
);

AND2x4_ASAP7_75t_L g7853 ( 
.A(n_7437),
.B(n_6857),
.Y(n_7853)
);

AND2x4_ASAP7_75t_L g7854 ( 
.A(n_7456),
.B(n_6865),
.Y(n_7854)
);

NAND2xp5_ASAP7_75t_L g7855 ( 
.A(n_7386),
.B(n_7387),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7256),
.Y(n_7856)
);

INVxp67_ASAP7_75t_SL g7857 ( 
.A(n_7205),
.Y(n_7857)
);

AOI221xp5_ASAP7_75t_L g7858 ( 
.A1(n_7173),
.A2(n_6923),
.B1(n_6933),
.B2(n_6919),
.C(n_6915),
.Y(n_7858)
);

BUFx2_ASAP7_75t_L g7859 ( 
.A(n_7325),
.Y(n_7859)
);

NAND2xp5_ASAP7_75t_L g7860 ( 
.A(n_7387),
.B(n_6888),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7257),
.Y(n_7861)
);

OA21x2_ASAP7_75t_L g7862 ( 
.A1(n_7091),
.A2(n_6977),
.B(n_6963),
.Y(n_7862)
);

OAI211xp5_ASAP7_75t_L g7863 ( 
.A1(n_7173),
.A2(n_7042),
.B(n_7071),
.C(n_6956),
.Y(n_7863)
);

BUFx6f_ASAP7_75t_L g7864 ( 
.A(n_7388),
.Y(n_7864)
);

OR2x6_ASAP7_75t_L g7865 ( 
.A(n_7116),
.B(n_3742),
.Y(n_7865)
);

AND2x2_ASAP7_75t_L g7866 ( 
.A(n_7453),
.B(n_6371),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7186),
.Y(n_7867)
);

OA21x2_ASAP7_75t_L g7868 ( 
.A1(n_7095),
.A2(n_6980),
.B(n_6963),
.Y(n_7868)
);

INVx2_ASAP7_75t_SL g7869 ( 
.A(n_7347),
.Y(n_7869)
);

INVx1_ASAP7_75t_L g7870 ( 
.A(n_7186),
.Y(n_7870)
);

AND2x2_ASAP7_75t_L g7871 ( 
.A(n_7455),
.B(n_6371),
.Y(n_7871)
);

INVx1_ASAP7_75t_L g7872 ( 
.A(n_7195),
.Y(n_7872)
);

OAI21x1_ASAP7_75t_L g7873 ( 
.A1(n_7242),
.A2(n_7071),
.B(n_6869),
.Y(n_7873)
);

A2O1A1Ixp33_ASAP7_75t_L g7874 ( 
.A1(n_7094),
.A2(n_6466),
.B(n_5705),
.C(n_6006),
.Y(n_7874)
);

AO21x2_ASAP7_75t_L g7875 ( 
.A1(n_7388),
.A2(n_6989),
.B(n_6987),
.Y(n_7875)
);

INVx2_ASAP7_75t_L g7876 ( 
.A(n_7207),
.Y(n_7876)
);

INVx2_ASAP7_75t_L g7877 ( 
.A(n_7207),
.Y(n_7877)
);

AOI21xp5_ASAP7_75t_L g7878 ( 
.A1(n_7183),
.A2(n_6869),
.B(n_6866),
.Y(n_7878)
);

OAI21xp33_ASAP7_75t_SL g7879 ( 
.A1(n_7344),
.A2(n_6298),
.B(n_6876),
.Y(n_7879)
);

HB1xp67_ASAP7_75t_L g7880 ( 
.A(n_7392),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7195),
.Y(n_7881)
);

INVx1_ASAP7_75t_L g7882 ( 
.A(n_7201),
.Y(n_7882)
);

AO21x2_ASAP7_75t_L g7883 ( 
.A1(n_7392),
.A2(n_6989),
.B(n_6987),
.Y(n_7883)
);

NAND2xp5_ASAP7_75t_L g7884 ( 
.A(n_7401),
.B(n_6876),
.Y(n_7884)
);

NAND2xp5_ASAP7_75t_L g7885 ( 
.A(n_7401),
.B(n_6880),
.Y(n_7885)
);

INVx2_ASAP7_75t_L g7886 ( 
.A(n_7789),
.Y(n_7886)
);

AO21x2_ASAP7_75t_L g7887 ( 
.A1(n_7528),
.A2(n_7338),
.B(n_7076),
.Y(n_7887)
);

NAND4xp75_ASAP7_75t_L g7888 ( 
.A(n_7574),
.B(n_7238),
.C(n_7232),
.D(n_7338),
.Y(n_7888)
);

NAND2xp5_ASAP7_75t_L g7889 ( 
.A(n_7513),
.B(n_7208),
.Y(n_7889)
);

NOR3xp33_ASAP7_75t_L g7890 ( 
.A(n_7560),
.B(n_7176),
.C(n_7174),
.Y(n_7890)
);

HB1xp67_ASAP7_75t_L g7891 ( 
.A(n_7576),
.Y(n_7891)
);

INVx1_ASAP7_75t_L g7892 ( 
.A(n_7602),
.Y(n_7892)
);

BUFx3_ASAP7_75t_L g7893 ( 
.A(n_7647),
.Y(n_7893)
);

NAND4xp75_ASAP7_75t_L g7894 ( 
.A(n_7571),
.B(n_7179),
.C(n_7158),
.D(n_7160),
.Y(n_7894)
);

OAI21xp5_ASAP7_75t_L g7895 ( 
.A1(n_7541),
.A2(n_7261),
.B(n_7202),
.Y(n_7895)
);

NOR2xp33_ASAP7_75t_L g7896 ( 
.A(n_7589),
.B(n_7151),
.Y(n_7896)
);

OR2x2_ASAP7_75t_L g7897 ( 
.A(n_7514),
.B(n_7231),
.Y(n_7897)
);

AOI221xp5_ASAP7_75t_L g7898 ( 
.A1(n_7517),
.A2(n_7183),
.B1(n_7328),
.B2(n_7201),
.C(n_7264),
.Y(n_7898)
);

NOR3xp33_ASAP7_75t_L g7899 ( 
.A(n_7660),
.B(n_7165),
.C(n_7161),
.Y(n_7899)
);

INVx2_ASAP7_75t_SL g7900 ( 
.A(n_7789),
.Y(n_7900)
);

NOR3xp33_ASAP7_75t_L g7901 ( 
.A(n_7777),
.B(n_7170),
.C(n_7189),
.Y(n_7901)
);

BUFx3_ASAP7_75t_L g7902 ( 
.A(n_7648),
.Y(n_7902)
);

AND2x2_ASAP7_75t_L g7903 ( 
.A(n_7548),
.B(n_7215),
.Y(n_7903)
);

HB1xp67_ASAP7_75t_L g7904 ( 
.A(n_7641),
.Y(n_7904)
);

OR2x2_ASAP7_75t_L g7905 ( 
.A(n_7714),
.B(n_7729),
.Y(n_7905)
);

AOI22xp33_ASAP7_75t_L g7906 ( 
.A1(n_7534),
.A2(n_7270),
.B1(n_7262),
.B2(n_7348),
.Y(n_7906)
);

AND2x2_ASAP7_75t_L g7907 ( 
.A(n_7573),
.B(n_7216),
.Y(n_7907)
);

INVxp67_ASAP7_75t_SL g7908 ( 
.A(n_7666),
.Y(n_7908)
);

INVx3_ASAP7_75t_L g7909 ( 
.A(n_7639),
.Y(n_7909)
);

AOI22xp33_ASAP7_75t_L g7910 ( 
.A1(n_7516),
.A2(n_7415),
.B1(n_7414),
.B2(n_7486),
.Y(n_7910)
);

AND2x2_ASAP7_75t_L g7911 ( 
.A(n_7575),
.B(n_7709),
.Y(n_7911)
);

AND2x4_ASAP7_75t_L g7912 ( 
.A(n_7785),
.B(n_7503),
.Y(n_7912)
);

NAND2xp5_ASAP7_75t_L g7913 ( 
.A(n_7644),
.B(n_7738),
.Y(n_7913)
);

NAND3xp33_ASAP7_75t_L g7914 ( 
.A(n_7580),
.B(n_7441),
.C(n_7250),
.Y(n_7914)
);

NAND3xp33_ASAP7_75t_L g7915 ( 
.A(n_7532),
.B(n_7321),
.C(n_7249),
.Y(n_7915)
);

AO21x2_ASAP7_75t_L g7916 ( 
.A1(n_7637),
.A2(n_7076),
.B(n_7282),
.Y(n_7916)
);

INVx1_ASAP7_75t_L g7917 ( 
.A(n_7668),
.Y(n_7917)
);

NAND2xp5_ASAP7_75t_L g7918 ( 
.A(n_7749),
.B(n_7208),
.Y(n_7918)
);

NAND2xp5_ASAP7_75t_L g7919 ( 
.A(n_7520),
.B(n_7217),
.Y(n_7919)
);

INVxp67_ASAP7_75t_SL g7920 ( 
.A(n_7765),
.Y(n_7920)
);

AND2x2_ASAP7_75t_L g7921 ( 
.A(n_7610),
.B(n_7224),
.Y(n_7921)
);

NOR3xp33_ASAP7_75t_L g7922 ( 
.A(n_7600),
.B(n_7498),
.C(n_7328),
.Y(n_7922)
);

NAND3xp33_ASAP7_75t_L g7923 ( 
.A(n_7565),
.B(n_7358),
.C(n_7323),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7512),
.Y(n_7924)
);

AOI221xp5_ASAP7_75t_L g7925 ( 
.A1(n_7829),
.A2(n_7268),
.B1(n_7275),
.B2(n_7266),
.C(n_7259),
.Y(n_7925)
);

NAND4xp75_ASAP7_75t_L g7926 ( 
.A(n_7546),
.B(n_7283),
.C(n_7286),
.D(n_7282),
.Y(n_7926)
);

NAND2xp5_ASAP7_75t_L g7927 ( 
.A(n_7859),
.B(n_7217),
.Y(n_7927)
);

AND2x2_ASAP7_75t_L g7928 ( 
.A(n_7564),
.B(n_7679),
.Y(n_7928)
);

OR2x2_ASAP7_75t_L g7929 ( 
.A(n_7572),
.B(n_7558),
.Y(n_7929)
);

NAND4xp75_ASAP7_75t_L g7930 ( 
.A(n_7533),
.B(n_7286),
.C(n_7326),
.D(n_7283),
.Y(n_7930)
);

AOI22xp5_ASAP7_75t_L g7931 ( 
.A1(n_7829),
.A2(n_7503),
.B1(n_7498),
.B2(n_7480),
.Y(n_7931)
);

OR2x2_ASAP7_75t_L g7932 ( 
.A(n_7695),
.B(n_7412),
.Y(n_7932)
);

AND2x2_ASAP7_75t_L g7933 ( 
.A(n_7570),
.B(n_7371),
.Y(n_7933)
);

NAND4xp75_ASAP7_75t_L g7934 ( 
.A(n_7633),
.B(n_7337),
.C(n_7326),
.D(n_7432),
.Y(n_7934)
);

AND2x2_ASAP7_75t_L g7935 ( 
.A(n_7557),
.B(n_7375),
.Y(n_7935)
);

XNOR2xp5_ASAP7_75t_L g7936 ( 
.A(n_7649),
.B(n_7480),
.Y(n_7936)
);

NAND3xp33_ASAP7_75t_L g7937 ( 
.A(n_7806),
.B(n_7440),
.C(n_7432),
.Y(n_7937)
);

OR2x2_ASAP7_75t_L g7938 ( 
.A(n_7568),
.B(n_7412),
.Y(n_7938)
);

AND2x2_ASAP7_75t_L g7939 ( 
.A(n_7523),
.B(n_7502),
.Y(n_7939)
);

AOI22xp33_ASAP7_75t_L g7940 ( 
.A1(n_7767),
.A2(n_7415),
.B1(n_7333),
.B2(n_7340),
.Y(n_7940)
);

NAND4xp75_ASAP7_75t_L g7941 ( 
.A(n_7686),
.B(n_7337),
.C(n_7465),
.D(n_7440),
.Y(n_7941)
);

OA21x2_ASAP7_75t_L g7942 ( 
.A1(n_7527),
.A2(n_7004),
.B(n_6999),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7512),
.Y(n_7943)
);

AOI22xp33_ASAP7_75t_L g7944 ( 
.A1(n_7683),
.A2(n_7460),
.B1(n_7279),
.B2(n_7280),
.Y(n_7944)
);

AND2x2_ASAP7_75t_L g7945 ( 
.A(n_7526),
.B(n_7409),
.Y(n_7945)
);

INVx3_ASAP7_75t_L g7946 ( 
.A(n_7639),
.Y(n_7946)
);

NOR3xp33_ASAP7_75t_L g7947 ( 
.A(n_7657),
.B(n_7287),
.C(n_7274),
.Y(n_7947)
);

AOI22xp33_ASAP7_75t_L g7948 ( 
.A1(n_7694),
.A2(n_7284),
.B1(n_7290),
.B2(n_7276),
.Y(n_7948)
);

INVx2_ASAP7_75t_L g7949 ( 
.A(n_7789),
.Y(n_7949)
);

OR2x2_ASAP7_75t_L g7950 ( 
.A(n_7566),
.B(n_7277),
.Y(n_7950)
);

NAND2xp5_ASAP7_75t_L g7951 ( 
.A(n_7608),
.B(n_7228),
.Y(n_7951)
);

AND2x2_ASAP7_75t_L g7952 ( 
.A(n_7601),
.B(n_7350),
.Y(n_7952)
);

AOI22xp33_ASAP7_75t_L g7953 ( 
.A1(n_7530),
.A2(n_7297),
.B1(n_7301),
.B2(n_7304),
.Y(n_7953)
);

NAND3xp33_ASAP7_75t_L g7954 ( 
.A(n_7583),
.B(n_7493),
.C(n_7465),
.Y(n_7954)
);

NOR2xp33_ASAP7_75t_L g7955 ( 
.A(n_7673),
.B(n_7698),
.Y(n_7955)
);

NOR3xp33_ASAP7_75t_L g7956 ( 
.A(n_7588),
.B(n_7287),
.C(n_7274),
.Y(n_7956)
);

NOR2xp33_ASAP7_75t_L g7957 ( 
.A(n_7585),
.B(n_7491),
.Y(n_7957)
);

AND2x4_ASAP7_75t_SL g7958 ( 
.A(n_7515),
.B(n_4879),
.Y(n_7958)
);

NAND2xp5_ASAP7_75t_L g7959 ( 
.A(n_7796),
.B(n_7228),
.Y(n_7959)
);

AND2x2_ASAP7_75t_L g7960 ( 
.A(n_7638),
.B(n_7491),
.Y(n_7960)
);

NAND4xp75_ASAP7_75t_L g7961 ( 
.A(n_7595),
.B(n_7696),
.C(n_7587),
.D(n_7662),
.Y(n_7961)
);

NOR3xp33_ASAP7_75t_L g7962 ( 
.A(n_7519),
.B(n_7322),
.C(n_7281),
.Y(n_7962)
);

AND2x2_ASAP7_75t_L g7963 ( 
.A(n_7559),
.B(n_7345),
.Y(n_7963)
);

NAND2xp5_ASAP7_75t_L g7964 ( 
.A(n_7803),
.B(n_7272),
.Y(n_7964)
);

INVx2_ASAP7_75t_L g7965 ( 
.A(n_7785),
.Y(n_7965)
);

NAND3xp33_ASAP7_75t_L g7966 ( 
.A(n_7590),
.B(n_7493),
.C(n_7281),
.Y(n_7966)
);

AND2x2_ASAP7_75t_L g7967 ( 
.A(n_7582),
.B(n_7613),
.Y(n_7967)
);

INVx1_ASAP7_75t_L g7968 ( 
.A(n_7518),
.Y(n_7968)
);

INVx1_ASAP7_75t_SL g7969 ( 
.A(n_7744),
.Y(n_7969)
);

NAND4xp75_ASAP7_75t_L g7970 ( 
.A(n_7692),
.B(n_7272),
.C(n_7509),
.D(n_7500),
.Y(n_7970)
);

AND2x2_ASAP7_75t_L g7971 ( 
.A(n_7640),
.B(n_7377),
.Y(n_7971)
);

AO21x2_ASAP7_75t_L g7972 ( 
.A1(n_7529),
.A2(n_7097),
.B(n_7095),
.Y(n_7972)
);

NOR2x1_ASAP7_75t_L g7973 ( 
.A(n_7535),
.B(n_7097),
.Y(n_7973)
);

NAND3xp33_ASAP7_75t_L g7974 ( 
.A(n_7551),
.B(n_7285),
.C(n_7278),
.Y(n_7974)
);

NAND3xp33_ASAP7_75t_L g7975 ( 
.A(n_7552),
.B(n_7294),
.C(n_7292),
.Y(n_7975)
);

CKINVDCx20_ASAP7_75t_R g7976 ( 
.A(n_7592),
.Y(n_7976)
);

OR2x2_ASAP7_75t_L g7977 ( 
.A(n_7555),
.B(n_7298),
.Y(n_7977)
);

NAND2xp5_ASAP7_75t_L g7978 ( 
.A(n_7653),
.B(n_7500),
.Y(n_7978)
);

AND2x2_ASAP7_75t_L g7979 ( 
.A(n_7642),
.B(n_7380),
.Y(n_7979)
);

OR2x2_ASAP7_75t_L g7980 ( 
.A(n_7577),
.B(n_7289),
.Y(n_7980)
);

AOI22xp33_ASAP7_75t_L g7981 ( 
.A1(n_7515),
.A2(n_7354),
.B1(n_7366),
.B2(n_7353),
.Y(n_7981)
);

AOI22xp33_ASAP7_75t_SL g7982 ( 
.A1(n_7627),
.A2(n_7444),
.B1(n_7462),
.B2(n_7435),
.Y(n_7982)
);

OA211x2_ASAP7_75t_L g7983 ( 
.A1(n_7616),
.A2(n_7221),
.B(n_7255),
.C(n_7219),
.Y(n_7983)
);

OAI211xp5_ASAP7_75t_SL g7984 ( 
.A1(n_7584),
.A2(n_7307),
.B(n_7312),
.C(n_7299),
.Y(n_7984)
);

OR2x2_ASAP7_75t_L g7985 ( 
.A(n_7739),
.B(n_7322),
.Y(n_7985)
);

NOR2x1_ASAP7_75t_SL g7986 ( 
.A(n_7634),
.B(n_7509),
.Y(n_7986)
);

OR2x2_ASAP7_75t_L g7987 ( 
.A(n_7556),
.B(n_7219),
.Y(n_7987)
);

NAND4xp75_ASAP7_75t_L g7988 ( 
.A(n_7543),
.B(n_7447),
.C(n_7507),
.D(n_7450),
.Y(n_7988)
);

NAND3xp33_ASAP7_75t_L g7989 ( 
.A(n_7596),
.B(n_7494),
.C(n_7492),
.Y(n_7989)
);

AND2x2_ASAP7_75t_L g7990 ( 
.A(n_7540),
.B(n_7393),
.Y(n_7990)
);

NAND4xp75_ASAP7_75t_L g7991 ( 
.A(n_7550),
.B(n_7814),
.C(n_7774),
.D(n_7620),
.Y(n_7991)
);

AND2x2_ASAP7_75t_L g7992 ( 
.A(n_7553),
.B(n_7396),
.Y(n_7992)
);

AND2x2_ASAP7_75t_L g7993 ( 
.A(n_7652),
.B(n_7397),
.Y(n_7993)
);

AND2x2_ASAP7_75t_L g7994 ( 
.A(n_7562),
.B(n_7400),
.Y(n_7994)
);

AND2x2_ASAP7_75t_L g7995 ( 
.A(n_7740),
.B(n_7419),
.Y(n_7995)
);

OR2x2_ASAP7_75t_L g7996 ( 
.A(n_7833),
.B(n_7221),
.Y(n_7996)
);

NAND3xp33_ASAP7_75t_L g7997 ( 
.A(n_7598),
.B(n_7464),
.C(n_7463),
.Y(n_7997)
);

AOI22xp5_ASAP7_75t_L g7998 ( 
.A1(n_7795),
.A2(n_7313),
.B1(n_7331),
.B2(n_7317),
.Y(n_7998)
);

NAND3xp33_ASAP7_75t_L g7999 ( 
.A(n_7678),
.B(n_7479),
.C(n_7469),
.Y(n_7999)
);

AND2x2_ASAP7_75t_L g8000 ( 
.A(n_7755),
.B(n_7425),
.Y(n_8000)
);

INVx2_ASAP7_75t_L g8001 ( 
.A(n_7812),
.Y(n_8001)
);

AND2x2_ASAP7_75t_L g8002 ( 
.A(n_7869),
.B(n_7426),
.Y(n_8002)
);

BUFx2_ASAP7_75t_L g8003 ( 
.A(n_7656),
.Y(n_8003)
);

NAND2xp5_ASAP7_75t_L g8004 ( 
.A(n_7841),
.B(n_7434),
.Y(n_8004)
);

NAND2xp5_ASAP7_75t_L g8005 ( 
.A(n_7816),
.B(n_7442),
.Y(n_8005)
);

OR2x2_ASAP7_75t_L g8006 ( 
.A(n_7522),
.B(n_7255),
.Y(n_8006)
);

AND2x2_ASAP7_75t_L g8007 ( 
.A(n_7801),
.B(n_7430),
.Y(n_8007)
);

AND2x2_ASAP7_75t_L g8008 ( 
.A(n_7728),
.B(n_7430),
.Y(n_8008)
);

NOR2xp33_ASAP7_75t_L g8009 ( 
.A(n_7547),
.B(n_7501),
.Y(n_8009)
);

NAND3xp33_ASAP7_75t_L g8010 ( 
.A(n_7800),
.B(n_7510),
.C(n_7336),
.Y(n_8010)
);

NAND3xp33_ASAP7_75t_L g8011 ( 
.A(n_7780),
.B(n_7452),
.C(n_7451),
.Y(n_8011)
);

XNOR2xp5_ASAP7_75t_L g8012 ( 
.A(n_7599),
.B(n_5193),
.Y(n_8012)
);

AOI22xp5_ASAP7_75t_L g8013 ( 
.A1(n_7619),
.A2(n_7334),
.B1(n_7351),
.B2(n_7342),
.Y(n_8013)
);

OR2x2_ASAP7_75t_L g8014 ( 
.A(n_7622),
.B(n_7314),
.Y(n_8014)
);

NAND4xp75_ASAP7_75t_L g8015 ( 
.A(n_7623),
.B(n_7357),
.C(n_7360),
.D(n_7352),
.Y(n_8015)
);

OR2x2_ASAP7_75t_L g8016 ( 
.A(n_7531),
.B(n_7315),
.Y(n_8016)
);

NAND2xp5_ASAP7_75t_L g8017 ( 
.A(n_7816),
.B(n_7362),
.Y(n_8017)
);

AOI22xp5_ASAP7_75t_L g8018 ( 
.A1(n_7629),
.A2(n_7376),
.B1(n_7379),
.B2(n_7373),
.Y(n_8018)
);

NAND2x1p5_ASAP7_75t_L g8019 ( 
.A(n_7656),
.B(n_7435),
.Y(n_8019)
);

INVx2_ASAP7_75t_L g8020 ( 
.A(n_7812),
.Y(n_8020)
);

AND2x2_ASAP7_75t_L g8021 ( 
.A(n_7625),
.B(n_7444),
.Y(n_8021)
);

NAND3xp33_ASAP7_75t_L g8022 ( 
.A(n_7703),
.B(n_7458),
.C(n_7454),
.Y(n_8022)
);

NAND2xp5_ASAP7_75t_L g8023 ( 
.A(n_7761),
.B(n_7381),
.Y(n_8023)
);

NAND4xp25_ASAP7_75t_L g8024 ( 
.A(n_7621),
.B(n_7495),
.C(n_7497),
.D(n_7467),
.Y(n_8024)
);

NAND4xp75_ASAP7_75t_L g8025 ( 
.A(n_7646),
.B(n_7398),
.C(n_7405),
.D(n_7391),
.Y(n_8025)
);

OR2x2_ASAP7_75t_L g8026 ( 
.A(n_7757),
.B(n_7329),
.Y(n_8026)
);

AND2x2_ASAP7_75t_L g8027 ( 
.A(n_7525),
.B(n_7462),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7525),
.B(n_7347),
.Y(n_8028)
);

NAND3xp33_ASAP7_75t_L g8029 ( 
.A(n_7667),
.B(n_7418),
.C(n_7417),
.Y(n_8029)
);

NAND3xp33_ASAP7_75t_L g8030 ( 
.A(n_7779),
.B(n_7427),
.C(n_7423),
.Y(n_8030)
);

NOR3xp33_ASAP7_75t_L g8031 ( 
.A(n_7826),
.B(n_7428),
.C(n_7369),
.Y(n_8031)
);

BUFx2_ASAP7_75t_L g8032 ( 
.A(n_7578),
.Y(n_8032)
);

XNOR2xp5_ASAP7_75t_L g8033 ( 
.A(n_7687),
.B(n_5294),
.Y(n_8033)
);

NAND2xp5_ASAP7_75t_L g8034 ( 
.A(n_7766),
.B(n_7477),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_7518),
.Y(n_8035)
);

INVx2_ASAP7_75t_SL g8036 ( 
.A(n_7669),
.Y(n_8036)
);

NAND3xp33_ASAP7_75t_L g8037 ( 
.A(n_7535),
.B(n_7477),
.C(n_7369),
.Y(n_8037)
);

OAI211xp5_ASAP7_75t_L g8038 ( 
.A1(n_7631),
.A2(n_7389),
.B(n_7406),
.C(n_7365),
.Y(n_8038)
);

NOR3xp33_ASAP7_75t_L g8039 ( 
.A(n_7628),
.B(n_7389),
.C(n_7365),
.Y(n_8039)
);

HB1xp67_ASAP7_75t_L g8040 ( 
.A(n_7864),
.Y(n_8040)
);

NAND3xp33_ASAP7_75t_L g8041 ( 
.A(n_7628),
.B(n_7416),
.C(n_7406),
.Y(n_8041)
);

NAND2xp5_ASAP7_75t_L g8042 ( 
.A(n_7721),
.B(n_7416),
.Y(n_8042)
);

OAI211xp5_ASAP7_75t_L g8043 ( 
.A1(n_7685),
.A2(n_7429),
.B(n_7433),
.C(n_7422),
.Y(n_8043)
);

XOR2x2_ASAP7_75t_L g8044 ( 
.A(n_7828),
.B(n_4985),
.Y(n_8044)
);

AND2x2_ASAP7_75t_L g8045 ( 
.A(n_7634),
.B(n_6361),
.Y(n_8045)
);

NAND3xp33_ASAP7_75t_L g8046 ( 
.A(n_7858),
.B(n_7429),
.C(n_7422),
.Y(n_8046)
);

AND2x2_ASAP7_75t_L g8047 ( 
.A(n_7865),
.B(n_6361),
.Y(n_8047)
);

OAI211xp5_ASAP7_75t_SL g8048 ( 
.A1(n_7594),
.A2(n_7484),
.B(n_7487),
.C(n_7468),
.Y(n_8048)
);

OAI211xp5_ASAP7_75t_SL g8049 ( 
.A1(n_7597),
.A2(n_7484),
.B(n_7487),
.C(n_7468),
.Y(n_8049)
);

NOR3xp33_ASAP7_75t_L g8050 ( 
.A(n_7605),
.B(n_7561),
.C(n_7536),
.Y(n_8050)
);

AND2x2_ASAP7_75t_L g8051 ( 
.A(n_7865),
.B(n_6373),
.Y(n_8051)
);

NOR2xp33_ASAP7_75t_L g8052 ( 
.A(n_7563),
.B(n_7370),
.Y(n_8052)
);

INVx2_ASAP7_75t_L g8053 ( 
.A(n_7864),
.Y(n_8053)
);

NOR2x1_ASAP7_75t_L g8054 ( 
.A(n_7521),
.B(n_7099),
.Y(n_8054)
);

NOR2xp33_ASAP7_75t_R g8055 ( 
.A(n_7586),
.B(n_5125),
.Y(n_8055)
);

AND2x4_ASAP7_75t_SL g8056 ( 
.A(n_7671),
.B(n_5350),
.Y(n_8056)
);

NAND3xp33_ASAP7_75t_L g8057 ( 
.A(n_7579),
.B(n_7449),
.C(n_7433),
.Y(n_8057)
);

AOI22xp33_ASAP7_75t_L g8058 ( 
.A1(n_7650),
.A2(n_5574),
.B1(n_6046),
.B2(n_7408),
.Y(n_8058)
);

NOR3xp33_ASAP7_75t_L g8059 ( 
.A(n_7797),
.B(n_7461),
.C(n_7449),
.Y(n_8059)
);

INVx1_ASAP7_75t_SL g8060 ( 
.A(n_7834),
.Y(n_8060)
);

OR2x2_ASAP7_75t_L g8061 ( 
.A(n_7636),
.B(n_7420),
.Y(n_8061)
);

NOR2xp33_ASAP7_75t_L g8062 ( 
.A(n_7611),
.B(n_7436),
.Y(n_8062)
);

AOI22xp5_ASAP7_75t_L g8063 ( 
.A1(n_7654),
.A2(n_6046),
.B1(n_5574),
.B2(n_5964),
.Y(n_8063)
);

AOI22xp33_ASAP7_75t_SL g8064 ( 
.A1(n_7549),
.A2(n_6046),
.B1(n_5188),
.B2(n_4942),
.Y(n_8064)
);

OR2x2_ASAP7_75t_L g8065 ( 
.A(n_7764),
.B(n_7023),
.Y(n_8065)
);

AOI22xp33_ASAP7_75t_L g8066 ( 
.A1(n_7770),
.A2(n_6046),
.B1(n_6919),
.B2(n_6915),
.Y(n_8066)
);

NAND3xp33_ASAP7_75t_L g8067 ( 
.A(n_7677),
.B(n_7466),
.C(n_7461),
.Y(n_8067)
);

INVx1_ASAP7_75t_L g8068 ( 
.A(n_7521),
.Y(n_8068)
);

XOR2x2_ASAP7_75t_L g8069 ( 
.A(n_7630),
.B(n_4985),
.Y(n_8069)
);

AOI22xp33_ASAP7_75t_L g8070 ( 
.A1(n_7727),
.A2(n_6933),
.B1(n_6937),
.B2(n_6923),
.Y(n_8070)
);

AOI22xp33_ASAP7_75t_L g8071 ( 
.A1(n_7772),
.A2(n_6955),
.B1(n_6956),
.B2(n_6937),
.Y(n_8071)
);

AND2x2_ASAP7_75t_L g8072 ( 
.A(n_7743),
.B(n_6373),
.Y(n_8072)
);

HB1xp67_ASAP7_75t_L g8073 ( 
.A(n_7864),
.Y(n_8073)
);

AND2x2_ASAP7_75t_L g8074 ( 
.A(n_7837),
.B(n_6390),
.Y(n_8074)
);

AOI22xp33_ASAP7_75t_L g8075 ( 
.A1(n_7866),
.A2(n_6955),
.B1(n_6888),
.B2(n_6889),
.Y(n_8075)
);

NOR2x1_ASAP7_75t_L g8076 ( 
.A(n_7524),
.B(n_7099),
.Y(n_8076)
);

OA211x2_ASAP7_75t_L g8077 ( 
.A1(n_7775),
.A2(n_7466),
.B(n_6192),
.C(n_4665),
.Y(n_8077)
);

OR2x2_ASAP7_75t_L g8078 ( 
.A(n_7754),
.B(n_7060),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7524),
.Y(n_8079)
);

OR2x2_ASAP7_75t_L g8080 ( 
.A(n_7768),
.B(n_7771),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_7537),
.Y(n_8081)
);

NAND4xp75_ASAP7_75t_L g8082 ( 
.A(n_7658),
.B(n_7112),
.C(n_7114),
.D(n_7102),
.Y(n_8082)
);

BUFx2_ASAP7_75t_L g8083 ( 
.A(n_7822),
.Y(n_8083)
);

HB1xp67_ASAP7_75t_L g8084 ( 
.A(n_7790),
.Y(n_8084)
);

AND2x4_ASAP7_75t_L g8085 ( 
.A(n_7822),
.B(n_6880),
.Y(n_8085)
);

AND2x2_ASAP7_75t_L g8086 ( 
.A(n_7871),
.B(n_6137),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_7537),
.Y(n_8087)
);

NAND2xp5_ASAP7_75t_L g8088 ( 
.A(n_7626),
.B(n_6889),
.Y(n_8088)
);

NAND2xp5_ASAP7_75t_L g8089 ( 
.A(n_7635),
.B(n_6137),
.Y(n_8089)
);

OA211x2_ASAP7_75t_L g8090 ( 
.A1(n_7855),
.A2(n_6192),
.B(n_5171),
.C(n_5170),
.Y(n_8090)
);

AOI22xp5_ASAP7_75t_L g8091 ( 
.A1(n_7661),
.A2(n_5964),
.B1(n_4942),
.B2(n_4918),
.Y(n_8091)
);

AO21x2_ASAP7_75t_L g8092 ( 
.A1(n_7836),
.A2(n_7112),
.B(n_7102),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_7538),
.Y(n_8093)
);

NAND4xp75_ASAP7_75t_L g8094 ( 
.A(n_7665),
.B(n_7121),
.C(n_7126),
.D(n_7114),
.Y(n_8094)
);

AND2x2_ASAP7_75t_L g8095 ( 
.A(n_7702),
.B(n_6138),
.Y(n_8095)
);

NAND2xp5_ASAP7_75t_L g8096 ( 
.A(n_7643),
.B(n_6569),
.Y(n_8096)
);

AND2x4_ASAP7_75t_L g8097 ( 
.A(n_7849),
.B(n_6298),
.Y(n_8097)
);

NAND3xp33_ASAP7_75t_L g8098 ( 
.A(n_7677),
.B(n_7126),
.C(n_7121),
.Y(n_8098)
);

AOI221xp5_ASAP7_75t_L g8099 ( 
.A1(n_7708),
.A2(n_7674),
.B1(n_7737),
.B2(n_7730),
.C(n_7663),
.Y(n_8099)
);

AOI22xp33_ASAP7_75t_L g8100 ( 
.A1(n_7611),
.A2(n_5964),
.B1(n_5052),
.B2(n_4905),
.Y(n_8100)
);

NAND2xp5_ASAP7_75t_L g8101 ( 
.A(n_7659),
.B(n_6576),
.Y(n_8101)
);

AND2x2_ASAP7_75t_L g8102 ( 
.A(n_7751),
.B(n_6138),
.Y(n_8102)
);

AND2x4_ASAP7_75t_L g8103 ( 
.A(n_7849),
.B(n_6144),
.Y(n_8103)
);

NOR2xp33_ASAP7_75t_L g8104 ( 
.A(n_7671),
.B(n_4985),
.Y(n_8104)
);

AND4x1_ASAP7_75t_L g8105 ( 
.A(n_7538),
.B(n_7544),
.C(n_7545),
.D(n_7567),
.Y(n_8105)
);

OR2x2_ASAP7_75t_L g8106 ( 
.A(n_7810),
.B(n_7062),
.Y(n_8106)
);

NOR3xp33_ASAP7_75t_L g8107 ( 
.A(n_7586),
.B(n_7632),
.C(n_7711),
.Y(n_8107)
);

NOR3xp33_ASAP7_75t_L g8108 ( 
.A(n_7632),
.B(n_6980),
.C(n_6999),
.Y(n_8108)
);

NAND4xp75_ASAP7_75t_L g8109 ( 
.A(n_7645),
.B(n_7581),
.C(n_7604),
.D(n_7591),
.Y(n_8109)
);

INVx3_ASAP7_75t_L g8110 ( 
.A(n_7677),
.Y(n_8110)
);

OR2x2_ASAP7_75t_L g8111 ( 
.A(n_7655),
.B(n_6192),
.Y(n_8111)
);

OR2x2_ASAP7_75t_L g8112 ( 
.A(n_7688),
.B(n_6192),
.Y(n_8112)
);

NOR2xp33_ASAP7_75t_L g8113 ( 
.A(n_7713),
.B(n_5360),
.Y(n_8113)
);

NAND3xp33_ASAP7_75t_SL g8114 ( 
.A(n_7682),
.B(n_5923),
.C(n_7004),
.Y(n_8114)
);

INVx1_ASAP7_75t_L g8115 ( 
.A(n_7544),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7690),
.Y(n_8116)
);

OR2x2_ASAP7_75t_L g8117 ( 
.A(n_7717),
.B(n_6356),
.Y(n_8117)
);

AND2x2_ASAP7_75t_L g8118 ( 
.A(n_7751),
.B(n_6144),
.Y(n_8118)
);

NAND3xp33_ASAP7_75t_SL g8119 ( 
.A(n_7769),
.B(n_7020),
.C(n_7005),
.Y(n_8119)
);

NOR2x1_ASAP7_75t_L g8120 ( 
.A(n_7545),
.B(n_7005),
.Y(n_8120)
);

NAND4xp75_ASAP7_75t_L g8121 ( 
.A(n_7615),
.B(n_7026),
.C(n_7027),
.D(n_7020),
.Y(n_8121)
);

OR2x2_ASAP7_75t_L g8122 ( 
.A(n_7720),
.B(n_6356),
.Y(n_8122)
);

AND2x2_ASAP7_75t_L g8123 ( 
.A(n_7664),
.B(n_6163),
.Y(n_8123)
);

OR2x2_ASAP7_75t_L g8124 ( 
.A(n_7786),
.B(n_6270),
.Y(n_8124)
);

OR2x2_ASAP7_75t_L g8125 ( 
.A(n_7787),
.B(n_6270),
.Y(n_8125)
);

OR2x2_ASAP7_75t_L g8126 ( 
.A(n_7793),
.B(n_6579),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_7715),
.B(n_6581),
.Y(n_8127)
);

NAND3xp33_ASAP7_75t_L g8128 ( 
.A(n_7863),
.B(n_7027),
.C(n_7026),
.Y(n_8128)
);

NAND3xp33_ASAP7_75t_L g8129 ( 
.A(n_7758),
.B(n_7029),
.C(n_4911),
.Y(n_8129)
);

OR2x2_ASAP7_75t_L g8130 ( 
.A(n_7799),
.B(n_6584),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_7836),
.Y(n_8131)
);

INVx2_ASAP7_75t_L g8132 ( 
.A(n_7690),
.Y(n_8132)
);

AND2x2_ASAP7_75t_L g8133 ( 
.A(n_7834),
.B(n_7853),
.Y(n_8133)
);

AOI22xp33_ASAP7_75t_SL g8134 ( 
.A1(n_7539),
.A2(n_4918),
.B1(n_4942),
.B2(n_5195),
.Y(n_8134)
);

AND2x2_ASAP7_75t_L g8135 ( 
.A(n_7853),
.B(n_7854),
.Y(n_8135)
);

AND2x2_ASAP7_75t_L g8136 ( 
.A(n_7854),
.B(n_6163),
.Y(n_8136)
);

NOR2xp33_ASAP7_75t_L g8137 ( 
.A(n_7670),
.B(n_6176),
.Y(n_8137)
);

AND2x2_ASAP7_75t_L g8138 ( 
.A(n_7672),
.B(n_6176),
.Y(n_8138)
);

NAND3xp33_ASAP7_75t_L g8139 ( 
.A(n_7807),
.B(n_7029),
.C(n_4911),
.Y(n_8139)
);

INVx1_ASAP7_75t_L g8140 ( 
.A(n_7792),
.Y(n_8140)
);

AND2x2_ASAP7_75t_L g8141 ( 
.A(n_7676),
.B(n_5790),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_7792),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7794),
.Y(n_8143)
);

INVx2_ASAP7_75t_L g8144 ( 
.A(n_7690),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7794),
.Y(n_8145)
);

AND2x2_ASAP7_75t_L g8146 ( 
.A(n_7857),
.B(n_5790),
.Y(n_8146)
);

NAND3xp33_ASAP7_75t_L g8147 ( 
.A(n_7809),
.B(n_7846),
.C(n_7815),
.Y(n_8147)
);

INVx1_ASAP7_75t_L g8148 ( 
.A(n_7808),
.Y(n_8148)
);

AND2x2_ASAP7_75t_L g8149 ( 
.A(n_7773),
.B(n_5790),
.Y(n_8149)
);

NAND4xp75_ASAP7_75t_L g8150 ( 
.A(n_7569),
.B(n_6081),
.C(n_6401),
.D(n_6359),
.Y(n_8150)
);

AND2x2_ASAP7_75t_L g8151 ( 
.A(n_7773),
.B(n_7603),
.Y(n_8151)
);

AND2x2_ASAP7_75t_L g8152 ( 
.A(n_7606),
.B(n_5833),
.Y(n_8152)
);

AND2x2_ASAP7_75t_L g8153 ( 
.A(n_7607),
.B(n_7760),
.Y(n_8153)
);

NAND2xp5_ASAP7_75t_L g8154 ( 
.A(n_7684),
.B(n_6048),
.Y(n_8154)
);

AOI221xp5_ASAP7_75t_L g8155 ( 
.A1(n_7838),
.A2(n_6571),
.B1(n_6562),
.B2(n_6618),
.C(n_6597),
.Y(n_8155)
);

AOI22xp33_ASAP7_75t_L g8156 ( 
.A1(n_7838),
.A2(n_5964),
.B1(n_5052),
.B2(n_4905),
.Y(n_8156)
);

NOR3xp33_ASAP7_75t_L g8157 ( 
.A(n_7745),
.B(n_5318),
.C(n_5297),
.Y(n_8157)
);

OAI211xp5_ASAP7_75t_SL g8158 ( 
.A1(n_7839),
.A2(n_6560),
.B(n_6552),
.C(n_5375),
.Y(n_8158)
);

OAI211xp5_ASAP7_75t_SL g8159 ( 
.A1(n_7839),
.A2(n_6560),
.B(n_6552),
.C(n_5418),
.Y(n_8159)
);

NAND3xp33_ASAP7_75t_L g8160 ( 
.A(n_7719),
.B(n_6081),
.C(n_6249),
.Y(n_8160)
);

AND2x2_ASAP7_75t_L g8161 ( 
.A(n_7680),
.B(n_5833),
.Y(n_8161)
);

NOR3xp33_ASAP7_75t_L g8162 ( 
.A(n_7746),
.B(n_5318),
.C(n_5297),
.Y(n_8162)
);

AO21x2_ASAP7_75t_L g8163 ( 
.A1(n_7618),
.A2(n_6203),
.B(n_6571),
.Y(n_8163)
);

AND2x2_ASAP7_75t_L g8164 ( 
.A(n_7680),
.B(n_5833),
.Y(n_8164)
);

AOI221xp5_ASAP7_75t_L g8165 ( 
.A1(n_7843),
.A2(n_6571),
.B1(n_6562),
.B2(n_6618),
.C(n_6597),
.Y(n_8165)
);

AND2x2_ASAP7_75t_L g8166 ( 
.A(n_7700),
.B(n_5833),
.Y(n_8166)
);

OAI211xp5_ASAP7_75t_L g8167 ( 
.A1(n_7878),
.A2(n_5736),
.B(n_5608),
.C(n_5368),
.Y(n_8167)
);

NOR3xp33_ASAP7_75t_L g8168 ( 
.A(n_7747),
.B(n_5318),
.C(n_5297),
.Y(n_8168)
);

AND2x2_ASAP7_75t_L g8169 ( 
.A(n_7701),
.B(n_5860),
.Y(n_8169)
);

NAND3xp33_ASAP7_75t_L g8170 ( 
.A(n_7722),
.B(n_6249),
.C(n_5964),
.Y(n_8170)
);

NAND4xp75_ASAP7_75t_L g8171 ( 
.A(n_7681),
.B(n_6401),
.C(n_6493),
.D(n_6359),
.Y(n_8171)
);

AND2x2_ASAP7_75t_L g8172 ( 
.A(n_7710),
.B(n_5860),
.Y(n_8172)
);

NOR2x1_ASAP7_75t_L g8173 ( 
.A(n_7808),
.B(n_6203),
.Y(n_8173)
);

NOR2x1_ASAP7_75t_L g8174 ( 
.A(n_7811),
.B(n_6203),
.Y(n_8174)
);

BUFx2_ASAP7_75t_L g8175 ( 
.A(n_7819),
.Y(n_8175)
);

NAND2xp5_ASAP7_75t_SL g8176 ( 
.A(n_7776),
.B(n_6025),
.Y(n_8176)
);

AOI22xp33_ASAP7_75t_SL g8177 ( 
.A1(n_7735),
.A2(n_4918),
.B1(n_4942),
.B2(n_5195),
.Y(n_8177)
);

NAND3xp33_ASAP7_75t_L g8178 ( 
.A(n_7750),
.B(n_4911),
.C(n_4872),
.Y(n_8178)
);

NAND2xp5_ASAP7_75t_L g8179 ( 
.A(n_7725),
.B(n_6048),
.Y(n_8179)
);

NOR3xp33_ASAP7_75t_L g8180 ( 
.A(n_7756),
.B(n_7763),
.C(n_7759),
.Y(n_8180)
);

OR2x2_ASAP7_75t_L g8181 ( 
.A(n_7804),
.B(n_5518),
.Y(n_8181)
);

NOR2xp33_ASAP7_75t_L g8182 ( 
.A(n_7705),
.B(n_5784),
.Y(n_8182)
);

AOI22xp33_ASAP7_75t_L g8183 ( 
.A1(n_7843),
.A2(n_4905),
.B1(n_6618),
.B2(n_6597),
.Y(n_8183)
);

NAND2xp5_ASAP7_75t_L g8184 ( 
.A(n_7726),
.B(n_7732),
.Y(n_8184)
);

NAND2xp5_ASAP7_75t_L g8185 ( 
.A(n_7736),
.B(n_6048),
.Y(n_8185)
);

NAND2xp5_ASAP7_75t_L g8186 ( 
.A(n_7742),
.B(n_6048),
.Y(n_8186)
);

INVx2_ASAP7_75t_L g8187 ( 
.A(n_7762),
.Y(n_8187)
);

AOI22xp33_ASAP7_75t_L g8188 ( 
.A1(n_7781),
.A2(n_4905),
.B1(n_6562),
.B2(n_4918),
.Y(n_8188)
);

AND2x2_ASAP7_75t_L g8189 ( 
.A(n_7823),
.B(n_7824),
.Y(n_8189)
);

NAND4xp75_ASAP7_75t_L g8190 ( 
.A(n_7752),
.B(n_6549),
.C(n_6401),
.D(n_6493),
.Y(n_8190)
);

AND2x2_ASAP7_75t_L g8191 ( 
.A(n_7880),
.B(n_6029),
.Y(n_8191)
);

BUFx3_ASAP7_75t_L g8192 ( 
.A(n_7614),
.Y(n_8192)
);

INVx2_ASAP7_75t_L g8193 ( 
.A(n_7788),
.Y(n_8193)
);

AND2x2_ASAP7_75t_L g8194 ( 
.A(n_7691),
.B(n_6029),
.Y(n_8194)
);

INVx1_ASAP7_75t_L g8195 ( 
.A(n_7811),
.Y(n_8195)
);

NAND2xp5_ASAP7_75t_L g8196 ( 
.A(n_7712),
.B(n_6053),
.Y(n_8196)
);

AOI221x1_ASAP7_75t_SL g8197 ( 
.A1(n_7782),
.A2(n_6133),
.B1(n_6140),
.B2(n_6122),
.C(n_6117),
.Y(n_8197)
);

AO21x2_ASAP7_75t_L g8198 ( 
.A1(n_7624),
.A2(n_6446),
.B(n_6122),
.Y(n_8198)
);

NAND2xp5_ASAP7_75t_L g8199 ( 
.A(n_7731),
.B(n_6053),
.Y(n_8199)
);

NOR3xp33_ASAP7_75t_L g8200 ( 
.A(n_7783),
.B(n_5318),
.C(n_5297),
.Y(n_8200)
);

NAND3xp33_ASAP7_75t_L g8201 ( 
.A(n_7784),
.B(n_4911),
.C(n_4872),
.Y(n_8201)
);

NAND4xp75_ASAP7_75t_L g8202 ( 
.A(n_7718),
.B(n_6493),
.C(n_6549),
.D(n_6359),
.Y(n_8202)
);

AOI22xp33_ASAP7_75t_L g8203 ( 
.A1(n_7867),
.A2(n_4905),
.B1(n_5034),
.B2(n_4944),
.Y(n_8203)
);

NAND3xp33_ASAP7_75t_L g8204 ( 
.A(n_7651),
.B(n_4983),
.C(n_4939),
.Y(n_8204)
);

AND2x2_ASAP7_75t_L g8205 ( 
.A(n_7805),
.B(n_6041),
.Y(n_8205)
);

AND2x2_ASAP7_75t_L g8206 ( 
.A(n_7825),
.B(n_6041),
.Y(n_8206)
);

AND2x2_ASAP7_75t_L g8207 ( 
.A(n_7827),
.B(n_5784),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_7813),
.Y(n_8208)
);

AND2x2_ASAP7_75t_L g8209 ( 
.A(n_7832),
.B(n_5784),
.Y(n_8209)
);

NAND3xp33_ASAP7_75t_L g8210 ( 
.A(n_7817),
.B(n_4983),
.C(n_4939),
.Y(n_8210)
);

INVx2_ASAP7_75t_L g8211 ( 
.A(n_8019),
.Y(n_8211)
);

OAI211xp5_ASAP7_75t_SL g8212 ( 
.A1(n_8099),
.A2(n_7870),
.B(n_7881),
.C(n_7872),
.Y(n_8212)
);

INVx1_ASAP7_75t_L g8213 ( 
.A(n_8120),
.Y(n_8213)
);

AOI22xp33_ASAP7_75t_L g8214 ( 
.A1(n_8147),
.A2(n_7689),
.B1(n_7699),
.B2(n_7697),
.Y(n_8214)
);

AOI22xp33_ASAP7_75t_L g8215 ( 
.A1(n_7901),
.A2(n_7706),
.B1(n_7707),
.B2(n_7867),
.Y(n_8215)
);

INVx2_ASAP7_75t_L g8216 ( 
.A(n_7912),
.Y(n_8216)
);

INVx4_ASAP7_75t_L g8217 ( 
.A(n_8110),
.Y(n_8217)
);

AND2x4_ASAP7_75t_SL g8218 ( 
.A(n_7976),
.B(n_7912),
.Y(n_8218)
);

AND2x2_ASAP7_75t_L g8219 ( 
.A(n_7911),
.B(n_7844),
.Y(n_8219)
);

AOI221xp5_ASAP7_75t_L g8220 ( 
.A1(n_7954),
.A2(n_7872),
.B1(n_7882),
.B2(n_7881),
.C(n_7870),
.Y(n_8220)
);

AND2x4_ASAP7_75t_L g8221 ( 
.A(n_8133),
.B(n_7617),
.Y(n_8221)
);

INVx1_ASAP7_75t_L g8222 ( 
.A(n_8175),
.Y(n_8222)
);

INVx1_ASAP7_75t_L g8223 ( 
.A(n_8054),
.Y(n_8223)
);

HB1xp67_ASAP7_75t_L g8224 ( 
.A(n_8105),
.Y(n_8224)
);

INVx2_ASAP7_75t_L g8225 ( 
.A(n_7986),
.Y(n_8225)
);

INVx1_ASAP7_75t_SL g8226 ( 
.A(n_8135),
.Y(n_8226)
);

OAI31xp33_ASAP7_75t_L g8227 ( 
.A1(n_8167),
.A2(n_7748),
.A3(n_7802),
.B(n_7845),
.Y(n_8227)
);

AND2x2_ASAP7_75t_L g8228 ( 
.A(n_7907),
.B(n_7850),
.Y(n_8228)
);

AND2x2_ASAP7_75t_L g8229 ( 
.A(n_7903),
.B(n_7876),
.Y(n_8229)
);

NAND2x1p5_ASAP7_75t_L g8230 ( 
.A(n_7969),
.B(n_7693),
.Y(n_8230)
);

INVx2_ASAP7_75t_L g8231 ( 
.A(n_8003),
.Y(n_8231)
);

INVx1_ASAP7_75t_L g8232 ( 
.A(n_8054),
.Y(n_8232)
);

NOR2xp33_ASAP7_75t_L g8233 ( 
.A(n_7893),
.B(n_7882),
.Y(n_8233)
);

INVx1_ASAP7_75t_L g8234 ( 
.A(n_8076),
.Y(n_8234)
);

INVx1_ASAP7_75t_L g8235 ( 
.A(n_8076),
.Y(n_8235)
);

INVx2_ASAP7_75t_SL g8236 ( 
.A(n_7909),
.Y(n_8236)
);

AND2x2_ASAP7_75t_L g8237 ( 
.A(n_7928),
.B(n_7877),
.Y(n_8237)
);

AOI322xp5_ASAP7_75t_L g8238 ( 
.A1(n_7925),
.A2(n_7830),
.A3(n_7835),
.B1(n_7831),
.B2(n_7733),
.C1(n_7724),
.C2(n_7723),
.Y(n_8238)
);

OAI22xp5_ASAP7_75t_L g8239 ( 
.A1(n_7894),
.A2(n_7860),
.B1(n_7884),
.B2(n_7842),
.Y(n_8239)
);

AND2x2_ASAP7_75t_L g8240 ( 
.A(n_7967),
.B(n_7830),
.Y(n_8240)
);

NAND2xp5_ASAP7_75t_L g8241 ( 
.A(n_8060),
.B(n_7885),
.Y(n_8241)
);

AND2x2_ASAP7_75t_L g8242 ( 
.A(n_8007),
.B(n_7831),
.Y(n_8242)
);

OR2x2_ASAP7_75t_L g8243 ( 
.A(n_7905),
.B(n_7835),
.Y(n_8243)
);

INVx4_ASAP7_75t_L g8244 ( 
.A(n_8110),
.Y(n_8244)
);

INVx2_ASAP7_75t_L g8245 ( 
.A(n_7900),
.Y(n_8245)
);

INVx2_ASAP7_75t_SL g8246 ( 
.A(n_7909),
.Y(n_8246)
);

AND2x2_ASAP7_75t_L g8247 ( 
.A(n_7921),
.B(n_7847),
.Y(n_8247)
);

INVx2_ASAP7_75t_L g8248 ( 
.A(n_7946),
.Y(n_8248)
);

INVx1_ASAP7_75t_L g8249 ( 
.A(n_8084),
.Y(n_8249)
);

OAI221xp5_ASAP7_75t_L g8250 ( 
.A1(n_7982),
.A2(n_7879),
.B1(n_7874),
.B2(n_7851),
.C(n_7852),
.Y(n_8250)
);

OR2x2_ASAP7_75t_L g8251 ( 
.A(n_7951),
.B(n_7847),
.Y(n_8251)
);

OR2x2_ASAP7_75t_L g8252 ( 
.A(n_7913),
.B(n_7848),
.Y(n_8252)
);

AND2x2_ASAP7_75t_L g8253 ( 
.A(n_7933),
.B(n_7848),
.Y(n_8253)
);

AOI222xp33_ASAP7_75t_L g8254 ( 
.A1(n_7898),
.A2(n_7818),
.B1(n_7821),
.B2(n_7820),
.C1(n_7813),
.C2(n_7851),
.Y(n_8254)
);

AND2x2_ASAP7_75t_L g8255 ( 
.A(n_7960),
.B(n_7852),
.Y(n_8255)
);

AOI221x1_ASAP7_75t_L g8256 ( 
.A1(n_8107),
.A2(n_7735),
.B1(n_7821),
.B2(n_7820),
.C(n_7818),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7891),
.Y(n_8257)
);

HB1xp67_ASAP7_75t_L g8258 ( 
.A(n_8105),
.Y(n_8258)
);

INVx1_ASAP7_75t_L g8259 ( 
.A(n_7904),
.Y(n_8259)
);

OAI31xp33_ASAP7_75t_L g8260 ( 
.A1(n_8043),
.A2(n_7861),
.A3(n_7856),
.B(n_5184),
.Y(n_8260)
);

HB1xp67_ASAP7_75t_L g8261 ( 
.A(n_7972),
.Y(n_8261)
);

NAND2xp5_ASAP7_75t_L g8262 ( 
.A(n_7920),
.B(n_7856),
.Y(n_8262)
);

INVx1_ASAP7_75t_L g8263 ( 
.A(n_7972),
.Y(n_8263)
);

NAND3xp33_ASAP7_75t_SL g8264 ( 
.A(n_7931),
.B(n_7861),
.C(n_7704),
.Y(n_8264)
);

AND2x2_ASAP7_75t_L g8265 ( 
.A(n_7939),
.B(n_7873),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_8189),
.Y(n_8266)
);

NAND2xp5_ASAP7_75t_L g8267 ( 
.A(n_8151),
.B(n_7883),
.Y(n_8267)
);

AND2x2_ASAP7_75t_L g8268 ( 
.A(n_7935),
.B(n_7542),
.Y(n_8268)
);

AND2x2_ASAP7_75t_L g8269 ( 
.A(n_8021),
.B(n_7554),
.Y(n_8269)
);

AND2x2_ASAP7_75t_SL g8270 ( 
.A(n_7899),
.B(n_7593),
.Y(n_8270)
);

INVx1_ASAP7_75t_L g8271 ( 
.A(n_8092),
.Y(n_8271)
);

NAND2x1_ASAP7_75t_L g8272 ( 
.A(n_7946),
.B(n_7593),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_8092),
.Y(n_8273)
);

INVx1_ASAP7_75t_L g8274 ( 
.A(n_7908),
.Y(n_8274)
);

INVx1_ASAP7_75t_L g8275 ( 
.A(n_8120),
.Y(n_8275)
);

INVx1_ASAP7_75t_SL g8276 ( 
.A(n_8083),
.Y(n_8276)
);

HB1xp67_ASAP7_75t_L g8277 ( 
.A(n_8040),
.Y(n_8277)
);

AND2x2_ASAP7_75t_L g8278 ( 
.A(n_7952),
.B(n_7875),
.Y(n_8278)
);

INVx2_ASAP7_75t_L g8279 ( 
.A(n_8036),
.Y(n_8279)
);

INVx2_ASAP7_75t_L g8280 ( 
.A(n_7886),
.Y(n_8280)
);

NAND2xp5_ASAP7_75t_SL g8281 ( 
.A(n_8064),
.B(n_6025),
.Y(n_8281)
);

AND2x2_ASAP7_75t_L g8282 ( 
.A(n_7963),
.B(n_8008),
.Y(n_8282)
);

INVx2_ASAP7_75t_L g8283 ( 
.A(n_7949),
.Y(n_8283)
);

INVx1_ASAP7_75t_L g8284 ( 
.A(n_7942),
.Y(n_8284)
);

BUFx3_ASAP7_75t_L g8285 ( 
.A(n_7902),
.Y(n_8285)
);

AND2x4_ASAP7_75t_L g8286 ( 
.A(n_8085),
.B(n_7612),
.Y(n_8286)
);

BUFx2_ASAP7_75t_L g8287 ( 
.A(n_8073),
.Y(n_8287)
);

NAND4xp25_ASAP7_75t_L g8288 ( 
.A(n_7906),
.B(n_7957),
.C(n_7890),
.D(n_7955),
.Y(n_8288)
);

INVx4_ASAP7_75t_L g8289 ( 
.A(n_7965),
.Y(n_8289)
);

INVx1_ASAP7_75t_L g8290 ( 
.A(n_7929),
.Y(n_8290)
);

NAND2xp5_ASAP7_75t_L g8291 ( 
.A(n_8002),
.B(n_7716),
.Y(n_8291)
);

HB1xp67_ASAP7_75t_L g8292 ( 
.A(n_7973),
.Y(n_8292)
);

INVx3_ASAP7_75t_L g8293 ( 
.A(n_8097),
.Y(n_8293)
);

OR2x2_ASAP7_75t_L g8294 ( 
.A(n_7889),
.B(n_7609),
.Y(n_8294)
);

AND2x2_ASAP7_75t_L g8295 ( 
.A(n_7993),
.B(n_7609),
.Y(n_8295)
);

NOR4xp25_ASAP7_75t_L g8296 ( 
.A(n_7937),
.B(n_7741),
.C(n_7753),
.D(n_7798),
.Y(n_8296)
);

NAND3xp33_ASAP7_75t_L g8297 ( 
.A(n_7966),
.B(n_7778),
.C(n_7734),
.Y(n_8297)
);

AND2x2_ASAP7_75t_L g8298 ( 
.A(n_7990),
.B(n_7675),
.Y(n_8298)
);

AND2x4_ASAP7_75t_L g8299 ( 
.A(n_8085),
.B(n_5801),
.Y(n_8299)
);

INVx2_ASAP7_75t_L g8300 ( 
.A(n_8097),
.Y(n_8300)
);

INVx1_ASAP7_75t_SL g8301 ( 
.A(n_8028),
.Y(n_8301)
);

INVx1_ASAP7_75t_SL g8302 ( 
.A(n_8056),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7932),
.Y(n_8303)
);

INVx2_ASAP7_75t_L g8304 ( 
.A(n_8103),
.Y(n_8304)
);

AOI22xp5_ASAP7_75t_SL g8305 ( 
.A1(n_7936),
.A2(n_7778),
.B1(n_7734),
.B2(n_7791),
.Y(n_8305)
);

HB1xp67_ASAP7_75t_L g8306 ( 
.A(n_7973),
.Y(n_8306)
);

INVx3_ASAP7_75t_L g8307 ( 
.A(n_8103),
.Y(n_8307)
);

HB1xp67_ASAP7_75t_L g8308 ( 
.A(n_7988),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_7992),
.B(n_7675),
.Y(n_8309)
);

NAND4xp25_ASAP7_75t_L g8310 ( 
.A(n_7895),
.B(n_5024),
.C(n_5369),
.D(n_4894),
.Y(n_8310)
);

AND2x2_ASAP7_75t_L g8311 ( 
.A(n_7971),
.B(n_7862),
.Y(n_8311)
);

INVx4_ASAP7_75t_L g8312 ( 
.A(n_8001),
.Y(n_8312)
);

OAI221xp5_ASAP7_75t_L g8313 ( 
.A1(n_8134),
.A2(n_7791),
.B1(n_5208),
.B2(n_5233),
.C(n_5195),
.Y(n_8313)
);

INVxp67_ASAP7_75t_SL g8314 ( 
.A(n_7927),
.Y(n_8314)
);

INVx1_ASAP7_75t_L g8315 ( 
.A(n_7924),
.Y(n_8315)
);

AND2x2_ASAP7_75t_L g8316 ( 
.A(n_7979),
.B(n_7862),
.Y(n_8316)
);

HB1xp67_ASAP7_75t_L g8317 ( 
.A(n_7991),
.Y(n_8317)
);

AND2x2_ASAP7_75t_L g8318 ( 
.A(n_7994),
.B(n_7868),
.Y(n_8318)
);

BUFx2_ASAP7_75t_L g8319 ( 
.A(n_8055),
.Y(n_8319)
);

INVx1_ASAP7_75t_L g8320 ( 
.A(n_7943),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_7968),
.Y(n_8321)
);

NAND3xp33_ASAP7_75t_L g8322 ( 
.A(n_8046),
.B(n_7868),
.C(n_7840),
.Y(n_8322)
);

OR2x2_ASAP7_75t_L g8323 ( 
.A(n_7918),
.B(n_7840),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_8035),
.Y(n_8324)
);

AND2x4_ASAP7_75t_L g8325 ( 
.A(n_8020),
.B(n_5801),
.Y(n_8325)
);

AND2x4_ASAP7_75t_L g8326 ( 
.A(n_8053),
.B(n_5801),
.Y(n_8326)
);

NAND3xp33_ASAP7_75t_SL g8327 ( 
.A(n_7931),
.B(n_5526),
.C(n_5430),
.Y(n_8327)
);

HB1xp67_ASAP7_75t_L g8328 ( 
.A(n_7930),
.Y(n_8328)
);

AND2x2_ASAP7_75t_L g8329 ( 
.A(n_7995),
.B(n_5687),
.Y(n_8329)
);

NAND2xp5_ASAP7_75t_L g8330 ( 
.A(n_8153),
.B(n_8000),
.Y(n_8330)
);

OAI31xp33_ASAP7_75t_SL g8331 ( 
.A1(n_8114),
.A2(n_6006),
.A3(n_6422),
.B(n_6291),
.Y(n_8331)
);

AOI22xp33_ASAP7_75t_L g8332 ( 
.A1(n_7983),
.A2(n_5233),
.B1(n_5208),
.B2(n_5330),
.Y(n_8332)
);

INVx1_ASAP7_75t_L g8333 ( 
.A(n_8068),
.Y(n_8333)
);

NAND2xp5_ASAP7_75t_SL g8334 ( 
.A(n_8032),
.B(n_6025),
.Y(n_8334)
);

INVx1_ASAP7_75t_SL g8335 ( 
.A(n_8146),
.Y(n_8335)
);

INVx1_ASAP7_75t_L g8336 ( 
.A(n_8079),
.Y(n_8336)
);

AND2x4_ASAP7_75t_L g8337 ( 
.A(n_8027),
.B(n_5801),
.Y(n_8337)
);

AND2x4_ASAP7_75t_L g8338 ( 
.A(n_8037),
.B(n_8192),
.Y(n_8338)
);

AND2x2_ASAP7_75t_L g8339 ( 
.A(n_7945),
.B(n_5687),
.Y(n_8339)
);

INVx1_ASAP7_75t_L g8340 ( 
.A(n_8081),
.Y(n_8340)
);

AND2x2_ASAP7_75t_L g8341 ( 
.A(n_7940),
.B(n_5803),
.Y(n_8341)
);

OR2x2_ASAP7_75t_L g8342 ( 
.A(n_7959),
.B(n_6117),
.Y(n_8342)
);

AND2x2_ASAP7_75t_L g8343 ( 
.A(n_7953),
.B(n_5803),
.Y(n_8343)
);

BUFx2_ASAP7_75t_L g8344 ( 
.A(n_8136),
.Y(n_8344)
);

INVx3_ASAP7_75t_L g8345 ( 
.A(n_8149),
.Y(n_8345)
);

BUFx12f_ASAP7_75t_L g8346 ( 
.A(n_7897),
.Y(n_8346)
);

AND2x2_ASAP7_75t_L g8347 ( 
.A(n_8152),
.B(n_5858),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_8087),
.Y(n_8348)
);

AND2x2_ASAP7_75t_L g8349 ( 
.A(n_8138),
.B(n_5858),
.Y(n_8349)
);

AOI33xp33_ASAP7_75t_L g8350 ( 
.A1(n_7910),
.A2(n_5362),
.A3(n_5342),
.B1(n_5338),
.B2(n_5421),
.B3(n_6133),
.Y(n_8350)
);

INVx1_ASAP7_75t_L g8351 ( 
.A(n_8093),
.Y(n_8351)
);

AOI21xp5_ASAP7_75t_SL g8352 ( 
.A1(n_7887),
.A2(n_5208),
.B(n_5233),
.Y(n_8352)
);

OR2x6_ASAP7_75t_L g8353 ( 
.A(n_7888),
.B(n_3742),
.Y(n_8353)
);

INVx2_ASAP7_75t_L g8354 ( 
.A(n_8161),
.Y(n_8354)
);

INVx2_ASAP7_75t_L g8355 ( 
.A(n_8164),
.Y(n_8355)
);

AND2x2_ASAP7_75t_L g8356 ( 
.A(n_7944),
.B(n_5671),
.Y(n_8356)
);

NAND2xp5_ASAP7_75t_L g8357 ( 
.A(n_8116),
.B(n_8132),
.Y(n_8357)
);

OR2x2_ASAP7_75t_L g8358 ( 
.A(n_7964),
.B(n_6140),
.Y(n_8358)
);

INVx1_ASAP7_75t_L g8359 ( 
.A(n_7942),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_8173),
.Y(n_8360)
);

HB1xp67_ASAP7_75t_L g8361 ( 
.A(n_7916),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_8115),
.Y(n_8362)
);

AND2x2_ASAP7_75t_L g8363 ( 
.A(n_7948),
.B(n_5671),
.Y(n_8363)
);

AND2x4_ASAP7_75t_L g8364 ( 
.A(n_7892),
.B(n_5808),
.Y(n_8364)
);

OR2x2_ASAP7_75t_L g8365 ( 
.A(n_8004),
.B(n_6142),
.Y(n_8365)
);

NAND2xp5_ASAP7_75t_L g8366 ( 
.A(n_8144),
.B(n_6053),
.Y(n_8366)
);

NAND2xp5_ASAP7_75t_L g8367 ( 
.A(n_7896),
.B(n_7922),
.Y(n_8367)
);

OAI33xp33_ASAP7_75t_L g8368 ( 
.A1(n_7997),
.A2(n_6172),
.A3(n_6153),
.B1(n_6174),
.B2(n_6169),
.B3(n_6142),
.Y(n_8368)
);

NAND2xp5_ASAP7_75t_L g8369 ( 
.A(n_7941),
.B(n_6053),
.Y(n_8369)
);

BUFx2_ASAP7_75t_L g8370 ( 
.A(n_7917),
.Y(n_8370)
);

OAI221xp5_ASAP7_75t_L g8371 ( 
.A1(n_7981),
.A2(n_5733),
.B1(n_5808),
.B2(n_5076),
.C(n_5207),
.Y(n_8371)
);

NAND2xp5_ASAP7_75t_L g8372 ( 
.A(n_8050),
.B(n_6153),
.Y(n_8372)
);

AND2x2_ASAP7_75t_L g8373 ( 
.A(n_8141),
.B(n_5683),
.Y(n_8373)
);

OAI33xp33_ASAP7_75t_L g8374 ( 
.A1(n_7984),
.A2(n_6175),
.A3(n_6172),
.B1(n_6178),
.B2(n_6174),
.B3(n_6169),
.Y(n_8374)
);

AOI221xp5_ASAP7_75t_L g8375 ( 
.A1(n_8197),
.A2(n_6446),
.B1(n_6256),
.B2(n_6247),
.C(n_6235),
.Y(n_8375)
);

OAI22xp5_ASAP7_75t_L g8376 ( 
.A1(n_7961),
.A2(n_5808),
.B1(n_5733),
.B2(n_5722),
.Y(n_8376)
);

INVx2_ASAP7_75t_SL g8377 ( 
.A(n_7958),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_8080),
.Y(n_8378)
);

AOI33xp33_ASAP7_75t_L g8379 ( 
.A1(n_7998),
.A2(n_6182),
.A3(n_6178),
.B1(n_6194),
.B2(n_6193),
.B3(n_6175),
.Y(n_8379)
);

AOI221x1_ASAP7_75t_L g8380 ( 
.A1(n_8108),
.A2(n_6193),
.B1(n_6195),
.B2(n_6194),
.C(n_6182),
.Y(n_8380)
);

AND2x4_ASAP7_75t_L g8381 ( 
.A(n_8098),
.B(n_5808),
.Y(n_8381)
);

BUFx2_ASAP7_75t_L g8382 ( 
.A(n_7978),
.Y(n_8382)
);

INVx2_ASAP7_75t_SL g8383 ( 
.A(n_8045),
.Y(n_8383)
);

AND2x2_ASAP7_75t_L g8384 ( 
.A(n_8123),
.B(n_5683),
.Y(n_8384)
);

OAI21xp5_ASAP7_75t_L g8385 ( 
.A1(n_8109),
.A2(n_5920),
.B(n_5878),
.Y(n_8385)
);

AND2x2_ASAP7_75t_L g8386 ( 
.A(n_8072),
.B(n_5870),
.Y(n_8386)
);

OR2x2_ASAP7_75t_L g8387 ( 
.A(n_7938),
.B(n_6195),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_8140),
.Y(n_8388)
);

AND2x4_ASAP7_75t_L g8389 ( 
.A(n_8029),
.B(n_5722),
.Y(n_8389)
);

INVx2_ASAP7_75t_L g8390 ( 
.A(n_8187),
.Y(n_8390)
);

AND2x2_ASAP7_75t_L g8391 ( 
.A(n_8169),
.B(n_5870),
.Y(n_8391)
);

AOI22xp33_ASAP7_75t_L g8392 ( 
.A1(n_7983),
.A2(n_5381),
.B1(n_5330),
.B2(n_4939),
.Y(n_8392)
);

HB1xp67_ASAP7_75t_L g8393 ( 
.A(n_7916),
.Y(n_8393)
);

OR2x2_ASAP7_75t_L g8394 ( 
.A(n_7919),
.B(n_6214),
.Y(n_8394)
);

NOR2xp67_ASAP7_75t_SL g8395 ( 
.A(n_7926),
.B(n_3742),
.Y(n_8395)
);

NAND2xp5_ASAP7_75t_L g8396 ( 
.A(n_7947),
.B(n_6214),
.Y(n_8396)
);

NAND2xp5_ASAP7_75t_L g8397 ( 
.A(n_8052),
.B(n_6216),
.Y(n_8397)
);

AND2x2_ASAP7_75t_L g8398 ( 
.A(n_8172),
.B(n_5914),
.Y(n_8398)
);

HB1xp67_ASAP7_75t_L g8399 ( 
.A(n_8082),
.Y(n_8399)
);

OAI211xp5_ASAP7_75t_L g8400 ( 
.A1(n_8177),
.A2(n_5736),
.B(n_5608),
.C(n_5330),
.Y(n_8400)
);

HB1xp67_ASAP7_75t_L g8401 ( 
.A(n_8094),
.Y(n_8401)
);

INVx1_ASAP7_75t_L g8402 ( 
.A(n_8142),
.Y(n_8402)
);

HB1xp67_ASAP7_75t_L g8403 ( 
.A(n_7934),
.Y(n_8403)
);

AND2x4_ASAP7_75t_L g8404 ( 
.A(n_7915),
.B(n_5722),
.Y(n_8404)
);

OAI31xp33_ASAP7_75t_SL g8405 ( 
.A1(n_8119),
.A2(n_6422),
.A3(n_6291),
.B(n_6243),
.Y(n_8405)
);

INVx2_ASAP7_75t_L g8406 ( 
.A(n_8086),
.Y(n_8406)
);

INVx1_ASAP7_75t_L g8407 ( 
.A(n_8173),
.Y(n_8407)
);

NAND2xp5_ASAP7_75t_SL g8408 ( 
.A(n_7977),
.B(n_6025),
.Y(n_8408)
);

INVx4_ASAP7_75t_L g8409 ( 
.A(n_8131),
.Y(n_8409)
);

AND2x2_ASAP7_75t_L g8410 ( 
.A(n_8047),
.B(n_5914),
.Y(n_8410)
);

NOR3xp33_ASAP7_75t_L g8411 ( 
.A(n_8204),
.B(n_8210),
.C(n_8139),
.Y(n_8411)
);

INVx2_ASAP7_75t_L g8412 ( 
.A(n_8193),
.Y(n_8412)
);

INVx5_ASAP7_75t_L g8413 ( 
.A(n_8044),
.Y(n_8413)
);

INVx6_ASAP7_75t_L g8414 ( 
.A(n_7987),
.Y(n_8414)
);

AND2x4_ASAP7_75t_L g8415 ( 
.A(n_8034),
.B(n_5722),
.Y(n_8415)
);

AOI22xp5_ASAP7_75t_L g8416 ( 
.A1(n_8182),
.A2(n_5347),
.B1(n_5381),
.B2(n_5330),
.Y(n_8416)
);

INVx2_ASAP7_75t_L g8417 ( 
.A(n_8074),
.Y(n_8417)
);

INVx1_ASAP7_75t_L g8418 ( 
.A(n_8143),
.Y(n_8418)
);

INVx1_ASAP7_75t_L g8419 ( 
.A(n_8145),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_8148),
.Y(n_8420)
);

INVx1_ASAP7_75t_L g8421 ( 
.A(n_8195),
.Y(n_8421)
);

CKINVDCx16_ASAP7_75t_R g8422 ( 
.A(n_7980),
.Y(n_8422)
);

INVxp67_ASAP7_75t_SL g8423 ( 
.A(n_8016),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_8174),
.Y(n_8424)
);

NAND2xp5_ASAP7_75t_L g8425 ( 
.A(n_7962),
.B(n_6216),
.Y(n_8425)
);

NAND3xp33_ASAP7_75t_L g8426 ( 
.A(n_7923),
.B(n_4983),
.C(n_4939),
.Y(n_8426)
);

AND2x4_ASAP7_75t_L g8427 ( 
.A(n_8208),
.B(n_6027),
.Y(n_8427)
);

INVx3_ASAP7_75t_L g8428 ( 
.A(n_8191),
.Y(n_8428)
);

NAND2xp5_ASAP7_75t_SL g8429 ( 
.A(n_8063),
.B(n_6027),
.Y(n_8429)
);

AND2x2_ASAP7_75t_L g8430 ( 
.A(n_8051),
.B(n_5916),
.Y(n_8430)
);

NAND2xp5_ASAP7_75t_L g8431 ( 
.A(n_8137),
.B(n_6227),
.Y(n_8431)
);

OAI21xp5_ASAP7_75t_L g8432 ( 
.A1(n_8022),
.A2(n_5920),
.B(n_5857),
.Y(n_8432)
);

NOR2xp67_ASAP7_75t_L g8433 ( 
.A(n_8067),
.B(n_6227),
.Y(n_8433)
);

OAI33xp33_ASAP7_75t_L g8434 ( 
.A1(n_7989),
.A2(n_6259),
.A3(n_6253),
.B1(n_6276),
.B2(n_6255),
.B3(n_6252),
.Y(n_8434)
);

OR2x2_ASAP7_75t_L g8435 ( 
.A(n_8184),
.B(n_6252),
.Y(n_8435)
);

INVx2_ASAP7_75t_L g8436 ( 
.A(n_8095),
.Y(n_8436)
);

INVx2_ASAP7_75t_L g8437 ( 
.A(n_8194),
.Y(n_8437)
);

AND2x2_ASAP7_75t_L g8438 ( 
.A(n_8166),
.B(n_5916),
.Y(n_8438)
);

INVx1_ASAP7_75t_L g8439 ( 
.A(n_8042),
.Y(n_8439)
);

OAI22xp5_ASAP7_75t_L g8440 ( 
.A1(n_8058),
.A2(n_8066),
.B1(n_7914),
.B2(n_8090),
.Y(n_8440)
);

AOI21xp5_ASAP7_75t_L g8441 ( 
.A1(n_7887),
.A2(n_6446),
.B(n_6255),
.Y(n_8441)
);

INVx2_ASAP7_75t_L g8442 ( 
.A(n_8102),
.Y(n_8442)
);

OR2x2_ASAP7_75t_L g8443 ( 
.A(n_8014),
.B(n_6253),
.Y(n_8443)
);

NAND2xp5_ASAP7_75t_L g8444 ( 
.A(n_8005),
.B(n_6259),
.Y(n_8444)
);

INVx2_ASAP7_75t_L g8445 ( 
.A(n_8118),
.Y(n_8445)
);

NAND2xp5_ASAP7_75t_L g8446 ( 
.A(n_8062),
.B(n_6276),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_8017),
.Y(n_8447)
);

HB1xp67_ASAP7_75t_L g8448 ( 
.A(n_7970),
.Y(n_8448)
);

OR2x2_ASAP7_75t_L g8449 ( 
.A(n_7985),
.B(n_6279),
.Y(n_8449)
);

NAND2xp5_ASAP7_75t_L g8450 ( 
.A(n_7956),
.B(n_6279),
.Y(n_8450)
);

AND2x4_ASAP7_75t_SL g8451 ( 
.A(n_8104),
.B(n_5381),
.Y(n_8451)
);

AOI222xp33_ASAP7_75t_L g8452 ( 
.A1(n_7999),
.A2(n_4568),
.B1(n_5198),
.B2(n_5209),
.C1(n_4983),
.C2(n_5401),
.Y(n_8452)
);

INVx5_ASAP7_75t_L g8453 ( 
.A(n_8069),
.Y(n_8453)
);

OAI31xp33_ASAP7_75t_SL g8454 ( 
.A1(n_8038),
.A2(n_6243),
.A3(n_5097),
.B(n_5261),
.Y(n_8454)
);

INVx1_ASAP7_75t_L g8455 ( 
.A(n_8026),
.Y(n_8455)
);

NAND2xp5_ASAP7_75t_L g8456 ( 
.A(n_8059),
.B(n_6281),
.Y(n_8456)
);

AND2x2_ASAP7_75t_L g8457 ( 
.A(n_8113),
.B(n_5922),
.Y(n_8457)
);

AND2x4_ASAP7_75t_L g8458 ( 
.A(n_8180),
.B(n_6027),
.Y(n_8458)
);

HB1xp67_ASAP7_75t_L g8459 ( 
.A(n_7996),
.Y(n_8459)
);

INVx1_ASAP7_75t_L g8460 ( 
.A(n_8023),
.Y(n_8460)
);

AOI31xp33_ASAP7_75t_SL g8461 ( 
.A1(n_8012),
.A2(n_6281),
.A3(n_6290),
.B(n_6285),
.Y(n_8461)
);

AND2x2_ASAP7_75t_L g8462 ( 
.A(n_8205),
.B(n_5922),
.Y(n_8462)
);

BUFx2_ASAP7_75t_L g8463 ( 
.A(n_8078),
.Y(n_8463)
);

INVx3_ASAP7_75t_L g8464 ( 
.A(n_8207),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_8015),
.Y(n_8465)
);

AND2x4_ASAP7_75t_L g8466 ( 
.A(n_8039),
.B(n_6027),
.Y(n_8466)
);

OR2x2_ASAP7_75t_L g8467 ( 
.A(n_8061),
.B(n_6285),
.Y(n_8467)
);

NAND2xp5_ASAP7_75t_L g8468 ( 
.A(n_8009),
.B(n_6290),
.Y(n_8468)
);

AND2x2_ASAP7_75t_L g8469 ( 
.A(n_8206),
.B(n_5928),
.Y(n_8469)
);

INVx4_ASAP7_75t_L g8470 ( 
.A(n_7950),
.Y(n_8470)
);

AND2x2_ASAP7_75t_L g8471 ( 
.A(n_8033),
.B(n_5928),
.Y(n_8471)
);

OAI33xp33_ASAP7_75t_L g8472 ( 
.A1(n_8048),
.A2(n_6332),
.A3(n_6307),
.B1(n_6338),
.B2(n_6324),
.B3(n_6305),
.Y(n_8472)
);

AND2x2_ASAP7_75t_L g8473 ( 
.A(n_8089),
.B(n_5938),
.Y(n_8473)
);

NAND2xp5_ASAP7_75t_L g8474 ( 
.A(n_7998),
.B(n_6305),
.Y(n_8474)
);

INVx1_ASAP7_75t_L g8475 ( 
.A(n_8025),
.Y(n_8475)
);

AND2x2_ASAP7_75t_L g8476 ( 
.A(n_8065),
.B(n_5938),
.Y(n_8476)
);

HB1xp67_ASAP7_75t_L g8477 ( 
.A(n_8121),
.Y(n_8477)
);

NAND4xp25_ASAP7_75t_L g8478 ( 
.A(n_8178),
.B(n_5063),
.C(n_5038),
.D(n_5224),
.Y(n_8478)
);

AND2x2_ASAP7_75t_L g8479 ( 
.A(n_8106),
.B(n_5975),
.Y(n_8479)
);

NAND3xp33_ASAP7_75t_L g8480 ( 
.A(n_8129),
.B(n_6324),
.C(n_6307),
.Y(n_8480)
);

BUFx2_ASAP7_75t_L g8481 ( 
.A(n_8209),
.Y(n_8481)
);

OR2x2_ASAP7_75t_L g8482 ( 
.A(n_8006),
.B(n_6332),
.Y(n_8482)
);

OAI221xp5_ASAP7_75t_L g8483 ( 
.A1(n_8201),
.A2(n_5204),
.B1(n_5401),
.B2(n_5381),
.C(n_5154),
.Y(n_8483)
);

AOI211xp5_ASAP7_75t_L g8484 ( 
.A1(n_8010),
.A2(n_5378),
.B(n_5388),
.C(n_5286),
.Y(n_8484)
);

INVx2_ASAP7_75t_L g8485 ( 
.A(n_8124),
.Y(n_8485)
);

AND2x4_ASAP7_75t_L g8486 ( 
.A(n_8030),
.B(n_6028),
.Y(n_8486)
);

INVx2_ASAP7_75t_L g8487 ( 
.A(n_8125),
.Y(n_8487)
);

INVx4_ASAP7_75t_L g8488 ( 
.A(n_8126),
.Y(n_8488)
);

AOI222xp33_ASAP7_75t_L g8489 ( 
.A1(n_8057),
.A2(n_5401),
.B1(n_5235),
.B2(n_6033),
.C1(n_6028),
.C2(n_4645),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_8130),
.Y(n_8490)
);

NOR2x1_ASAP7_75t_L g8491 ( 
.A(n_8041),
.B(n_6585),
.Y(n_8491)
);

HB1xp67_ASAP7_75t_L g8492 ( 
.A(n_8088),
.Y(n_8492)
);

INVx1_ASAP7_75t_L g8493 ( 
.A(n_7974),
.Y(n_8493)
);

OAI31xp33_ASAP7_75t_SL g8494 ( 
.A1(n_8049),
.A2(n_6028),
.A3(n_6033),
.B(n_4851),
.Y(n_8494)
);

NAND4xp25_ASAP7_75t_L g8495 ( 
.A(n_8011),
.B(n_3746),
.C(n_3748),
.D(n_5090),
.Y(n_8495)
);

INVx2_ASAP7_75t_L g8496 ( 
.A(n_8181),
.Y(n_8496)
);

INVx2_ASAP7_75t_SL g8497 ( 
.A(n_8196),
.Y(n_8497)
);

AOI33xp33_ASAP7_75t_L g8498 ( 
.A1(n_8075),
.A2(n_6365),
.A3(n_6346),
.B1(n_6367),
.B2(n_6350),
.B3(n_6338),
.Y(n_8498)
);

NAND2xp5_ASAP7_75t_L g8499 ( 
.A(n_8031),
.B(n_6346),
.Y(n_8499)
);

AND2x2_ASAP7_75t_L g8500 ( 
.A(n_8157),
.B(n_5975),
.Y(n_8500)
);

AND2x4_ASAP7_75t_L g8501 ( 
.A(n_7974),
.B(n_6028),
.Y(n_8501)
);

NOR3xp33_ASAP7_75t_SL g8502 ( 
.A(n_8024),
.B(n_5276),
.C(n_4855),
.Y(n_8502)
);

AND2x4_ASAP7_75t_L g8503 ( 
.A(n_7975),
.B(n_6033),
.Y(n_8503)
);

AOI22xp5_ASAP7_75t_L g8504 ( 
.A1(n_8090),
.A2(n_5347),
.B1(n_6033),
.B2(n_5036),
.Y(n_8504)
);

INVx2_ASAP7_75t_L g8505 ( 
.A(n_8198),
.Y(n_8505)
);

AOI322xp5_ASAP7_75t_L g8506 ( 
.A1(n_8013),
.A2(n_8018),
.A3(n_8203),
.B1(n_8174),
.B2(n_8165),
.C1(n_8155),
.C2(n_8070),
.Y(n_8506)
);

OAI33xp33_ASAP7_75t_L g8507 ( 
.A1(n_7975),
.A2(n_6391),
.A3(n_6365),
.B1(n_6397),
.B2(n_6367),
.B3(n_6350),
.Y(n_8507)
);

AOI21xp33_ASAP7_75t_L g8508 ( 
.A1(n_8176),
.A2(n_6397),
.B(n_6391),
.Y(n_8508)
);

AOI211xp5_ASAP7_75t_L g8509 ( 
.A1(n_8162),
.A2(n_4592),
.B(n_5373),
.C(n_5262),
.Y(n_8509)
);

AOI22xp33_ASAP7_75t_L g8510 ( 
.A1(n_8077),
.A2(n_4567),
.B1(n_4976),
.B2(n_4896),
.Y(n_8510)
);

INVx3_ASAP7_75t_L g8511 ( 
.A(n_8217),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8261),
.Y(n_8512)
);

HB1xp67_ASAP7_75t_L g8513 ( 
.A(n_8272),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_8271),
.Y(n_8514)
);

NAND2xp5_ASAP7_75t_L g8515 ( 
.A(n_8422),
.B(n_8013),
.Y(n_8515)
);

A2O1A1O1Ixp25_ASAP7_75t_L g8516 ( 
.A1(n_8250),
.A2(n_8077),
.B(n_8127),
.C(n_8199),
.D(n_8096),
.Y(n_8516)
);

HB1xp67_ASAP7_75t_L g8517 ( 
.A(n_8224),
.Y(n_8517)
);

CKINVDCx16_ASAP7_75t_R g8518 ( 
.A(n_8346),
.Y(n_8518)
);

INVx2_ASAP7_75t_L g8519 ( 
.A(n_8286),
.Y(n_8519)
);

INVx1_ASAP7_75t_L g8520 ( 
.A(n_8273),
.Y(n_8520)
);

AND2x2_ASAP7_75t_L g8521 ( 
.A(n_8218),
.B(n_8282),
.Y(n_8521)
);

OR2x2_ASAP7_75t_L g8522 ( 
.A(n_8231),
.B(n_8101),
.Y(n_8522)
);

BUFx2_ASAP7_75t_L g8523 ( 
.A(n_8258),
.Y(n_8523)
);

AND2x2_ASAP7_75t_L g8524 ( 
.A(n_8216),
.B(n_8168),
.Y(n_8524)
);

INVx2_ASAP7_75t_L g8525 ( 
.A(n_8286),
.Y(n_8525)
);

AND2x2_ASAP7_75t_L g8526 ( 
.A(n_8219),
.B(n_8200),
.Y(n_8526)
);

INVx1_ASAP7_75t_L g8527 ( 
.A(n_8263),
.Y(n_8527)
);

AND2x2_ASAP7_75t_L g8528 ( 
.A(n_8228),
.B(n_8018),
.Y(n_8528)
);

INVx2_ASAP7_75t_L g8529 ( 
.A(n_8307),
.Y(n_8529)
);

INVx1_ASAP7_75t_L g8530 ( 
.A(n_8292),
.Y(n_8530)
);

AOI21xp33_ASAP7_75t_L g8531 ( 
.A1(n_8270),
.A2(n_8112),
.B(n_8111),
.Y(n_8531)
);

AND2x2_ASAP7_75t_L g8532 ( 
.A(n_8229),
.B(n_8071),
.Y(n_8532)
);

INVx2_ASAP7_75t_L g8533 ( 
.A(n_8307),
.Y(n_8533)
);

INVx1_ASAP7_75t_L g8534 ( 
.A(n_8306),
.Y(n_8534)
);

NAND2xp5_ASAP7_75t_L g8535 ( 
.A(n_8236),
.B(n_8154),
.Y(n_8535)
);

AND2x2_ASAP7_75t_L g8536 ( 
.A(n_8237),
.B(n_8344),
.Y(n_8536)
);

INVx2_ASAP7_75t_L g8537 ( 
.A(n_8293),
.Y(n_8537)
);

OR2x2_ASAP7_75t_L g8538 ( 
.A(n_8463),
.B(n_8179),
.Y(n_8538)
);

AOI22xp5_ASAP7_75t_L g8539 ( 
.A1(n_8317),
.A2(n_8100),
.B1(n_8156),
.B2(n_8063),
.Y(n_8539)
);

BUFx3_ASAP7_75t_L g8540 ( 
.A(n_8221),
.Y(n_8540)
);

AOI221xp5_ASAP7_75t_L g8541 ( 
.A1(n_8296),
.A2(n_8128),
.B1(n_8170),
.B2(n_8160),
.C(n_8183),
.Y(n_8541)
);

OR2x2_ASAP7_75t_L g8542 ( 
.A(n_8470),
.B(n_8276),
.Y(n_8542)
);

AND2x2_ASAP7_75t_L g8543 ( 
.A(n_8226),
.B(n_8185),
.Y(n_8543)
);

AND2x2_ASAP7_75t_L g8544 ( 
.A(n_8423),
.B(n_8186),
.Y(n_8544)
);

AOI221xp5_ASAP7_75t_L g8545 ( 
.A1(n_8493),
.A2(n_8170),
.B1(n_8160),
.B2(n_8159),
.C(n_8158),
.Y(n_8545)
);

NAND2xp5_ASAP7_75t_L g8546 ( 
.A(n_8246),
.B(n_8117),
.Y(n_8546)
);

NAND2xp5_ASAP7_75t_L g8547 ( 
.A(n_8221),
.B(n_8289),
.Y(n_8547)
);

NAND2xp5_ASAP7_75t_L g8548 ( 
.A(n_8289),
.B(n_8122),
.Y(n_8548)
);

AND2x2_ASAP7_75t_L g8549 ( 
.A(n_8301),
.B(n_8091),
.Y(n_8549)
);

NAND3xp33_ASAP7_75t_L g8550 ( 
.A(n_8256),
.B(n_8188),
.C(n_8091),
.Y(n_8550)
);

NAND2xp5_ASAP7_75t_L g8551 ( 
.A(n_8312),
.B(n_8150),
.Y(n_8551)
);

OR2x2_ASAP7_75t_L g8552 ( 
.A(n_8470),
.B(n_8198),
.Y(n_8552)
);

INVx2_ASAP7_75t_L g8553 ( 
.A(n_8293),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_8361),
.Y(n_8554)
);

NOR3x1_ASAP7_75t_L g8555 ( 
.A(n_8426),
.B(n_8202),
.C(n_8190),
.Y(n_8555)
);

INVx3_ASAP7_75t_R g8556 ( 
.A(n_8287),
.Y(n_8556)
);

INVx1_ASAP7_75t_SL g8557 ( 
.A(n_8414),
.Y(n_8557)
);

NAND2xp5_ASAP7_75t_L g8558 ( 
.A(n_8312),
.B(n_8171),
.Y(n_8558)
);

AND2x2_ASAP7_75t_L g8559 ( 
.A(n_8211),
.B(n_6403),
.Y(n_8559)
);

INVx2_ASAP7_75t_L g8560 ( 
.A(n_8217),
.Y(n_8560)
);

OAI32xp33_ASAP7_75t_L g8561 ( 
.A1(n_8393),
.A2(n_8163),
.A3(n_5461),
.B1(n_5462),
.B2(n_5460),
.Y(n_8561)
);

XNOR2x2_ASAP7_75t_L g8562 ( 
.A(n_8322),
.B(n_8163),
.Y(n_8562)
);

AND2x2_ASAP7_75t_L g8563 ( 
.A(n_8255),
.B(n_6403),
.Y(n_8563)
);

OR2x2_ASAP7_75t_L g8564 ( 
.A(n_8335),
.B(n_6404),
.Y(n_8564)
);

OR2x2_ASAP7_75t_L g8565 ( 
.A(n_8243),
.B(n_6404),
.Y(n_8565)
);

INVx2_ASAP7_75t_L g8566 ( 
.A(n_8244),
.Y(n_8566)
);

INVx2_ASAP7_75t_SL g8567 ( 
.A(n_8414),
.Y(n_8567)
);

NAND2xp5_ASAP7_75t_L g8568 ( 
.A(n_8338),
.B(n_6593),
.Y(n_8568)
);

NAND4xp25_ASAP7_75t_L g8569 ( 
.A(n_8411),
.B(n_3746),
.C(n_3748),
.D(n_4896),
.Y(n_8569)
);

NAND3xp33_ASAP7_75t_L g8570 ( 
.A(n_8506),
.B(n_6414),
.C(n_6412),
.Y(n_8570)
);

AND2x2_ASAP7_75t_L g8571 ( 
.A(n_8285),
.B(n_6412),
.Y(n_8571)
);

INVx1_ASAP7_75t_L g8572 ( 
.A(n_8213),
.Y(n_8572)
);

OAI211xp5_ASAP7_75t_L g8573 ( 
.A1(n_8227),
.A2(n_4925),
.B(n_4927),
.C(n_6549),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_8213),
.Y(n_8574)
);

BUFx3_ASAP7_75t_L g8575 ( 
.A(n_8225),
.Y(n_8575)
);

AND2x2_ASAP7_75t_L g8576 ( 
.A(n_8302),
.B(n_6414),
.Y(n_8576)
);

INVxp67_ASAP7_75t_SL g8577 ( 
.A(n_8230),
.Y(n_8577)
);

INVxp67_ASAP7_75t_SL g8578 ( 
.A(n_8305),
.Y(n_8578)
);

INVx1_ASAP7_75t_L g8579 ( 
.A(n_8284),
.Y(n_8579)
);

INVx1_ASAP7_75t_L g8580 ( 
.A(n_8284),
.Y(n_8580)
);

NAND2xp5_ASAP7_75t_L g8581 ( 
.A(n_8338),
.B(n_6525),
.Y(n_8581)
);

INVx1_ASAP7_75t_L g8582 ( 
.A(n_8359),
.Y(n_8582)
);

OR2x6_ASAP7_75t_L g8583 ( 
.A(n_8319),
.B(n_3746),
.Y(n_8583)
);

NOR2xp33_ASAP7_75t_L g8584 ( 
.A(n_8288),
.B(n_4900),
.Y(n_8584)
);

AND2x2_ASAP7_75t_L g8585 ( 
.A(n_8428),
.B(n_6423),
.Y(n_8585)
);

OR2x2_ASAP7_75t_L g8586 ( 
.A(n_8428),
.B(n_6432),
.Y(n_8586)
);

INVx1_ASAP7_75t_L g8587 ( 
.A(n_8359),
.Y(n_8587)
);

NAND2xp5_ASAP7_75t_L g8588 ( 
.A(n_8248),
.B(n_8279),
.Y(n_8588)
);

OAI21xp33_ASAP7_75t_L g8589 ( 
.A1(n_8454),
.A2(n_6424),
.B(n_6423),
.Y(n_8589)
);

NAND2xp5_ASAP7_75t_L g8590 ( 
.A(n_8308),
.B(n_6529),
.Y(n_8590)
);

AND2x2_ASAP7_75t_L g8591 ( 
.A(n_8437),
.B(n_6424),
.Y(n_8591)
);

AND2x2_ASAP7_75t_L g8592 ( 
.A(n_8345),
.B(n_6432),
.Y(n_8592)
);

AND2x2_ASAP7_75t_L g8593 ( 
.A(n_8345),
.B(n_6441),
.Y(n_8593)
);

AND2x2_ASAP7_75t_L g8594 ( 
.A(n_8240),
.B(n_6441),
.Y(n_8594)
);

OR2x2_ASAP7_75t_L g8595 ( 
.A(n_8266),
.B(n_6451),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_8275),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_8360),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_8360),
.Y(n_8598)
);

NAND2xp5_ASAP7_75t_L g8599 ( 
.A(n_8448),
.B(n_8244),
.Y(n_8599)
);

NAND2x1_ASAP7_75t_SL g8600 ( 
.A(n_8501),
.B(n_6451),
.Y(n_8600)
);

INVx2_ASAP7_75t_L g8601 ( 
.A(n_8501),
.Y(n_8601)
);

NAND2xp5_ASAP7_75t_L g8602 ( 
.A(n_8242),
.B(n_8245),
.Y(n_8602)
);

NOR2xp33_ASAP7_75t_L g8603 ( 
.A(n_8453),
.B(n_4900),
.Y(n_8603)
);

NAND2x1p5_ASAP7_75t_L g8604 ( 
.A(n_8413),
.B(n_3748),
.Y(n_8604)
);

AND2x2_ASAP7_75t_L g8605 ( 
.A(n_8383),
.B(n_6442),
.Y(n_8605)
);

NAND2xp5_ASAP7_75t_L g8606 ( 
.A(n_8399),
.B(n_8401),
.Y(n_8606)
);

INVx2_ASAP7_75t_L g8607 ( 
.A(n_8503),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_8223),
.Y(n_8608)
);

NAND2x1p5_ASAP7_75t_L g8609 ( 
.A(n_8413),
.B(n_4978),
.Y(n_8609)
);

INVx1_ASAP7_75t_L g8610 ( 
.A(n_8232),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_8234),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_8235),
.Y(n_8612)
);

AND2x2_ASAP7_75t_L g8613 ( 
.A(n_8471),
.B(n_6442),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_8277),
.Y(n_8614)
);

AND2x2_ASAP7_75t_L g8615 ( 
.A(n_8304),
.B(n_6453),
.Y(n_8615)
);

NAND2xp5_ASAP7_75t_L g8616 ( 
.A(n_8328),
.B(n_6567),
.Y(n_8616)
);

NAND2xp5_ASAP7_75t_L g8617 ( 
.A(n_8247),
.B(n_8300),
.Y(n_8617)
);

INVx2_ASAP7_75t_L g8618 ( 
.A(n_8503),
.Y(n_8618)
);

INVx1_ASAP7_75t_L g8619 ( 
.A(n_8253),
.Y(n_8619)
);

INVx1_ASAP7_75t_L g8620 ( 
.A(n_8370),
.Y(n_8620)
);

INVx1_ASAP7_75t_L g8621 ( 
.A(n_8459),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_8274),
.Y(n_8622)
);

NAND2xp5_ASAP7_75t_L g8623 ( 
.A(n_8222),
.B(n_8403),
.Y(n_8623)
);

NAND2xp5_ASAP7_75t_L g8624 ( 
.A(n_8257),
.B(n_6567),
.Y(n_8624)
);

INVx1_ASAP7_75t_L g8625 ( 
.A(n_8241),
.Y(n_8625)
);

OR2x2_ASAP7_75t_L g8626 ( 
.A(n_8357),
.B(n_8406),
.Y(n_8626)
);

OR2x2_ASAP7_75t_L g8627 ( 
.A(n_8259),
.B(n_6469),
.Y(n_8627)
);

INVx1_ASAP7_75t_SL g8628 ( 
.A(n_8265),
.Y(n_8628)
);

AND2x2_ASAP7_75t_L g8629 ( 
.A(n_8436),
.B(n_6453),
.Y(n_8629)
);

INVx1_ASAP7_75t_SL g8630 ( 
.A(n_8268),
.Y(n_8630)
);

NOR2xp67_ASAP7_75t_L g8631 ( 
.A(n_8488),
.B(n_6459),
.Y(n_8631)
);

INVx2_ASAP7_75t_L g8632 ( 
.A(n_8404),
.Y(n_8632)
);

INVx1_ASAP7_75t_L g8633 ( 
.A(n_8262),
.Y(n_8633)
);

INVx2_ASAP7_75t_L g8634 ( 
.A(n_8404),
.Y(n_8634)
);

AND2x2_ASAP7_75t_L g8635 ( 
.A(n_8415),
.B(n_6459),
.Y(n_8635)
);

AND2x2_ASAP7_75t_L g8636 ( 
.A(n_8415),
.B(n_6469),
.Y(n_8636)
);

INVx1_ASAP7_75t_L g8637 ( 
.A(n_8251),
.Y(n_8637)
);

INVx1_ASAP7_75t_L g8638 ( 
.A(n_8252),
.Y(n_8638)
);

HB1xp67_ASAP7_75t_L g8639 ( 
.A(n_8298),
.Y(n_8639)
);

AND2x2_ASAP7_75t_L g8640 ( 
.A(n_8417),
.B(n_6471),
.Y(n_8640)
);

BUFx3_ASAP7_75t_L g8641 ( 
.A(n_8481),
.Y(n_8641)
);

INVx3_ASAP7_75t_L g8642 ( 
.A(n_8299),
.Y(n_8642)
);

AND2x2_ASAP7_75t_L g8643 ( 
.A(n_8442),
.B(n_6471),
.Y(n_8643)
);

INVxp67_ASAP7_75t_SL g8644 ( 
.A(n_8395),
.Y(n_8644)
);

INVx1_ASAP7_75t_L g8645 ( 
.A(n_8407),
.Y(n_8645)
);

INVxp67_ASAP7_75t_L g8646 ( 
.A(n_8330),
.Y(n_8646)
);

AND2x2_ASAP7_75t_L g8647 ( 
.A(n_8445),
.B(n_6472),
.Y(n_8647)
);

NAND2x1_ASAP7_75t_L g8648 ( 
.A(n_8352),
.B(n_6472),
.Y(n_8648)
);

INVx1_ASAP7_75t_L g8649 ( 
.A(n_8407),
.Y(n_8649)
);

INVx2_ASAP7_75t_L g8650 ( 
.A(n_8381),
.Y(n_8650)
);

INVx2_ASAP7_75t_L g8651 ( 
.A(n_8381),
.Y(n_8651)
);

NAND2xp5_ASAP7_75t_L g8652 ( 
.A(n_8280),
.B(n_6615),
.Y(n_8652)
);

INVx1_ASAP7_75t_L g8653 ( 
.A(n_8424),
.Y(n_8653)
);

BUFx2_ASAP7_75t_L g8654 ( 
.A(n_8488),
.Y(n_8654)
);

OR2x6_ASAP7_75t_L g8655 ( 
.A(n_8382),
.B(n_4900),
.Y(n_8655)
);

INVx1_ASAP7_75t_L g8656 ( 
.A(n_8424),
.Y(n_8656)
);

INVx1_ASAP7_75t_L g8657 ( 
.A(n_8505),
.Y(n_8657)
);

INVx1_ASAP7_75t_L g8658 ( 
.A(n_8297),
.Y(n_8658)
);

INVx2_ASAP7_75t_SL g8659 ( 
.A(n_8299),
.Y(n_8659)
);

AND2x2_ASAP7_75t_L g8660 ( 
.A(n_8453),
.B(n_6478),
.Y(n_8660)
);

NOR2x1_ASAP7_75t_L g8661 ( 
.A(n_8409),
.B(n_6478),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_8283),
.Y(n_8662)
);

INVx1_ASAP7_75t_L g8663 ( 
.A(n_8249),
.Y(n_8663)
);

INVx2_ASAP7_75t_SL g8664 ( 
.A(n_8427),
.Y(n_8664)
);

NAND2xp5_ASAP7_75t_L g8665 ( 
.A(n_8278),
.B(n_6486),
.Y(n_8665)
);

NAND2xp5_ASAP7_75t_L g8666 ( 
.A(n_8303),
.B(n_6486),
.Y(n_8666)
);

AND2x2_ASAP7_75t_L g8667 ( 
.A(n_8453),
.B(n_6489),
.Y(n_8667)
);

BUFx2_ASAP7_75t_L g8668 ( 
.A(n_8311),
.Y(n_8668)
);

NAND2xp5_ASAP7_75t_L g8669 ( 
.A(n_8464),
.B(n_6517),
.Y(n_8669)
);

INVx1_ASAP7_75t_L g8670 ( 
.A(n_8316),
.Y(n_8670)
);

OR2x6_ASAP7_75t_L g8671 ( 
.A(n_8290),
.B(n_4900),
.Y(n_8671)
);

NAND2x1p5_ASAP7_75t_L g8672 ( 
.A(n_8413),
.B(n_4978),
.Y(n_8672)
);

INVx1_ASAP7_75t_L g8673 ( 
.A(n_8318),
.Y(n_8673)
);

AND2x2_ASAP7_75t_L g8674 ( 
.A(n_8457),
.B(n_6489),
.Y(n_8674)
);

NAND2xp5_ASAP7_75t_L g8675 ( 
.A(n_8464),
.B(n_6528),
.Y(n_8675)
);

AOI22xp5_ASAP7_75t_L g8676 ( 
.A1(n_8353),
.A2(n_5036),
.B1(n_5095),
.B2(n_4899),
.Y(n_8676)
);

NAND2xp5_ASAP7_75t_L g8677 ( 
.A(n_8309),
.B(n_6528),
.Y(n_8677)
);

AND2x2_ASAP7_75t_L g8678 ( 
.A(n_8354),
.B(n_6497),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_L g8679 ( 
.A(n_8295),
.B(n_6529),
.Y(n_8679)
);

INVx2_ASAP7_75t_L g8680 ( 
.A(n_8389),
.Y(n_8680)
);

NAND2xp5_ASAP7_75t_L g8681 ( 
.A(n_8314),
.B(n_6535),
.Y(n_8681)
);

BUFx2_ASAP7_75t_L g8682 ( 
.A(n_8389),
.Y(n_8682)
);

INVx2_ASAP7_75t_L g8683 ( 
.A(n_8427),
.Y(n_8683)
);

NAND2xp5_ASAP7_75t_L g8684 ( 
.A(n_8458),
.B(n_6535),
.Y(n_8684)
);

INVx1_ASAP7_75t_L g8685 ( 
.A(n_8409),
.Y(n_8685)
);

XNOR2x1_ASAP7_75t_L g8686 ( 
.A(n_8353),
.B(n_4896),
.Y(n_8686)
);

INVxp67_ASAP7_75t_SL g8687 ( 
.A(n_8323),
.Y(n_8687)
);

OAI21xp33_ASAP7_75t_L g8688 ( 
.A1(n_8495),
.A2(n_6500),
.B(n_6497),
.Y(n_8688)
);

INVxp67_ASAP7_75t_SL g8689 ( 
.A(n_8291),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8492),
.Y(n_8690)
);

NAND3xp33_ASAP7_75t_L g8691 ( 
.A(n_8220),
.B(n_6504),
.C(n_6500),
.Y(n_8691)
);

AND2x2_ASAP7_75t_L g8692 ( 
.A(n_8355),
.B(n_6504),
.Y(n_8692)
);

NAND2xp5_ASAP7_75t_SL g8693 ( 
.A(n_8486),
.B(n_4899),
.Y(n_8693)
);

AND2x2_ASAP7_75t_L g8694 ( 
.A(n_8485),
.B(n_8487),
.Y(n_8694)
);

INVx1_ASAP7_75t_L g8695 ( 
.A(n_8294),
.Y(n_8695)
);

AND2x2_ASAP7_75t_L g8696 ( 
.A(n_8377),
.B(n_6506),
.Y(n_8696)
);

INVxp67_ASAP7_75t_L g8697 ( 
.A(n_8477),
.Y(n_8697)
);

NAND2xp5_ASAP7_75t_L g8698 ( 
.A(n_8458),
.B(n_6585),
.Y(n_8698)
);

HB1xp67_ASAP7_75t_L g8699 ( 
.A(n_8433),
.Y(n_8699)
);

NAND2xp5_ASAP7_75t_L g8700 ( 
.A(n_8239),
.B(n_6593),
.Y(n_8700)
);

NAND3xp33_ASAP7_75t_L g8701 ( 
.A(n_8254),
.B(n_6507),
.C(n_6506),
.Y(n_8701)
);

INVx1_ASAP7_75t_L g8702 ( 
.A(n_8390),
.Y(n_8702)
);

OR2x2_ASAP7_75t_L g8703 ( 
.A(n_8378),
.B(n_6516),
.Y(n_8703)
);

INVx1_ASAP7_75t_L g8704 ( 
.A(n_8412),
.Y(n_8704)
);

INVx1_ASAP7_75t_L g8705 ( 
.A(n_8491),
.Y(n_8705)
);

NAND2xp5_ASAP7_75t_SL g8706 ( 
.A(n_8486),
.B(n_4899),
.Y(n_8706)
);

INVx2_ASAP7_75t_L g8707 ( 
.A(n_8339),
.Y(n_8707)
);

OR2x2_ASAP7_75t_L g8708 ( 
.A(n_8455),
.B(n_6516),
.Y(n_8708)
);

INVxp67_ASAP7_75t_L g8709 ( 
.A(n_8269),
.Y(n_8709)
);

INVxp67_ASAP7_75t_L g8710 ( 
.A(n_8233),
.Y(n_8710)
);

NAND2x2_ASAP7_75t_L g8711 ( 
.A(n_8367),
.B(n_4976),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8443),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_8387),
.Y(n_8713)
);

INVx1_ASAP7_75t_L g8714 ( 
.A(n_8372),
.Y(n_8714)
);

AOI22xp5_ASAP7_75t_L g8715 ( 
.A1(n_8465),
.A2(n_4899),
.B1(n_5095),
.B2(n_5036),
.Y(n_8715)
);

AND2x2_ASAP7_75t_L g8716 ( 
.A(n_8341),
.B(n_6507),
.Y(n_8716)
);

INVx1_ASAP7_75t_L g8717 ( 
.A(n_8396),
.Y(n_8717)
);

AND2x2_ASAP7_75t_L g8718 ( 
.A(n_8363),
.B(n_6517),
.Y(n_8718)
);

INVx1_ASAP7_75t_L g8719 ( 
.A(n_8342),
.Y(n_8719)
);

OR2x2_ASAP7_75t_L g8720 ( 
.A(n_8475),
.B(n_6554),
.Y(n_8720)
);

OR2x2_ASAP7_75t_L g8721 ( 
.A(n_8397),
.B(n_6554),
.Y(n_8721)
);

INVx3_ASAP7_75t_L g8722 ( 
.A(n_8325),
.Y(n_8722)
);

AND2x2_ASAP7_75t_L g8723 ( 
.A(n_8356),
.B(n_6525),
.Y(n_8723)
);

NAND2xp5_ASAP7_75t_L g8724 ( 
.A(n_8215),
.B(n_6557),
.Y(n_8724)
);

INVx1_ASAP7_75t_L g8725 ( 
.A(n_8358),
.Y(n_8725)
);

HB1xp67_ASAP7_75t_L g8726 ( 
.A(n_8267),
.Y(n_8726)
);

OR2x2_ASAP7_75t_L g8727 ( 
.A(n_8497),
.B(n_6563),
.Y(n_8727)
);

NAND2xp5_ASAP7_75t_L g8728 ( 
.A(n_8238),
.B(n_6557),
.Y(n_8728)
);

BUFx3_ASAP7_75t_L g8729 ( 
.A(n_8451),
.Y(n_8729)
);

INVx1_ASAP7_75t_L g8730 ( 
.A(n_8467),
.Y(n_8730)
);

INVx1_ASAP7_75t_L g8731 ( 
.A(n_8474),
.Y(n_8731)
);

HB1xp67_ASAP7_75t_L g8732 ( 
.A(n_8466),
.Y(n_8732)
);

OR2x2_ASAP7_75t_L g8733 ( 
.A(n_8365),
.B(n_6565),
.Y(n_8733)
);

INVx2_ASAP7_75t_L g8734 ( 
.A(n_8325),
.Y(n_8734)
);

INVx1_ASAP7_75t_L g8735 ( 
.A(n_8449),
.Y(n_8735)
);

OR2x2_ASAP7_75t_L g8736 ( 
.A(n_8496),
.B(n_6565),
.Y(n_8736)
);

NAND2xp5_ASAP7_75t_L g8737 ( 
.A(n_8364),
.B(n_8260),
.Y(n_8737)
);

INVx1_ASAP7_75t_L g8738 ( 
.A(n_8435),
.Y(n_8738)
);

AOI221xp5_ASAP7_75t_L g8739 ( 
.A1(n_8264),
.A2(n_6256),
.B1(n_6247),
.B2(n_6235),
.C(n_6563),
.Y(n_8739)
);

OR2x2_ASAP7_75t_L g8740 ( 
.A(n_8431),
.B(n_8444),
.Y(n_8740)
);

INVx1_ASAP7_75t_SL g8741 ( 
.A(n_8466),
.Y(n_8741)
);

AND2x2_ASAP7_75t_L g8742 ( 
.A(n_8337),
.B(n_6610),
.Y(n_8742)
);

BUFx3_ASAP7_75t_L g8743 ( 
.A(n_8490),
.Y(n_8743)
);

NAND2xp5_ASAP7_75t_L g8744 ( 
.A(n_8364),
.B(n_8214),
.Y(n_8744)
);

NAND2xp5_ASAP7_75t_L g8745 ( 
.A(n_8343),
.B(n_6610),
.Y(n_8745)
);

NAND2xp5_ASAP7_75t_L g8746 ( 
.A(n_8326),
.B(n_6613),
.Y(n_8746)
);

NAND2xp5_ASAP7_75t_L g8747 ( 
.A(n_8326),
.B(n_6613),
.Y(n_8747)
);

NOR2xp33_ASAP7_75t_L g8748 ( 
.A(n_8447),
.B(n_6615),
.Y(n_8748)
);

INVx1_ASAP7_75t_L g8749 ( 
.A(n_8394),
.Y(n_8749)
);

INVx2_ASAP7_75t_L g8750 ( 
.A(n_8329),
.Y(n_8750)
);

INVx1_ASAP7_75t_L g8751 ( 
.A(n_8482),
.Y(n_8751)
);

HB1xp67_ASAP7_75t_L g8752 ( 
.A(n_8334),
.Y(n_8752)
);

NAND2xp5_ASAP7_75t_L g8753 ( 
.A(n_8439),
.B(n_6015),
.Y(n_8753)
);

NAND2xp5_ASAP7_75t_L g8754 ( 
.A(n_8460),
.B(n_6030),
.Y(n_8754)
);

NAND2xp5_ASAP7_75t_L g8755 ( 
.A(n_8369),
.B(n_6032),
.Y(n_8755)
);

INVx1_ASAP7_75t_SL g8756 ( 
.A(n_8337),
.Y(n_8756)
);

NAND2xp5_ASAP7_75t_L g8757 ( 
.A(n_8440),
.B(n_6045),
.Y(n_8757)
);

INVx2_ASAP7_75t_L g8758 ( 
.A(n_8349),
.Y(n_8758)
);

OR2x2_ASAP7_75t_L g8759 ( 
.A(n_8446),
.B(n_6316),
.Y(n_8759)
);

NAND2xp5_ASAP7_75t_L g8760 ( 
.A(n_8479),
.B(n_5655),
.Y(n_8760)
);

AND3x2_ASAP7_75t_L g8761 ( 
.A(n_8315),
.B(n_4763),
.C(n_4686),
.Y(n_8761)
);

INVx1_ASAP7_75t_L g8762 ( 
.A(n_8320),
.Y(n_8762)
);

NOR2xp33_ASAP7_75t_SL g8763 ( 
.A(n_8313),
.B(n_4899),
.Y(n_8763)
);

AND2x2_ASAP7_75t_L g8764 ( 
.A(n_8476),
.B(n_4849),
.Y(n_8764)
);

INVx1_ASAP7_75t_L g8765 ( 
.A(n_8321),
.Y(n_8765)
);

INVx1_ASAP7_75t_L g8766 ( 
.A(n_8324),
.Y(n_8766)
);

INVxp67_ASAP7_75t_L g8767 ( 
.A(n_8654),
.Y(n_8767)
);

AO21x1_ASAP7_75t_L g8768 ( 
.A1(n_8578),
.A2(n_8658),
.B(n_8552),
.Y(n_8768)
);

XOR2x2_ASAP7_75t_L g8769 ( 
.A(n_8521),
.B(n_8281),
.Y(n_8769)
);

AND2x2_ASAP7_75t_L g8770 ( 
.A(n_8536),
.B(n_8473),
.Y(n_8770)
);

OA21x2_ASAP7_75t_L g8771 ( 
.A1(n_8658),
.A2(n_8441),
.B(n_8375),
.Y(n_8771)
);

INVx1_ASAP7_75t_L g8772 ( 
.A(n_8562),
.Y(n_8772)
);

INVx1_ASAP7_75t_L g8773 ( 
.A(n_8512),
.Y(n_8773)
);

OAI22xp33_ASAP7_75t_L g8774 ( 
.A1(n_8516),
.A2(n_8504),
.B1(n_8310),
.B2(n_8385),
.Y(n_8774)
);

INVx1_ASAP7_75t_L g8775 ( 
.A(n_8682),
.Y(n_8775)
);

INVx1_ASAP7_75t_L g8776 ( 
.A(n_8732),
.Y(n_8776)
);

NAND2xp5_ASAP7_75t_L g8777 ( 
.A(n_8540),
.B(n_8333),
.Y(n_8777)
);

INVx1_ASAP7_75t_L g8778 ( 
.A(n_8513),
.Y(n_8778)
);

O2A1O1Ixp33_ASAP7_75t_L g8779 ( 
.A1(n_8515),
.A2(n_8212),
.B(n_8461),
.C(n_8340),
.Y(n_8779)
);

INVx1_ASAP7_75t_L g8780 ( 
.A(n_8542),
.Y(n_8780)
);

AOI22xp5_ASAP7_75t_L g8781 ( 
.A1(n_8518),
.A2(n_8376),
.B1(n_8416),
.B2(n_8429),
.Y(n_8781)
);

NOR2xp33_ASAP7_75t_L g8782 ( 
.A(n_8557),
.B(n_8408),
.Y(n_8782)
);

AND2x4_ASAP7_75t_L g8783 ( 
.A(n_8567),
.B(n_8336),
.Y(n_8783)
);

INVx1_ASAP7_75t_SL g8784 ( 
.A(n_8547),
.Y(n_8784)
);

NAND3xp33_ASAP7_75t_L g8785 ( 
.A(n_8541),
.B(n_8332),
.C(n_8405),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_8668),
.Y(n_8786)
);

INVx2_ASAP7_75t_SL g8787 ( 
.A(n_8600),
.Y(n_8787)
);

INVx1_ASAP7_75t_L g8788 ( 
.A(n_8601),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_8607),
.Y(n_8789)
);

AOI32xp33_ASAP7_75t_L g8790 ( 
.A1(n_8545),
.A2(n_8392),
.A3(n_8500),
.B1(n_8425),
.B2(n_8499),
.Y(n_8790)
);

INVx2_ASAP7_75t_SL g8791 ( 
.A(n_8641),
.Y(n_8791)
);

OAI22xp33_ASAP7_75t_L g8792 ( 
.A1(n_8577),
.A2(n_8371),
.B1(n_8483),
.B2(n_8478),
.Y(n_8792)
);

NOR2xp33_ASAP7_75t_SL g8793 ( 
.A(n_8528),
.B(n_8366),
.Y(n_8793)
);

AND2x2_ASAP7_75t_L g8794 ( 
.A(n_8532),
.B(n_8386),
.Y(n_8794)
);

AND2x2_ASAP7_75t_L g8795 ( 
.A(n_8575),
.B(n_8410),
.Y(n_8795)
);

OAI22xp5_ASAP7_75t_L g8796 ( 
.A1(n_8697),
.A2(n_8484),
.B1(n_8509),
.B2(n_8502),
.Y(n_8796)
);

INVx1_ASAP7_75t_L g8797 ( 
.A(n_8618),
.Y(n_8797)
);

AOI22xp5_ASAP7_75t_L g8798 ( 
.A1(n_8573),
.A2(n_8603),
.B1(n_8763),
.B2(n_8584),
.Y(n_8798)
);

INVx2_ASAP7_75t_L g8799 ( 
.A(n_8511),
.Y(n_8799)
);

INVx1_ASAP7_75t_L g8800 ( 
.A(n_8579),
.Y(n_8800)
);

INVx1_ASAP7_75t_L g8801 ( 
.A(n_8580),
.Y(n_8801)
);

AND2x2_ASAP7_75t_L g8802 ( 
.A(n_8694),
.B(n_8430),
.Y(n_8802)
);

OAI21xp5_ASAP7_75t_L g8803 ( 
.A1(n_8550),
.A2(n_8480),
.B(n_8450),
.Y(n_8803)
);

AOI22xp5_ASAP7_75t_L g8804 ( 
.A1(n_8630),
.A2(n_8327),
.B1(n_8452),
.B2(n_8489),
.Y(n_8804)
);

OAI21xp5_ASAP7_75t_L g8805 ( 
.A1(n_8709),
.A2(n_8468),
.B(n_8456),
.Y(n_8805)
);

OAI22xp33_ASAP7_75t_L g8806 ( 
.A1(n_8728),
.A2(n_8432),
.B1(n_8351),
.B2(n_8362),
.Y(n_8806)
);

INVx1_ASAP7_75t_L g8807 ( 
.A(n_8582),
.Y(n_8807)
);

INVx2_ASAP7_75t_L g8808 ( 
.A(n_8511),
.Y(n_8808)
);

INVx1_ASAP7_75t_SL g8809 ( 
.A(n_8628),
.Y(n_8809)
);

AND2x2_ASAP7_75t_L g8810 ( 
.A(n_8543),
.B(n_8632),
.Y(n_8810)
);

NAND4xp75_ASAP7_75t_L g8811 ( 
.A(n_8555),
.B(n_8348),
.C(n_8402),
.D(n_8388),
.Y(n_8811)
);

INVx1_ASAP7_75t_L g8812 ( 
.A(n_8587),
.Y(n_8812)
);

AOI21xp5_ASAP7_75t_L g8813 ( 
.A1(n_8687),
.A2(n_8739),
.B(n_8648),
.Y(n_8813)
);

AND2x4_ASAP7_75t_L g8814 ( 
.A(n_8664),
.B(n_8418),
.Y(n_8814)
);

NAND2xp5_ASAP7_75t_L g8815 ( 
.A(n_8639),
.B(n_8419),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_8519),
.Y(n_8816)
);

INVxp67_ASAP7_75t_SL g8817 ( 
.A(n_8604),
.Y(n_8817)
);

INVx2_ASAP7_75t_L g8818 ( 
.A(n_8722),
.Y(n_8818)
);

AND2x2_ASAP7_75t_L g8819 ( 
.A(n_8634),
.B(n_8347),
.Y(n_8819)
);

NAND2xp5_ASAP7_75t_L g8820 ( 
.A(n_8670),
.B(n_8420),
.Y(n_8820)
);

OAI22xp5_ASAP7_75t_L g8821 ( 
.A1(n_8539),
.A2(n_8510),
.B1(n_8384),
.B2(n_8398),
.Y(n_8821)
);

OR2x2_ASAP7_75t_L g8822 ( 
.A(n_8529),
.B(n_8421),
.Y(n_8822)
);

A2O1A1Ixp33_ASAP7_75t_L g8823 ( 
.A1(n_8705),
.A2(n_8331),
.B(n_8494),
.C(n_8400),
.Y(n_8823)
);

NAND2xp5_ASAP7_75t_L g8824 ( 
.A(n_8673),
.B(n_8391),
.Y(n_8824)
);

CKINVDCx16_ASAP7_75t_R g8825 ( 
.A(n_8743),
.Y(n_8825)
);

NAND2xp5_ASAP7_75t_L g8826 ( 
.A(n_8533),
.B(n_8537),
.Y(n_8826)
);

INVx1_ASAP7_75t_L g8827 ( 
.A(n_8525),
.Y(n_8827)
);

AOI32xp33_ASAP7_75t_L g8828 ( 
.A1(n_8523),
.A2(n_8373),
.A3(n_8438),
.B1(n_8469),
.B2(n_8462),
.Y(n_8828)
);

OAI22xp33_ASAP7_75t_R g8829 ( 
.A1(n_8741),
.A2(n_8368),
.B1(n_8434),
.B2(n_8507),
.Y(n_8829)
);

AND2x4_ASAP7_75t_L g8830 ( 
.A(n_8722),
.B(n_8380),
.Y(n_8830)
);

AND2x2_ASAP7_75t_L g8831 ( 
.A(n_8752),
.B(n_8350),
.Y(n_8831)
);

INVx1_ASAP7_75t_L g8832 ( 
.A(n_8617),
.Y(n_8832)
);

INVx1_ASAP7_75t_L g8833 ( 
.A(n_8553),
.Y(n_8833)
);

INVx1_ASAP7_75t_L g8834 ( 
.A(n_8517),
.Y(n_8834)
);

INVx1_ASAP7_75t_L g8835 ( 
.A(n_8699),
.Y(n_8835)
);

NOR2xp67_ASAP7_75t_R g8836 ( 
.A(n_8620),
.B(n_8374),
.Y(n_8836)
);

INVx1_ASAP7_75t_L g8837 ( 
.A(n_8661),
.Y(n_8837)
);

INVx1_ASAP7_75t_L g8838 ( 
.A(n_8680),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_8642),
.Y(n_8839)
);

INVx1_ASAP7_75t_L g8840 ( 
.A(n_8599),
.Y(n_8840)
);

A2O1A1Ixp33_ASAP7_75t_L g8841 ( 
.A1(n_8695),
.A2(n_8508),
.B(n_8379),
.C(n_8498),
.Y(n_8841)
);

OAI22xp5_ASAP7_75t_L g8842 ( 
.A1(n_8606),
.A2(n_5416),
.B1(n_5431),
.B2(n_5373),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_8631),
.Y(n_8843)
);

AOI22xp5_ASAP7_75t_L g8844 ( 
.A1(n_8644),
.A2(n_8472),
.B1(n_4899),
.B2(n_5095),
.Y(n_8844)
);

BUFx2_ASAP7_75t_L g8845 ( 
.A(n_8560),
.Y(n_8845)
);

AOI22xp5_ASAP7_75t_L g8846 ( 
.A1(n_8549),
.A2(n_5095),
.B1(n_5148),
.B2(n_5036),
.Y(n_8846)
);

INVx2_ASAP7_75t_L g8847 ( 
.A(n_8642),
.Y(n_8847)
);

NOR3xp33_ASAP7_75t_L g8848 ( 
.A(n_8646),
.B(n_5004),
.C(n_4976),
.Y(n_8848)
);

AOI222xp33_ASAP7_75t_L g8849 ( 
.A1(n_8695),
.A2(n_5461),
.B1(n_5458),
.B2(n_5463),
.C1(n_5462),
.C2(n_5460),
.Y(n_8849)
);

INVx2_ASAP7_75t_L g8850 ( 
.A(n_8566),
.Y(n_8850)
);

INVx1_ASAP7_75t_L g8851 ( 
.A(n_8538),
.Y(n_8851)
);

AOI32xp33_ASAP7_75t_L g8852 ( 
.A1(n_8686),
.A2(n_5354),
.A3(n_5314),
.B1(n_5307),
.B2(n_5416),
.Y(n_8852)
);

INVx1_ASAP7_75t_L g8853 ( 
.A(n_8512),
.Y(n_8853)
);

OAI22xp5_ASAP7_75t_L g8854 ( 
.A1(n_8676),
.A2(n_5416),
.B1(n_5431),
.B2(n_5373),
.Y(n_8854)
);

AND2x2_ASAP7_75t_L g8855 ( 
.A(n_8576),
.B(n_4849),
.Y(n_8855)
);

HB1xp67_ASAP7_75t_L g8856 ( 
.A(n_8556),
.Y(n_8856)
);

OR2x2_ASAP7_75t_L g8857 ( 
.A(n_8602),
.B(n_6509),
.Y(n_8857)
);

AND2x2_ASAP7_75t_L g8858 ( 
.A(n_8544),
.B(n_4761),
.Y(n_8858)
);

OAI21xp33_ASAP7_75t_L g8859 ( 
.A1(n_8569),
.A2(n_5043),
.B(n_5004),
.Y(n_8859)
);

INVx2_ASAP7_75t_L g8860 ( 
.A(n_8683),
.Y(n_8860)
);

INVx2_ASAP7_75t_L g8861 ( 
.A(n_8609),
.Y(n_8861)
);

INVx2_ASAP7_75t_L g8862 ( 
.A(n_8672),
.Y(n_8862)
);

NAND2xp5_ASAP7_75t_L g8863 ( 
.A(n_8756),
.B(n_5657),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_8548),
.Y(n_8864)
);

INVx1_ASAP7_75t_L g8865 ( 
.A(n_8614),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_8619),
.Y(n_8866)
);

INVx2_ASAP7_75t_L g8867 ( 
.A(n_8734),
.Y(n_8867)
);

OAI32xp33_ASAP7_75t_L g8868 ( 
.A1(n_8551),
.A2(n_5463),
.A3(n_5461),
.B1(n_5462),
.B2(n_5460),
.Y(n_8868)
);

INVxp67_ASAP7_75t_SL g8869 ( 
.A(n_8621),
.Y(n_8869)
);

NAND2xp5_ASAP7_75t_L g8870 ( 
.A(n_8659),
.B(n_5657),
.Y(n_8870)
);

NAND2xp5_ASAP7_75t_L g8871 ( 
.A(n_8650),
.B(n_5659),
.Y(n_8871)
);

INVx1_ASAP7_75t_L g8872 ( 
.A(n_8588),
.Y(n_8872)
);

INVx1_ASAP7_75t_L g8873 ( 
.A(n_8626),
.Y(n_8873)
);

HB1xp67_ASAP7_75t_L g8874 ( 
.A(n_8685),
.Y(n_8874)
);

NAND2xp5_ASAP7_75t_L g8875 ( 
.A(n_8651),
.B(n_5659),
.Y(n_8875)
);

AND2x2_ASAP7_75t_SL g8876 ( 
.A(n_8660),
.B(n_4978),
.Y(n_8876)
);

AND2x2_ASAP7_75t_L g8877 ( 
.A(n_8750),
.B(n_8707),
.Y(n_8877)
);

AOI321xp33_ASAP7_75t_L g8878 ( 
.A1(n_8623),
.A2(n_4626),
.A3(n_4358),
.B1(n_4342),
.B2(n_4386),
.C(n_4370),
.Y(n_8878)
);

OR2x2_ASAP7_75t_L g8879 ( 
.A(n_8546),
.B(n_6509),
.Y(n_8879)
);

NAND2xp5_ASAP7_75t_L g8880 ( 
.A(n_8667),
.B(n_5665),
.Y(n_8880)
);

OR2x2_ASAP7_75t_L g8881 ( 
.A(n_8758),
.B(n_6509),
.Y(n_8881)
);

INVx2_ASAP7_75t_L g8882 ( 
.A(n_8583),
.Y(n_8882)
);

HB1xp67_ASAP7_75t_L g8883 ( 
.A(n_8583),
.Y(n_8883)
);

OR2x2_ASAP7_75t_L g8884 ( 
.A(n_8522),
.B(n_6316),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_8514),
.Y(n_8885)
);

NAND2xp5_ASAP7_75t_L g8886 ( 
.A(n_8662),
.B(n_5665),
.Y(n_8886)
);

AND2x4_ASAP7_75t_SL g8887 ( 
.A(n_8655),
.B(n_5036),
.Y(n_8887)
);

AND2x2_ASAP7_75t_L g8888 ( 
.A(n_8524),
.B(n_4761),
.Y(n_8888)
);

INVx1_ASAP7_75t_L g8889 ( 
.A(n_8514),
.Y(n_8889)
);

AO221x1_ASAP7_75t_L g8890 ( 
.A1(n_8710),
.A2(n_5148),
.B1(n_5191),
.B2(n_5095),
.C(n_5036),
.Y(n_8890)
);

AOI22xp5_ASAP7_75t_L g8891 ( 
.A1(n_8737),
.A2(n_8526),
.B1(n_8757),
.B2(n_8613),
.Y(n_8891)
);

NAND2xp5_ASAP7_75t_L g8892 ( 
.A(n_8696),
.B(n_5666),
.Y(n_8892)
);

INVx1_ASAP7_75t_L g8893 ( 
.A(n_8520),
.Y(n_8893)
);

NAND2xp5_ASAP7_75t_L g8894 ( 
.A(n_8712),
.B(n_5666),
.Y(n_8894)
);

OAI22xp5_ASAP7_75t_L g8895 ( 
.A1(n_8711),
.A2(n_8715),
.B1(n_8744),
.B2(n_8625),
.Y(n_8895)
);

INVx2_ASAP7_75t_SL g8896 ( 
.A(n_8655),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8520),
.Y(n_8897)
);

INVx1_ASAP7_75t_L g8898 ( 
.A(n_8527),
.Y(n_8898)
);

NOR2xp67_ASAP7_75t_SL g8899 ( 
.A(n_8638),
.B(n_5095),
.Y(n_8899)
);

NAND2xp5_ASAP7_75t_L g8900 ( 
.A(n_8730),
.B(n_5676),
.Y(n_8900)
);

INVx1_ASAP7_75t_L g8901 ( 
.A(n_8527),
.Y(n_8901)
);

AND2x2_ASAP7_75t_L g8902 ( 
.A(n_8729),
.B(n_4778),
.Y(n_8902)
);

BUFx2_ASAP7_75t_SL g8903 ( 
.A(n_8690),
.Y(n_8903)
);

OAI31xp33_ASAP7_75t_L g8904 ( 
.A1(n_8558),
.A2(n_8531),
.A3(n_8589),
.B(n_8570),
.Y(n_8904)
);

INVx2_ASAP7_75t_L g8905 ( 
.A(n_8586),
.Y(n_8905)
);

AOI32xp33_ASAP7_75t_L g8906 ( 
.A1(n_8663),
.A2(n_5354),
.A3(n_5314),
.B1(n_5307),
.B2(n_5431),
.Y(n_8906)
);

INVx1_ASAP7_75t_L g8907 ( 
.A(n_8657),
.Y(n_8907)
);

OAI22xp5_ASAP7_75t_L g8908 ( 
.A1(n_8535),
.A2(n_5383),
.B1(n_5262),
.B2(n_5336),
.Y(n_8908)
);

OAI22xp5_ASAP7_75t_L g8909 ( 
.A1(n_8637),
.A2(n_5383),
.B1(n_5262),
.B2(n_5336),
.Y(n_8909)
);

AND2x2_ASAP7_75t_L g8910 ( 
.A(n_8571),
.B(n_4778),
.Y(n_8910)
);

INVx2_ASAP7_75t_L g8911 ( 
.A(n_8564),
.Y(n_8911)
);

OAI22xp5_ASAP7_75t_L g8912 ( 
.A1(n_8701),
.A2(n_5383),
.B1(n_5321),
.B2(n_5336),
.Y(n_8912)
);

INVx2_ASAP7_75t_SL g8913 ( 
.A(n_8592),
.Y(n_8913)
);

AND2x2_ASAP7_75t_L g8914 ( 
.A(n_8605),
.B(n_4781),
.Y(n_8914)
);

NAND2xp5_ASAP7_75t_L g8915 ( 
.A(n_8594),
.B(n_5676),
.Y(n_8915)
);

INVx1_ASAP7_75t_L g8916 ( 
.A(n_8657),
.Y(n_8916)
);

AND2x2_ASAP7_75t_L g8917 ( 
.A(n_8671),
.B(n_4781),
.Y(n_8917)
);

OAI32xp33_ASAP7_75t_L g8918 ( 
.A1(n_8554),
.A2(n_5463),
.A3(n_5458),
.B1(n_5901),
.B2(n_5830),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_8530),
.Y(n_8919)
);

NAND2xp5_ASAP7_75t_L g8920 ( 
.A(n_8735),
.B(n_5685),
.Y(n_8920)
);

AOI32xp33_ASAP7_75t_L g8921 ( 
.A1(n_8731),
.A2(n_8534),
.A3(n_8622),
.B1(n_8716),
.B2(n_8718),
.Y(n_8921)
);

INVx1_ASAP7_75t_L g8922 ( 
.A(n_8563),
.Y(n_8922)
);

INVx2_ASAP7_75t_L g8923 ( 
.A(n_8593),
.Y(n_8923)
);

AND2x2_ASAP7_75t_SL g8924 ( 
.A(n_8751),
.B(n_4978),
.Y(n_8924)
);

INVx1_ASAP7_75t_L g8925 ( 
.A(n_8597),
.Y(n_8925)
);

INVx1_ASAP7_75t_L g8926 ( 
.A(n_8597),
.Y(n_8926)
);

AND2x2_ASAP7_75t_L g8927 ( 
.A(n_8671),
.B(n_5235),
.Y(n_8927)
);

INVxp67_ASAP7_75t_L g8928 ( 
.A(n_8693),
.Y(n_8928)
);

BUFx3_ASAP7_75t_L g8929 ( 
.A(n_8713),
.Y(n_8929)
);

OAI32xp33_ASAP7_75t_L g8930 ( 
.A1(n_8700),
.A2(n_5458),
.A3(n_5901),
.B1(n_5909),
.B2(n_5830),
.Y(n_8930)
);

OAI22xp33_ASAP7_75t_L g8931 ( 
.A1(n_8724),
.A2(n_5191),
.B1(n_5277),
.B2(n_5148),
.Y(n_8931)
);

INVx2_ASAP7_75t_L g8932 ( 
.A(n_8585),
.Y(n_8932)
);

INVx1_ASAP7_75t_L g8933 ( 
.A(n_8598),
.Y(n_8933)
);

INVx1_ASAP7_75t_L g8934 ( 
.A(n_8598),
.Y(n_8934)
);

OAI22xp5_ASAP7_75t_L g8935 ( 
.A1(n_8720),
.A2(n_5321),
.B1(n_5399),
.B2(n_5336),
.Y(n_8935)
);

INVx2_ASAP7_75t_L g8936 ( 
.A(n_8565),
.Y(n_8936)
);

AOI32xp33_ASAP7_75t_L g8937 ( 
.A1(n_8723),
.A2(n_5354),
.A3(n_5314),
.B1(n_5878),
.B2(n_5857),
.Y(n_8937)
);

NOR2xp67_ASAP7_75t_L g8938 ( 
.A(n_8691),
.B(n_5685),
.Y(n_8938)
);

OAI22xp33_ASAP7_75t_SL g8939 ( 
.A1(n_8706),
.A2(n_5100),
.B1(n_5149),
.B2(n_4943),
.Y(n_8939)
);

INVxp67_ASAP7_75t_L g8940 ( 
.A(n_8726),
.Y(n_8940)
);

INVx1_ASAP7_75t_L g8941 ( 
.A(n_8645),
.Y(n_8941)
);

INVx1_ASAP7_75t_L g8942 ( 
.A(n_8645),
.Y(n_8942)
);

INVx1_ASAP7_75t_L g8943 ( 
.A(n_8649),
.Y(n_8943)
);

AND2x2_ASAP7_75t_L g8944 ( 
.A(n_8615),
.B(n_8559),
.Y(n_8944)
);

INVx2_ASAP7_75t_L g8945 ( 
.A(n_8764),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8649),
.Y(n_8946)
);

INVx1_ASAP7_75t_L g8947 ( 
.A(n_8653),
.Y(n_8947)
);

INVx2_ASAP7_75t_L g8948 ( 
.A(n_8736),
.Y(n_8948)
);

INVx1_ASAP7_75t_L g8949 ( 
.A(n_8653),
.Y(n_8949)
);

OAI322xp33_ASAP7_75t_L g8950 ( 
.A1(n_8590),
.A2(n_5439),
.A3(n_5450),
.B1(n_5446),
.B2(n_5485),
.C1(n_5474),
.C2(n_5471),
.Y(n_8950)
);

AOI22x1_ASAP7_75t_L g8951 ( 
.A1(n_8689),
.A2(n_8719),
.B1(n_8725),
.B2(n_8738),
.Y(n_8951)
);

INVx1_ASAP7_75t_SL g8952 ( 
.A(n_8708),
.Y(n_8952)
);

NAND2xp5_ASAP7_75t_L g8953 ( 
.A(n_8702),
.B(n_5689),
.Y(n_8953)
);

INVx2_ASAP7_75t_L g8954 ( 
.A(n_8635),
.Y(n_8954)
);

AND2x2_ASAP7_75t_L g8955 ( 
.A(n_8633),
.B(n_5817),
.Y(n_8955)
);

OAI22xp5_ASAP7_75t_L g8956 ( 
.A1(n_8616),
.A2(n_8745),
.B1(n_8755),
.B2(n_8740),
.Y(n_8956)
);

NAND2xp5_ASAP7_75t_L g8957 ( 
.A(n_8704),
.B(n_5689),
.Y(n_8957)
);

INVx1_ASAP7_75t_L g8958 ( 
.A(n_8656),
.Y(n_8958)
);

OAI22xp5_ASAP7_75t_L g8959 ( 
.A1(n_8568),
.A2(n_5336),
.B1(n_5399),
.B2(n_5321),
.Y(n_8959)
);

AOI32xp33_ASAP7_75t_L g8960 ( 
.A1(n_8714),
.A2(n_5364),
.A3(n_5323),
.B1(n_4875),
.B2(n_4910),
.Y(n_8960)
);

INVx1_ASAP7_75t_L g8961 ( 
.A(n_8656),
.Y(n_8961)
);

INVx1_ASAP7_75t_L g8962 ( 
.A(n_8581),
.Y(n_8962)
);

INVx1_ASAP7_75t_L g8963 ( 
.A(n_8596),
.Y(n_8963)
);

OAI222xp33_ASAP7_75t_L g8964 ( 
.A1(n_8717),
.A2(n_5791),
.B1(n_4941),
.B2(n_5149),
.C1(n_5151),
.C2(n_5100),
.Y(n_8964)
);

NAND2xp5_ASAP7_75t_L g8965 ( 
.A(n_8643),
.B(n_5693),
.Y(n_8965)
);

AOI21xp5_ASAP7_75t_L g8966 ( 
.A1(n_8677),
.A2(n_8679),
.B(n_8684),
.Y(n_8966)
);

INVx1_ASAP7_75t_L g8967 ( 
.A(n_8596),
.Y(n_8967)
);

OAI32xp33_ASAP7_75t_L g8968 ( 
.A1(n_8572),
.A2(n_5901),
.A3(n_5913),
.B1(n_5912),
.B2(n_5909),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_L g8969 ( 
.A(n_8647),
.B(n_5693),
.Y(n_8969)
);

OAI21xp33_ASAP7_75t_L g8970 ( 
.A1(n_8688),
.A2(n_5043),
.B(n_5004),
.Y(n_8970)
);

AND2x2_ASAP7_75t_L g8971 ( 
.A(n_8678),
.B(n_5820),
.Y(n_8971)
);

OAI22xp33_ASAP7_75t_SL g8972 ( 
.A1(n_8698),
.A2(n_5100),
.B1(n_5149),
.B2(n_4943),
.Y(n_8972)
);

INVxp67_ASAP7_75t_L g8973 ( 
.A(n_8669),
.Y(n_8973)
);

OAI22xp5_ASAP7_75t_L g8974 ( 
.A1(n_8749),
.A2(n_5336),
.B1(n_5399),
.B2(n_5321),
.Y(n_8974)
);

INVx1_ASAP7_75t_L g8975 ( 
.A(n_8574),
.Y(n_8975)
);

INVx1_ASAP7_75t_L g8976 ( 
.A(n_8675),
.Y(n_8976)
);

NAND2xp5_ASAP7_75t_L g8977 ( 
.A(n_8692),
.B(n_5694),
.Y(n_8977)
);

OAI21xp33_ASAP7_75t_L g8978 ( 
.A1(n_8674),
.A2(n_5046),
.B(n_5043),
.Y(n_8978)
);

AOI211xp5_ASAP7_75t_L g8979 ( 
.A1(n_8748),
.A2(n_5191),
.B(n_5277),
.C(n_5148),
.Y(n_8979)
);

INVx1_ASAP7_75t_L g8980 ( 
.A(n_8595),
.Y(n_8980)
);

O2A1O1Ixp33_ASAP7_75t_L g8981 ( 
.A1(n_8608),
.A2(n_6247),
.B(n_6256),
.C(n_6235),
.Y(n_8981)
);

INVxp67_ASAP7_75t_L g8982 ( 
.A(n_8591),
.Y(n_8982)
);

OR2x2_ASAP7_75t_L g8983 ( 
.A(n_8703),
.B(n_6316),
.Y(n_8983)
);

OAI22xp5_ASAP7_75t_L g8984 ( 
.A1(n_8753),
.A2(n_5399),
.B1(n_5364),
.B2(n_5323),
.Y(n_8984)
);

AOI22xp5_ASAP7_75t_L g8985 ( 
.A1(n_8629),
.A2(n_5191),
.B1(n_5277),
.B2(n_5148),
.Y(n_8985)
);

OR2x2_ASAP7_75t_L g8986 ( 
.A(n_8666),
.B(n_6336),
.Y(n_8986)
);

NOR2x1p5_ASAP7_75t_SL g8987 ( 
.A(n_8627),
.B(n_5658),
.Y(n_8987)
);

NAND3xp33_ASAP7_75t_L g8988 ( 
.A(n_8610),
.B(n_6249),
.C(n_6568),
.Y(n_8988)
);

NAND2x1p5_ASAP7_75t_L g8989 ( 
.A(n_8727),
.B(n_5057),
.Y(n_8989)
);

INVx2_ASAP7_75t_L g8990 ( 
.A(n_8636),
.Y(n_8990)
);

AND2x2_ASAP7_75t_L g8991 ( 
.A(n_8640),
.B(n_5820),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_8611),
.Y(n_8992)
);

NAND2xp5_ASAP7_75t_L g8993 ( 
.A(n_8742),
.B(n_5694),
.Y(n_8993)
);

AND2x2_ASAP7_75t_L g8994 ( 
.A(n_8612),
.B(n_5836),
.Y(n_8994)
);

INVx2_ASAP7_75t_L g8995 ( 
.A(n_8733),
.Y(n_8995)
);

OR2x2_ASAP7_75t_L g8996 ( 
.A(n_8681),
.B(n_6336),
.Y(n_8996)
);

INVx1_ASAP7_75t_L g8997 ( 
.A(n_8652),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_8665),
.Y(n_8998)
);

INVx1_ASAP7_75t_L g8999 ( 
.A(n_8624),
.Y(n_8999)
);

INVx1_ASAP7_75t_L g9000 ( 
.A(n_8762),
.Y(n_9000)
);

INVx1_ASAP7_75t_SL g9001 ( 
.A(n_8721),
.Y(n_9001)
);

AND2x4_ASAP7_75t_L g9002 ( 
.A(n_8814),
.B(n_8766),
.Y(n_9002)
);

AOI22xp33_ASAP7_75t_L g9003 ( 
.A1(n_8772),
.A2(n_8761),
.B1(n_8765),
.B2(n_8762),
.Y(n_9003)
);

AND2x4_ASAP7_75t_SL g9004 ( 
.A(n_8795),
.B(n_8765),
.Y(n_9004)
);

INVx1_ASAP7_75t_SL g9005 ( 
.A(n_8769),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8830),
.Y(n_9006)
);

INVx1_ASAP7_75t_L g9007 ( 
.A(n_8830),
.Y(n_9007)
);

AND2x2_ASAP7_75t_L g9008 ( 
.A(n_8794),
.B(n_8754),
.Y(n_9008)
);

INVx1_ASAP7_75t_L g9009 ( 
.A(n_8856),
.Y(n_9009)
);

AOI22xp33_ASAP7_75t_L g9010 ( 
.A1(n_8772),
.A2(n_8760),
.B1(n_8747),
.B2(n_8746),
.Y(n_9010)
);

OR2x2_ASAP7_75t_L g9011 ( 
.A(n_8825),
.B(n_8759),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_8775),
.Y(n_9012)
);

INVx1_ASAP7_75t_SL g9013 ( 
.A(n_8814),
.Y(n_9013)
);

BUFx2_ASAP7_75t_L g9014 ( 
.A(n_8783),
.Y(n_9014)
);

OAI21x1_ASAP7_75t_L g9015 ( 
.A1(n_8837),
.A2(n_8561),
.B(n_5565),
.Y(n_9015)
);

INVxp33_ASAP7_75t_SL g9016 ( 
.A(n_8793),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_8770),
.Y(n_9017)
);

INVx1_ASAP7_75t_L g9018 ( 
.A(n_8776),
.Y(n_9018)
);

INVx1_ASAP7_75t_SL g9019 ( 
.A(n_8809),
.Y(n_9019)
);

AOI22xp33_ASAP7_75t_L g9020 ( 
.A1(n_8768),
.A2(n_5191),
.B1(n_5277),
.B2(n_5148),
.Y(n_9020)
);

NAND2xp5_ASAP7_75t_L g9021 ( 
.A(n_8786),
.B(n_8561),
.Y(n_9021)
);

NAND2xp33_ASAP7_75t_SL g9022 ( 
.A(n_8899),
.B(n_5191),
.Y(n_9022)
);

INVx1_ASAP7_75t_L g9023 ( 
.A(n_8819),
.Y(n_9023)
);

AND2x2_ASAP7_75t_L g9024 ( 
.A(n_8802),
.B(n_5836),
.Y(n_9024)
);

OR2x6_ASAP7_75t_L g9025 ( 
.A(n_8903),
.B(n_5277),
.Y(n_9025)
);

AND2x2_ASAP7_75t_L g9026 ( 
.A(n_8810),
.B(n_8877),
.Y(n_9026)
);

NAND2xp33_ASAP7_75t_R g9027 ( 
.A(n_8783),
.B(n_8845),
.Y(n_9027)
);

OR2x2_ASAP7_75t_L g9028 ( 
.A(n_8839),
.B(n_6336),
.Y(n_9028)
);

NOR2xp33_ASAP7_75t_L g9029 ( 
.A(n_8767),
.B(n_5046),
.Y(n_9029)
);

NOR2xp33_ASAP7_75t_R g9030 ( 
.A(n_8791),
.B(n_5046),
.Y(n_9030)
);

AND2x4_ASAP7_75t_L g9031 ( 
.A(n_8817),
.B(n_5439),
.Y(n_9031)
);

OR2x2_ASAP7_75t_L g9032 ( 
.A(n_8847),
.B(n_5446),
.Y(n_9032)
);

INVxp67_ASAP7_75t_R g9033 ( 
.A(n_8883),
.Y(n_9033)
);

OR2x2_ASAP7_75t_L g9034 ( 
.A(n_8818),
.B(n_5450),
.Y(n_9034)
);

INVx1_ASAP7_75t_L g9035 ( 
.A(n_8874),
.Y(n_9035)
);

INVx1_ASAP7_75t_SL g9036 ( 
.A(n_8952),
.Y(n_9036)
);

INVx1_ASAP7_75t_L g9037 ( 
.A(n_8799),
.Y(n_9037)
);

NAND2xp5_ASAP7_75t_L g9038 ( 
.A(n_8808),
.B(n_5703),
.Y(n_9038)
);

AOI22xp33_ASAP7_75t_L g9039 ( 
.A1(n_8785),
.A2(n_5313),
.B1(n_5277),
.B2(n_5065),
.Y(n_9039)
);

AND2x2_ASAP7_75t_L g9040 ( 
.A(n_8860),
.B(n_5842),
.Y(n_9040)
);

HB1xp67_ASAP7_75t_L g9041 ( 
.A(n_8787),
.Y(n_9041)
);

INVx1_ASAP7_75t_L g9042 ( 
.A(n_8778),
.Y(n_9042)
);

INVx2_ASAP7_75t_L g9043 ( 
.A(n_8929),
.Y(n_9043)
);

INVx1_ASAP7_75t_L g9044 ( 
.A(n_8824),
.Y(n_9044)
);

INVxp67_ASAP7_75t_SL g9045 ( 
.A(n_8782),
.Y(n_9045)
);

INVx1_ASAP7_75t_L g9046 ( 
.A(n_8826),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8869),
.Y(n_9047)
);

INVx1_ASAP7_75t_L g9048 ( 
.A(n_8834),
.Y(n_9048)
);

INVx1_ASAP7_75t_L g9049 ( 
.A(n_8944),
.Y(n_9049)
);

NAND2xp5_ASAP7_75t_L g9050 ( 
.A(n_8913),
.B(n_8828),
.Y(n_9050)
);

NOR2xp33_ASAP7_75t_L g9051 ( 
.A(n_8784),
.B(n_5059),
.Y(n_9051)
);

AND2x4_ASAP7_75t_SL g9052 ( 
.A(n_8780),
.B(n_5313),
.Y(n_9052)
);

AND2x4_ASAP7_75t_L g9053 ( 
.A(n_8867),
.B(n_5471),
.Y(n_9053)
);

AND2x2_ASAP7_75t_SL g9054 ( 
.A(n_8924),
.B(n_5057),
.Y(n_9054)
);

INVx2_ASAP7_75t_L g9055 ( 
.A(n_8902),
.Y(n_9055)
);

INVx2_ASAP7_75t_L g9056 ( 
.A(n_8910),
.Y(n_9056)
);

INVxp67_ASAP7_75t_L g9057 ( 
.A(n_8836),
.Y(n_9057)
);

INVx2_ASAP7_75t_L g9058 ( 
.A(n_8858),
.Y(n_9058)
);

INVx2_ASAP7_75t_L g9059 ( 
.A(n_8888),
.Y(n_9059)
);

INVx1_ASAP7_75t_L g9060 ( 
.A(n_8815),
.Y(n_9060)
);

NOR2x1_ASAP7_75t_L g9061 ( 
.A(n_8843),
.B(n_8811),
.Y(n_9061)
);

AND2x2_ASAP7_75t_L g9062 ( 
.A(n_8838),
.B(n_5842),
.Y(n_9062)
);

INVx1_ASAP7_75t_L g9063 ( 
.A(n_8816),
.Y(n_9063)
);

INVx1_ASAP7_75t_L g9064 ( 
.A(n_8827),
.Y(n_9064)
);

AO21x2_ASAP7_75t_L g9065 ( 
.A1(n_8773),
.A2(n_6351),
.B(n_6337),
.Y(n_9065)
);

INVx2_ASAP7_75t_L g9066 ( 
.A(n_8923),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8788),
.Y(n_9067)
);

NOR2xp33_ASAP7_75t_L g9068 ( 
.A(n_8922),
.B(n_5059),
.Y(n_9068)
);

NAND2xp5_ASAP7_75t_L g9069 ( 
.A(n_8789),
.B(n_5703),
.Y(n_9069)
);

OR2x2_ASAP7_75t_L g9070 ( 
.A(n_8797),
.B(n_5474),
.Y(n_9070)
);

INVx1_ASAP7_75t_L g9071 ( 
.A(n_8822),
.Y(n_9071)
);

INVx2_ASAP7_75t_SL g9072 ( 
.A(n_8887),
.Y(n_9072)
);

OR2x2_ASAP7_75t_L g9073 ( 
.A(n_8932),
.B(n_5485),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_8777),
.Y(n_9074)
);

INVx2_ASAP7_75t_L g9075 ( 
.A(n_8914),
.Y(n_9075)
);

AND2x2_ASAP7_75t_L g9076 ( 
.A(n_8945),
.B(n_5850),
.Y(n_9076)
);

NAND2xp5_ASAP7_75t_L g9077 ( 
.A(n_8835),
.B(n_5706),
.Y(n_9077)
);

INVx1_ASAP7_75t_SL g9078 ( 
.A(n_8876),
.Y(n_9078)
);

AOI22xp33_ASAP7_75t_L g9079 ( 
.A1(n_8803),
.A2(n_5313),
.B1(n_5065),
.B2(n_5059),
.Y(n_9079)
);

INVx1_ASAP7_75t_L g9080 ( 
.A(n_8773),
.Y(n_9080)
);

AOI22xp33_ASAP7_75t_L g9081 ( 
.A1(n_8774),
.A2(n_5313),
.B1(n_5065),
.B2(n_6405),
.Y(n_9081)
);

OAI221xp5_ASAP7_75t_L g9082 ( 
.A1(n_8904),
.A2(n_5151),
.B1(n_5331),
.B2(n_5268),
.C(n_4943),
.Y(n_9082)
);

INVx1_ASAP7_75t_L g9083 ( 
.A(n_8850),
.Y(n_9083)
);

NOR2xp33_ASAP7_75t_L g9084 ( 
.A(n_8833),
.B(n_5313),
.Y(n_9084)
);

INVx3_ASAP7_75t_L g9085 ( 
.A(n_8905),
.Y(n_9085)
);

AOI22xp5_ASAP7_75t_L g9086 ( 
.A1(n_8821),
.A2(n_5313),
.B1(n_5399),
.B2(n_5028),
.Y(n_9086)
);

NAND2xp5_ASAP7_75t_L g9087 ( 
.A(n_8954),
.B(n_5706),
.Y(n_9087)
);

AO21x2_ASAP7_75t_L g9088 ( 
.A1(n_8813),
.A2(n_6337),
.B(n_6351),
.Y(n_9088)
);

INVx1_ASAP7_75t_L g9089 ( 
.A(n_8820),
.Y(n_9089)
);

AND2x2_ASAP7_75t_L g9090 ( 
.A(n_8851),
.B(n_5850),
.Y(n_9090)
);

HB1xp67_ASAP7_75t_L g9091 ( 
.A(n_8911),
.Y(n_9091)
);

INVxp67_ASAP7_75t_SL g9092 ( 
.A(n_8779),
.Y(n_9092)
);

AND2x2_ASAP7_75t_L g9093 ( 
.A(n_8882),
.B(n_5867),
.Y(n_9093)
);

CKINVDCx16_ASAP7_75t_R g9094 ( 
.A(n_8891),
.Y(n_9094)
);

INVx1_ASAP7_75t_SL g9095 ( 
.A(n_9001),
.Y(n_9095)
);

BUFx3_ASAP7_75t_L g9096 ( 
.A(n_8990),
.Y(n_9096)
);

AND2x2_ASAP7_75t_L g9097 ( 
.A(n_8840),
.B(n_5867),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_8853),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_8925),
.Y(n_9099)
);

INVx3_ASAP7_75t_L g9100 ( 
.A(n_8936),
.Y(n_9100)
);

INVx1_ASAP7_75t_SL g9101 ( 
.A(n_8927),
.Y(n_9101)
);

INVx4_ASAP7_75t_L g9102 ( 
.A(n_9000),
.Y(n_9102)
);

AND2x2_ASAP7_75t_L g9103 ( 
.A(n_8873),
.B(n_5874),
.Y(n_9103)
);

BUFx3_ASAP7_75t_L g9104 ( 
.A(n_8865),
.Y(n_9104)
);

INVx1_ASAP7_75t_SL g9105 ( 
.A(n_8948),
.Y(n_9105)
);

NOR2x1_ASAP7_75t_L g9106 ( 
.A(n_8771),
.B(n_6495),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_8926),
.Y(n_9107)
);

NAND2xp5_ASAP7_75t_L g9108 ( 
.A(n_8921),
.B(n_5714),
.Y(n_9108)
);

INVx1_ASAP7_75t_SL g9109 ( 
.A(n_8995),
.Y(n_9109)
);

OR2x2_ASAP7_75t_L g9110 ( 
.A(n_8866),
.B(n_5488),
.Y(n_9110)
);

INVx1_ASAP7_75t_L g9111 ( 
.A(n_8933),
.Y(n_9111)
);

NAND2xp5_ASAP7_75t_L g9112 ( 
.A(n_8928),
.B(n_5714),
.Y(n_9112)
);

NOR2xp33_ASAP7_75t_L g9113 ( 
.A(n_8982),
.B(n_5057),
.Y(n_9113)
);

HB1xp67_ASAP7_75t_L g9114 ( 
.A(n_8771),
.Y(n_9114)
);

INVx1_ASAP7_75t_L g9115 ( 
.A(n_8934),
.Y(n_9115)
);

NOR2xp33_ASAP7_75t_L g9116 ( 
.A(n_8940),
.B(n_5057),
.Y(n_9116)
);

INVx1_ASAP7_75t_L g9117 ( 
.A(n_8941),
.Y(n_9117)
);

INVx2_ASAP7_75t_L g9118 ( 
.A(n_8951),
.Y(n_9118)
);

CKINVDCx16_ASAP7_75t_R g9119 ( 
.A(n_8831),
.Y(n_9119)
);

INVx1_ASAP7_75t_SL g9120 ( 
.A(n_8980),
.Y(n_9120)
);

AND2x2_ASAP7_75t_L g9121 ( 
.A(n_8781),
.B(n_8864),
.Y(n_9121)
);

OR2x6_ASAP7_75t_L g9122 ( 
.A(n_8861),
.B(n_5151),
.Y(n_9122)
);

INVxp67_ASAP7_75t_L g9123 ( 
.A(n_8919),
.Y(n_9123)
);

NAND2xp5_ASAP7_75t_L g9124 ( 
.A(n_8896),
.B(n_5715),
.Y(n_9124)
);

AND2x2_ASAP7_75t_L g9125 ( 
.A(n_8832),
.B(n_5874),
.Y(n_9125)
);

BUFx3_ASAP7_75t_L g9126 ( 
.A(n_8862),
.Y(n_9126)
);

INVx2_ASAP7_75t_L g9127 ( 
.A(n_8951),
.Y(n_9127)
);

HB1xp67_ASAP7_75t_L g9128 ( 
.A(n_8800),
.Y(n_9128)
);

INVx1_ASAP7_75t_L g9129 ( 
.A(n_8942),
.Y(n_9129)
);

INVx1_ASAP7_75t_L g9130 ( 
.A(n_8943),
.Y(n_9130)
);

OAI22xp5_ASAP7_75t_L g9131 ( 
.A1(n_8804),
.A2(n_5491),
.B1(n_5494),
.B2(n_5488),
.Y(n_9131)
);

INVx1_ASAP7_75t_L g9132 ( 
.A(n_8946),
.Y(n_9132)
);

HB1xp67_ASAP7_75t_L g9133 ( 
.A(n_8801),
.Y(n_9133)
);

AOI22x1_ASAP7_75t_L g9134 ( 
.A1(n_8807),
.A2(n_5268),
.B1(n_5331),
.B2(n_5491),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_8855),
.Y(n_9135)
);

INVx1_ASAP7_75t_SL g9136 ( 
.A(n_8879),
.Y(n_9136)
);

NAND2xp5_ASAP7_75t_L g9137 ( 
.A(n_8790),
.B(n_5715),
.Y(n_9137)
);

HB1xp67_ASAP7_75t_L g9138 ( 
.A(n_8812),
.Y(n_9138)
);

AND2x4_ASAP7_75t_L g9139 ( 
.A(n_8872),
.B(n_5494),
.Y(n_9139)
);

NAND2xp5_ASAP7_75t_L g9140 ( 
.A(n_8823),
.B(n_5716),
.Y(n_9140)
);

OR2x2_ASAP7_75t_L g9141 ( 
.A(n_8841),
.B(n_5495),
.Y(n_9141)
);

INVx2_ASAP7_75t_L g9142 ( 
.A(n_8917),
.Y(n_9142)
);

INVx3_ASAP7_75t_L g9143 ( 
.A(n_8881),
.Y(n_9143)
);

INVx2_ASAP7_75t_SL g9144 ( 
.A(n_8890),
.Y(n_9144)
);

AND2x2_ASAP7_75t_L g9145 ( 
.A(n_8805),
.B(n_8798),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_8989),
.Y(n_9146)
);

INVx1_ASAP7_75t_L g9147 ( 
.A(n_8947),
.Y(n_9147)
);

INVx1_ASAP7_75t_L g9148 ( 
.A(n_8949),
.Y(n_9148)
);

AND2x2_ASAP7_75t_SL g9149 ( 
.A(n_8848),
.B(n_8999),
.Y(n_9149)
);

INVx1_ASAP7_75t_SL g9150 ( 
.A(n_8863),
.Y(n_9150)
);

AND2x2_ASAP7_75t_L g9151 ( 
.A(n_8973),
.B(n_5875),
.Y(n_9151)
);

NAND2xp5_ASAP7_75t_L g9152 ( 
.A(n_8806),
.B(n_5716),
.Y(n_9152)
);

NAND2xp5_ASAP7_75t_L g9153 ( 
.A(n_8966),
.B(n_5717),
.Y(n_9153)
);

OAI22xp5_ASAP7_75t_L g9154 ( 
.A1(n_8846),
.A2(n_5495),
.B1(n_5508),
.B2(n_5497),
.Y(n_9154)
);

INVx1_ASAP7_75t_SL g9155 ( 
.A(n_8857),
.Y(n_9155)
);

OR2x2_ASAP7_75t_L g9156 ( 
.A(n_8956),
.B(n_5497),
.Y(n_9156)
);

INVx1_ASAP7_75t_L g9157 ( 
.A(n_8958),
.Y(n_9157)
);

INVx1_ASAP7_75t_L g9158 ( 
.A(n_8961),
.Y(n_9158)
);

NAND2xp5_ASAP7_75t_L g9159 ( 
.A(n_8792),
.B(n_5717),
.Y(n_9159)
);

BUFx3_ASAP7_75t_L g9160 ( 
.A(n_8976),
.Y(n_9160)
);

INVx1_ASAP7_75t_L g9161 ( 
.A(n_8907),
.Y(n_9161)
);

NOR2x1_ASAP7_75t_L g9162 ( 
.A(n_8963),
.B(n_6495),
.Y(n_9162)
);

NAND2xp33_ASAP7_75t_SL g9163 ( 
.A(n_8880),
.B(n_5399),
.Y(n_9163)
);

INVx2_ASAP7_75t_L g9164 ( 
.A(n_8971),
.Y(n_9164)
);

INVx4_ASAP7_75t_L g9165 ( 
.A(n_8967),
.Y(n_9165)
);

INVx1_ASAP7_75t_L g9166 ( 
.A(n_8916),
.Y(n_9166)
);

INVx1_ASAP7_75t_L g9167 ( 
.A(n_8885),
.Y(n_9167)
);

AND2x2_ASAP7_75t_L g9168 ( 
.A(n_8962),
.B(n_5875),
.Y(n_9168)
);

INVx4_ASAP7_75t_L g9169 ( 
.A(n_8975),
.Y(n_9169)
);

AND2x2_ASAP7_75t_L g9170 ( 
.A(n_8998),
.B(n_5880),
.Y(n_9170)
);

AOI22xp33_ASAP7_75t_L g9171 ( 
.A1(n_8829),
.A2(n_6405),
.B1(n_5796),
.B2(n_5798),
.Y(n_9171)
);

INVx1_ASAP7_75t_L g9172 ( 
.A(n_8889),
.Y(n_9172)
);

OR2x2_ASAP7_75t_L g9173 ( 
.A(n_8870),
.B(n_5508),
.Y(n_9173)
);

INVx2_ASAP7_75t_L g9174 ( 
.A(n_8991),
.Y(n_9174)
);

INVx1_ASAP7_75t_L g9175 ( 
.A(n_8893),
.Y(n_9175)
);

OR2x2_ASAP7_75t_L g9176 ( 
.A(n_8997),
.B(n_5512),
.Y(n_9176)
);

NAND2xp5_ASAP7_75t_L g9177 ( 
.A(n_8992),
.B(n_5719),
.Y(n_9177)
);

AOI22xp33_ASAP7_75t_SL g9178 ( 
.A1(n_8796),
.A2(n_6352),
.B1(n_5028),
.B2(n_5376),
.Y(n_9178)
);

INVx1_ASAP7_75t_SL g9179 ( 
.A(n_8955),
.Y(n_9179)
);

AND2x2_ASAP7_75t_L g9180 ( 
.A(n_8895),
.B(n_5880),
.Y(n_9180)
);

INVx1_ASAP7_75t_L g9181 ( 
.A(n_8987),
.Y(n_9181)
);

NAND2xp5_ASAP7_75t_L g9182 ( 
.A(n_8970),
.B(n_5719),
.Y(n_9182)
);

INVx1_ASAP7_75t_SL g9183 ( 
.A(n_8871),
.Y(n_9183)
);

AND2x2_ASAP7_75t_L g9184 ( 
.A(n_8978),
.B(n_5885),
.Y(n_9184)
);

AOI22xp33_ASAP7_75t_L g9185 ( 
.A1(n_8859),
.A2(n_6405),
.B1(n_5798),
.B2(n_6352),
.Y(n_9185)
);

OR2x2_ASAP7_75t_L g9186 ( 
.A(n_8892),
.B(n_5512),
.Y(n_9186)
);

INVx1_ASAP7_75t_L g9187 ( 
.A(n_8897),
.Y(n_9187)
);

INVx1_ASAP7_75t_L g9188 ( 
.A(n_8898),
.Y(n_9188)
);

NAND2xp5_ASAP7_75t_L g9189 ( 
.A(n_8994),
.B(n_5724),
.Y(n_9189)
);

INVx6_ASAP7_75t_L g9190 ( 
.A(n_8884),
.Y(n_9190)
);

INVx1_ASAP7_75t_SL g9191 ( 
.A(n_8875),
.Y(n_9191)
);

AND2x2_ASAP7_75t_L g9192 ( 
.A(n_8844),
.B(n_5885),
.Y(n_9192)
);

INVx1_ASAP7_75t_SL g9193 ( 
.A(n_8894),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_9014),
.Y(n_9194)
);

INVx1_ASAP7_75t_L g9195 ( 
.A(n_9114),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_SL g9196 ( 
.A(n_9013),
.B(n_8931),
.Y(n_9196)
);

AOI21xp5_ASAP7_75t_L g9197 ( 
.A1(n_9057),
.A2(n_8920),
.B(n_8900),
.Y(n_9197)
);

AOI22xp33_ASAP7_75t_L g9198 ( 
.A1(n_9092),
.A2(n_8842),
.B1(n_8908),
.B2(n_8909),
.Y(n_9198)
);

NAND2xp5_ASAP7_75t_L g9199 ( 
.A(n_9006),
.B(n_8901),
.Y(n_9199)
);

INVx1_ASAP7_75t_L g9200 ( 
.A(n_9181),
.Y(n_9200)
);

OAI21xp33_ASAP7_75t_L g9201 ( 
.A1(n_9016),
.A2(n_8852),
.B(n_8906),
.Y(n_9201)
);

AND2x2_ASAP7_75t_L g9202 ( 
.A(n_9033),
.B(n_8979),
.Y(n_9202)
);

OAI22xp5_ASAP7_75t_L g9203 ( 
.A1(n_9005),
.A2(n_8985),
.B1(n_8854),
.B2(n_8912),
.Y(n_9203)
);

INVx1_ASAP7_75t_L g9204 ( 
.A(n_9181),
.Y(n_9204)
);

AND2x2_ASAP7_75t_L g9205 ( 
.A(n_9026),
.B(n_8938),
.Y(n_9205)
);

NOR2xp33_ASAP7_75t_L g9206 ( 
.A(n_9094),
.B(n_8886),
.Y(n_9206)
);

OAI221xp5_ASAP7_75t_L g9207 ( 
.A1(n_9003),
.A2(n_8960),
.B1(n_8984),
.B2(n_8953),
.C(n_8957),
.Y(n_9207)
);

OAI22xp5_ASAP7_75t_L g9208 ( 
.A1(n_9039),
.A2(n_8915),
.B1(n_8969),
.B2(n_8965),
.Y(n_9208)
);

AND2x2_ASAP7_75t_L g9209 ( 
.A(n_9017),
.B(n_8977),
.Y(n_9209)
);

INVx1_ASAP7_75t_L g9210 ( 
.A(n_9007),
.Y(n_9210)
);

OAI22xp5_ASAP7_75t_L g9211 ( 
.A1(n_9081),
.A2(n_9086),
.B1(n_9079),
.B2(n_9045),
.Y(n_9211)
);

INVx2_ASAP7_75t_L g9212 ( 
.A(n_9002),
.Y(n_9212)
);

INVx1_ASAP7_75t_L g9213 ( 
.A(n_9002),
.Y(n_9213)
);

NAND3xp33_ASAP7_75t_L g9214 ( 
.A(n_9027),
.B(n_8996),
.C(n_8986),
.Y(n_9214)
);

AND2x2_ASAP7_75t_L g9215 ( 
.A(n_9023),
.B(n_8993),
.Y(n_9215)
);

NOR3xp33_ASAP7_75t_L g9216 ( 
.A(n_9050),
.B(n_8974),
.C(n_8935),
.Y(n_9216)
);

INVx2_ASAP7_75t_L g9217 ( 
.A(n_9004),
.Y(n_9217)
);

INVx1_ASAP7_75t_L g9218 ( 
.A(n_9091),
.Y(n_9218)
);

INVx1_ASAP7_75t_L g9219 ( 
.A(n_9009),
.Y(n_9219)
);

INVx1_ASAP7_75t_L g9220 ( 
.A(n_9085),
.Y(n_9220)
);

INVx2_ASAP7_75t_SL g9221 ( 
.A(n_9025),
.Y(n_9221)
);

NAND2xp5_ASAP7_75t_L g9222 ( 
.A(n_9085),
.B(n_8937),
.Y(n_9222)
);

INVx1_ASAP7_75t_L g9223 ( 
.A(n_9100),
.Y(n_9223)
);

HB1xp67_ASAP7_75t_L g9224 ( 
.A(n_9025),
.Y(n_9224)
);

NAND2xp5_ASAP7_75t_L g9225 ( 
.A(n_9019),
.B(n_8959),
.Y(n_9225)
);

NAND2xp5_ASAP7_75t_SL g9226 ( 
.A(n_9100),
.B(n_8939),
.Y(n_9226)
);

OAI21xp33_ASAP7_75t_L g9227 ( 
.A1(n_9036),
.A2(n_8972),
.B(n_8983),
.Y(n_9227)
);

INVx1_ASAP7_75t_L g9228 ( 
.A(n_9041),
.Y(n_9228)
);

AOI22xp33_ASAP7_75t_L g9229 ( 
.A1(n_9126),
.A2(n_8988),
.B1(n_8950),
.B2(n_8849),
.Y(n_9229)
);

INVx1_ASAP7_75t_L g9230 ( 
.A(n_9096),
.Y(n_9230)
);

NAND2xp5_ASAP7_75t_L g9231 ( 
.A(n_9109),
.B(n_9119),
.Y(n_9231)
);

NAND2xp5_ASAP7_75t_SL g9232 ( 
.A(n_9095),
.B(n_8981),
.Y(n_9232)
);

NAND2xp33_ASAP7_75t_SL g9233 ( 
.A(n_9030),
.B(n_8868),
.Y(n_9233)
);

INVx2_ASAP7_75t_L g9234 ( 
.A(n_9059),
.Y(n_9234)
);

INVx1_ASAP7_75t_L g9235 ( 
.A(n_9035),
.Y(n_9235)
);

OR2x2_ASAP7_75t_L g9236 ( 
.A(n_9105),
.B(n_8878),
.Y(n_9236)
);

AOI22xp5_ASAP7_75t_L g9237 ( 
.A1(n_9051),
.A2(n_8868),
.B1(n_6495),
.B2(n_6505),
.Y(n_9237)
);

AOI21xp33_ASAP7_75t_SL g9238 ( 
.A1(n_9144),
.A2(n_8930),
.B(n_8918),
.Y(n_9238)
);

NOR2xp33_ASAP7_75t_SL g9239 ( 
.A(n_9120),
.B(n_8964),
.Y(n_9239)
);

AOI22xp5_ASAP7_75t_L g9240 ( 
.A1(n_9121),
.A2(n_6505),
.B1(n_6447),
.B2(n_5376),
.Y(n_9240)
);

NOR2x1_ASAP7_75t_L g9241 ( 
.A(n_9118),
.B(n_8918),
.Y(n_9241)
);

AND2x2_ASAP7_75t_L g9242 ( 
.A(n_9008),
.B(n_8930),
.Y(n_9242)
);

OAI22xp5_ASAP7_75t_L g9243 ( 
.A1(n_9020),
.A2(n_5515),
.B1(n_5531),
.B2(n_5520),
.Y(n_9243)
);

AOI221xp5_ASAP7_75t_L g9244 ( 
.A1(n_9127),
.A2(n_8968),
.B1(n_6505),
.B2(n_6447),
.C(n_6353),
.Y(n_9244)
);

AOI21xp5_ASAP7_75t_L g9245 ( 
.A1(n_9106),
.A2(n_8968),
.B(n_6351),
.Y(n_9245)
);

INVx2_ASAP7_75t_L g9246 ( 
.A(n_9043),
.Y(n_9246)
);

OAI221xp5_ASAP7_75t_L g9247 ( 
.A1(n_9178),
.A2(n_5331),
.B1(n_5268),
.B2(n_4941),
.C(n_6568),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_9049),
.Y(n_9248)
);

OR2x2_ASAP7_75t_L g9249 ( 
.A(n_9055),
.B(n_5658),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_9047),
.Y(n_9250)
);

AOI21xp33_ASAP7_75t_L g9251 ( 
.A1(n_9011),
.A2(n_6447),
.B(n_6353),
.Y(n_9251)
);

AND2x2_ASAP7_75t_L g9252 ( 
.A(n_9058),
.B(n_5889),
.Y(n_9252)
);

NAND2xp5_ASAP7_75t_SL g9253 ( 
.A(n_9071),
.B(n_5515),
.Y(n_9253)
);

AOI21xp33_ASAP7_75t_L g9254 ( 
.A1(n_9116),
.A2(n_6353),
.B(n_6337),
.Y(n_9254)
);

OR2x2_ASAP7_75t_L g9255 ( 
.A(n_9056),
.B(n_5658),
.Y(n_9255)
);

OAI22xp5_ASAP7_75t_L g9256 ( 
.A1(n_9082),
.A2(n_5520),
.B1(n_5541),
.B2(n_5531),
.Y(n_9256)
);

AND2x2_ASAP7_75t_L g9257 ( 
.A(n_9075),
.B(n_5889),
.Y(n_9257)
);

OAI22xp5_ASAP7_75t_L g9258 ( 
.A1(n_9012),
.A2(n_5541),
.B1(n_5547),
.B2(n_5545),
.Y(n_9258)
);

OR2x2_ASAP7_75t_L g9259 ( 
.A(n_9066),
.B(n_5660),
.Y(n_9259)
);

NAND2xp5_ASAP7_75t_L g9260 ( 
.A(n_9072),
.B(n_5724),
.Y(n_9260)
);

INVx1_ASAP7_75t_L g9261 ( 
.A(n_9061),
.Y(n_9261)
);

OAI22xp5_ASAP7_75t_L g9262 ( 
.A1(n_9101),
.A2(n_9037),
.B1(n_9018),
.B2(n_9142),
.Y(n_9262)
);

NAND2xp33_ASAP7_75t_L g9263 ( 
.A(n_9128),
.B(n_5895),
.Y(n_9263)
);

NAND2xp5_ASAP7_75t_L g9264 ( 
.A(n_9179),
.B(n_9042),
.Y(n_9264)
);

AOI22xp5_ASAP7_75t_L g9265 ( 
.A1(n_9029),
.A2(n_5219),
.B1(n_5798),
.B2(n_6375),
.Y(n_9265)
);

AOI221xp5_ASAP7_75t_L g9266 ( 
.A1(n_9131),
.A2(n_6375),
.B1(n_5664),
.B2(n_5669),
.C(n_5661),
.Y(n_9266)
);

INVx1_ASAP7_75t_L g9267 ( 
.A(n_9133),
.Y(n_9267)
);

INVx1_ASAP7_75t_L g9268 ( 
.A(n_9138),
.Y(n_9268)
);

AO21x1_ASAP7_75t_L g9269 ( 
.A1(n_9102),
.A2(n_5661),
.B(n_5660),
.Y(n_9269)
);

NAND2xp5_ASAP7_75t_L g9270 ( 
.A(n_9135),
.B(n_5726),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_9021),
.Y(n_9271)
);

INVx1_ASAP7_75t_L g9272 ( 
.A(n_9080),
.Y(n_9272)
);

NAND2xp5_ASAP7_75t_L g9273 ( 
.A(n_9052),
.B(n_5726),
.Y(n_9273)
);

AOI322xp5_ASAP7_75t_L g9274 ( 
.A1(n_9145),
.A2(n_9113),
.A3(n_9137),
.B1(n_9140),
.B2(n_9159),
.C1(n_9068),
.C2(n_9060),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_9104),
.Y(n_9275)
);

INVx1_ASAP7_75t_L g9276 ( 
.A(n_9190),
.Y(n_9276)
);

NOR2x1_ASAP7_75t_L g9277 ( 
.A(n_9102),
.B(n_6375),
.Y(n_9277)
);

NAND2xp5_ASAP7_75t_SL g9278 ( 
.A(n_9169),
.B(n_5545),
.Y(n_9278)
);

INVxp67_ASAP7_75t_L g9279 ( 
.A(n_9084),
.Y(n_9279)
);

OR2x2_ASAP7_75t_L g9280 ( 
.A(n_9083),
.B(n_9164),
.Y(n_9280)
);

NAND3xp33_ASAP7_75t_L g9281 ( 
.A(n_9010),
.B(n_6568),
.C(n_6352),
.Y(n_9281)
);

INVx1_ASAP7_75t_L g9282 ( 
.A(n_9190),
.Y(n_9282)
);

NOR2xp33_ASAP7_75t_SL g9283 ( 
.A(n_9169),
.B(n_4231),
.Y(n_9283)
);

NOR2x1_ASAP7_75t_L g9284 ( 
.A(n_9165),
.B(n_9187),
.Y(n_9284)
);

INVx1_ASAP7_75t_L g9285 ( 
.A(n_9048),
.Y(n_9285)
);

OR2x2_ASAP7_75t_L g9286 ( 
.A(n_9174),
.B(n_5660),
.Y(n_9286)
);

INVxp67_ASAP7_75t_SL g9287 ( 
.A(n_9187),
.Y(n_9287)
);

NOR2x1_ASAP7_75t_L g9288 ( 
.A(n_9165),
.B(n_5547),
.Y(n_9288)
);

HB1xp67_ASAP7_75t_L g9289 ( 
.A(n_9188),
.Y(n_9289)
);

OAI22xp5_ASAP7_75t_L g9290 ( 
.A1(n_9078),
.A2(n_5550),
.B1(n_5559),
.B2(n_5552),
.Y(n_9290)
);

INVx1_ASAP7_75t_L g9291 ( 
.A(n_9063),
.Y(n_9291)
);

INVx1_ASAP7_75t_L g9292 ( 
.A(n_9064),
.Y(n_9292)
);

OAI221xp5_ASAP7_75t_L g9293 ( 
.A1(n_9123),
.A2(n_5219),
.B1(n_3754),
.B2(n_4268),
.C(n_5244),
.Y(n_9293)
);

AOI21xp5_ASAP7_75t_L g9294 ( 
.A1(n_9054),
.A2(n_5552),
.B(n_5550),
.Y(n_9294)
);

NAND2xp5_ASAP7_75t_L g9295 ( 
.A(n_9067),
.B(n_5734),
.Y(n_9295)
);

AOI21xp5_ASAP7_75t_L g9296 ( 
.A1(n_9022),
.A2(n_5577),
.B(n_5559),
.Y(n_9296)
);

INVx3_ASAP7_75t_L g9297 ( 
.A(n_9031),
.Y(n_9297)
);

INVx1_ASAP7_75t_L g9298 ( 
.A(n_9188),
.Y(n_9298)
);

AND2x2_ASAP7_75t_L g9299 ( 
.A(n_9044),
.B(n_5895),
.Y(n_9299)
);

AOI21xp5_ASAP7_75t_L g9300 ( 
.A1(n_9153),
.A2(n_5578),
.B(n_5576),
.Y(n_9300)
);

OAI221xp5_ASAP7_75t_L g9301 ( 
.A1(n_9141),
.A2(n_3754),
.B1(n_4268),
.B2(n_5244),
.C(n_4367),
.Y(n_9301)
);

INVx1_ASAP7_75t_L g9302 ( 
.A(n_9098),
.Y(n_9302)
);

INVx1_ASAP7_75t_L g9303 ( 
.A(n_9180),
.Y(n_9303)
);

AOI22xp5_ASAP7_75t_L g9304 ( 
.A1(n_9074),
.A2(n_5577),
.B1(n_5578),
.B2(n_5576),
.Y(n_9304)
);

XNOR2xp5_ASAP7_75t_L g9305 ( 
.A(n_9149),
.B(n_5791),
.Y(n_9305)
);

NAND2xp5_ASAP7_75t_SL g9306 ( 
.A(n_9031),
.B(n_5664),
.Y(n_9306)
);

OAI21xp33_ASAP7_75t_SL g9307 ( 
.A1(n_9015),
.A2(n_5565),
.B(n_5564),
.Y(n_9307)
);

OAI22xp33_ASAP7_75t_L g9308 ( 
.A1(n_9122),
.A2(n_5903),
.B1(n_5909),
.B2(n_5830),
.Y(n_9308)
);

AOI32xp33_ASAP7_75t_L g9309 ( 
.A1(n_9046),
.A2(n_4898),
.A3(n_4910),
.B1(n_4875),
.B2(n_4853),
.Y(n_9309)
);

NOR2xp33_ASAP7_75t_L g9310 ( 
.A(n_9150),
.B(n_5896),
.Y(n_9310)
);

INVx1_ASAP7_75t_L g9311 ( 
.A(n_9143),
.Y(n_9311)
);

XNOR2xp5_ASAP7_75t_L g9312 ( 
.A(n_9183),
.B(n_5288),
.Y(n_9312)
);

AOI22xp5_ASAP7_75t_L g9313 ( 
.A1(n_9146),
.A2(n_5664),
.B1(n_5669),
.B2(n_5661),
.Y(n_9313)
);

AOI21xp5_ASAP7_75t_L g9314 ( 
.A1(n_9163),
.A2(n_5673),
.B(n_5669),
.Y(n_9314)
);

AND2x2_ASAP7_75t_L g9315 ( 
.A(n_9160),
.B(n_5896),
.Y(n_9315)
);

INVx3_ASAP7_75t_L g9316 ( 
.A(n_9053),
.Y(n_9316)
);

INVx1_ASAP7_75t_L g9317 ( 
.A(n_9143),
.Y(n_9317)
);

NAND2xp5_ASAP7_75t_L g9318 ( 
.A(n_9062),
.B(n_5734),
.Y(n_9318)
);

INVx2_ASAP7_75t_L g9319 ( 
.A(n_9122),
.Y(n_9319)
);

AOI22xp5_ASAP7_75t_L g9320 ( 
.A1(n_9089),
.A2(n_9191),
.B1(n_9193),
.B2(n_9024),
.Y(n_9320)
);

AND2x2_ASAP7_75t_L g9321 ( 
.A(n_9090),
.B(n_5944),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_9161),
.Y(n_9322)
);

NAND2xp5_ASAP7_75t_L g9323 ( 
.A(n_9040),
.B(n_5739),
.Y(n_9323)
);

OAI32xp33_ASAP7_75t_L g9324 ( 
.A1(n_9152),
.A2(n_5942),
.A3(n_5913),
.B1(n_5919),
.B2(n_5912),
.Y(n_9324)
);

INVx1_ASAP7_75t_L g9325 ( 
.A(n_9166),
.Y(n_9325)
);

OAI221xp5_ASAP7_75t_L g9326 ( 
.A1(n_9108),
.A2(n_3754),
.B1(n_4268),
.B2(n_4367),
.C(n_4366),
.Y(n_9326)
);

INVx2_ASAP7_75t_L g9327 ( 
.A(n_9053),
.Y(n_9327)
);

AND2x2_ASAP7_75t_L g9328 ( 
.A(n_9093),
.B(n_5944),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_9099),
.Y(n_9329)
);

NAND2xp5_ASAP7_75t_L g9330 ( 
.A(n_9103),
.B(n_5739),
.Y(n_9330)
);

AND2x4_ASAP7_75t_L g9331 ( 
.A(n_9167),
.B(n_5673),
.Y(n_9331)
);

OAI31xp33_ASAP7_75t_SL g9332 ( 
.A1(n_9162),
.A2(n_5564),
.A3(n_5841),
.B(n_5824),
.Y(n_9332)
);

OAI22xp5_ASAP7_75t_L g9333 ( 
.A1(n_9171),
.A2(n_9185),
.B1(n_9182),
.B2(n_9156),
.Y(n_9333)
);

OAI22xp33_ASAP7_75t_L g9334 ( 
.A1(n_9112),
.A2(n_5912),
.B1(n_5913),
.B2(n_5903),
.Y(n_9334)
);

NAND2xp5_ASAP7_75t_L g9335 ( 
.A(n_9172),
.B(n_5740),
.Y(n_9335)
);

NAND2xp5_ASAP7_75t_L g9336 ( 
.A(n_9175),
.B(n_5740),
.Y(n_9336)
);

NOR3xp33_ASAP7_75t_SL g9337 ( 
.A(n_9107),
.B(n_4639),
.C(n_4540),
.Y(n_9337)
);

NAND2xp5_ASAP7_75t_SL g9338 ( 
.A(n_9136),
.B(n_5673),
.Y(n_9338)
);

INVx1_ASAP7_75t_L g9339 ( 
.A(n_9111),
.Y(n_9339)
);

NAND2xp5_ASAP7_75t_L g9340 ( 
.A(n_9076),
.B(n_9115),
.Y(n_9340)
);

NAND2x1p5_ASAP7_75t_L g9341 ( 
.A(n_9155),
.B(n_3755),
.Y(n_9341)
);

AND2x2_ASAP7_75t_L g9342 ( 
.A(n_9097),
.B(n_5948),
.Y(n_9342)
);

INVx1_ASAP7_75t_L g9343 ( 
.A(n_9117),
.Y(n_9343)
);

NOR2xp33_ASAP7_75t_L g9344 ( 
.A(n_9124),
.B(n_5948),
.Y(n_9344)
);

NAND2xp5_ASAP7_75t_L g9345 ( 
.A(n_9129),
.B(n_5742),
.Y(n_9345)
);

INVx1_ASAP7_75t_L g9346 ( 
.A(n_9130),
.Y(n_9346)
);

AOI221xp5_ASAP7_75t_L g9347 ( 
.A1(n_9132),
.A2(n_5691),
.B1(n_5692),
.B2(n_5688),
.C(n_5680),
.Y(n_9347)
);

OAI21xp5_ASAP7_75t_SL g9348 ( 
.A1(n_9184),
.A2(n_4268),
.B(n_4366),
.Y(n_9348)
);

INVx1_ASAP7_75t_L g9349 ( 
.A(n_9147),
.Y(n_9349)
);

INVx1_ASAP7_75t_L g9350 ( 
.A(n_9148),
.Y(n_9350)
);

INVx1_ASAP7_75t_L g9351 ( 
.A(n_9157),
.Y(n_9351)
);

AOI21xp5_ASAP7_75t_L g9352 ( 
.A1(n_9088),
.A2(n_9077),
.B(n_9158),
.Y(n_9352)
);

AOI21xp5_ASAP7_75t_L g9353 ( 
.A1(n_9087),
.A2(n_5688),
.B(n_5680),
.Y(n_9353)
);

AOI21xp5_ASAP7_75t_L g9354 ( 
.A1(n_9069),
.A2(n_5688),
.B(n_5680),
.Y(n_9354)
);

INVx1_ASAP7_75t_L g9355 ( 
.A(n_9038),
.Y(n_9355)
);

NAND2xp5_ASAP7_75t_L g9356 ( 
.A(n_9170),
.B(n_9168),
.Y(n_9356)
);

O2A1O1Ixp33_ASAP7_75t_L g9357 ( 
.A1(n_9028),
.A2(n_6342),
.B(n_6345),
.C(n_6341),
.Y(n_9357)
);

INVx1_ASAP7_75t_SL g9358 ( 
.A(n_9032),
.Y(n_9358)
);

OAI22xp33_ASAP7_75t_L g9359 ( 
.A1(n_9034),
.A2(n_5919),
.B1(n_5932),
.B2(n_5903),
.Y(n_9359)
);

NOR4xp25_ASAP7_75t_L g9360 ( 
.A(n_9177),
.B(n_9125),
.C(n_9070),
.D(n_9110),
.Y(n_9360)
);

AOI21xp33_ASAP7_75t_L g9361 ( 
.A1(n_9073),
.A2(n_6342),
.B(n_6341),
.Y(n_9361)
);

INVx2_ASAP7_75t_SL g9362 ( 
.A(n_9139),
.Y(n_9362)
);

AO22x1_ASAP7_75t_L g9363 ( 
.A1(n_9139),
.A2(n_5692),
.B1(n_5697),
.B2(n_5691),
.Y(n_9363)
);

AND2x2_ASAP7_75t_L g9364 ( 
.A(n_9151),
.B(n_5950),
.Y(n_9364)
);

NOR4xp25_ASAP7_75t_L g9365 ( 
.A(n_9176),
.B(n_5692),
.C(n_5697),
.D(n_5691),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_9065),
.Y(n_9366)
);

OAI221xp5_ASAP7_75t_L g9367 ( 
.A1(n_9186),
.A2(n_3754),
.B1(n_4367),
.B2(n_4366),
.C(n_6341),
.Y(n_9367)
);

OAI322xp33_ASAP7_75t_L g9368 ( 
.A1(n_9173),
.A2(n_5701),
.A3(n_5709),
.B1(n_5713),
.B2(n_5712),
.C1(n_5697),
.C2(n_5919),
.Y(n_9368)
);

INVx1_ASAP7_75t_L g9369 ( 
.A(n_9189),
.Y(n_9369)
);

NOR2xp33_ASAP7_75t_L g9370 ( 
.A(n_9192),
.B(n_5950),
.Y(n_9370)
);

NOR2xp33_ASAP7_75t_L g9371 ( 
.A(n_9154),
.B(n_5958),
.Y(n_9371)
);

NAND3xp33_ASAP7_75t_SL g9372 ( 
.A(n_9134),
.B(n_4675),
.C(n_4517),
.Y(n_9372)
);

INVx1_ASAP7_75t_L g9373 ( 
.A(n_9134),
.Y(n_9373)
);

AND2x2_ASAP7_75t_L g9374 ( 
.A(n_9033),
.B(n_5958),
.Y(n_9374)
);

INVx2_ASAP7_75t_L g9375 ( 
.A(n_9212),
.Y(n_9375)
);

INVx1_ASAP7_75t_SL g9376 ( 
.A(n_9213),
.Y(n_9376)
);

NOR2x1_ASAP7_75t_L g9377 ( 
.A(n_9195),
.B(n_9284),
.Y(n_9377)
);

OAI21xp5_ASAP7_75t_L g9378 ( 
.A1(n_9231),
.A2(n_5824),
.B(n_5800),
.Y(n_9378)
);

AOI21xp33_ASAP7_75t_L g9379 ( 
.A1(n_9276),
.A2(n_6210),
.B(n_6204),
.Y(n_9379)
);

AND2x2_ASAP7_75t_L g9380 ( 
.A(n_9194),
.B(n_5963),
.Y(n_9380)
);

OR2x6_ASAP7_75t_L g9381 ( 
.A(n_9217),
.B(n_3754),
.Y(n_9381)
);

AOI22xp33_ASAP7_75t_L g9382 ( 
.A1(n_9261),
.A2(n_3738),
.B1(n_6210),
.B2(n_6204),
.Y(n_9382)
);

AOI21xp5_ASAP7_75t_L g9383 ( 
.A1(n_9232),
.A2(n_6210),
.B(n_6204),
.Y(n_9383)
);

NAND2xp5_ASAP7_75t_L g9384 ( 
.A(n_9210),
.B(n_5963),
.Y(n_9384)
);

INVx2_ASAP7_75t_L g9385 ( 
.A(n_9297),
.Y(n_9385)
);

AOI22xp5_ASAP7_75t_L g9386 ( 
.A1(n_9239),
.A2(n_5701),
.B1(n_5712),
.B2(n_5709),
.Y(n_9386)
);

AOI322xp5_ASAP7_75t_L g9387 ( 
.A1(n_9271),
.A2(n_5932),
.A3(n_5939),
.B1(n_5942),
.B2(n_5940),
.C1(n_5935),
.C2(n_5713),
.Y(n_9387)
);

OR2x2_ASAP7_75t_L g9388 ( 
.A(n_9199),
.B(n_5701),
.Y(n_9388)
);

BUFx3_ASAP7_75t_L g9389 ( 
.A(n_9218),
.Y(n_9389)
);

NAND2xp33_ASAP7_75t_SL g9390 ( 
.A(n_9220),
.B(n_3738),
.Y(n_9390)
);

INVx1_ASAP7_75t_L g9391 ( 
.A(n_9284),
.Y(n_9391)
);

INVx1_ASAP7_75t_SL g9392 ( 
.A(n_9205),
.Y(n_9392)
);

NAND2xp5_ASAP7_75t_L g9393 ( 
.A(n_9223),
.B(n_5974),
.Y(n_9393)
);

AOI21xp33_ASAP7_75t_SL g9394 ( 
.A1(n_9362),
.A2(n_6345),
.B(n_6342),
.Y(n_9394)
);

OAI22xp5_ASAP7_75t_L g9395 ( 
.A1(n_9198),
.A2(n_5712),
.B1(n_5713),
.B2(n_5709),
.Y(n_9395)
);

NAND2xp5_ASAP7_75t_L g9396 ( 
.A(n_9228),
.B(n_5974),
.Y(n_9396)
);

AOI222xp33_ASAP7_75t_L g9397 ( 
.A1(n_9305),
.A2(n_5940),
.B1(n_5935),
.B2(n_5942),
.C1(n_5939),
.C2(n_5932),
.Y(n_9397)
);

INVxp67_ASAP7_75t_SL g9398 ( 
.A(n_9297),
.Y(n_9398)
);

INVxp67_ASAP7_75t_L g9399 ( 
.A(n_9283),
.Y(n_9399)
);

OAI221xp5_ASAP7_75t_SL g9400 ( 
.A1(n_9227),
.A2(n_4426),
.B1(n_4517),
.B2(n_4875),
.C(n_4853),
.Y(n_9400)
);

NAND2xp5_ASAP7_75t_L g9401 ( 
.A(n_9234),
.B(n_5976),
.Y(n_9401)
);

OAI22xp33_ASAP7_75t_L g9402 ( 
.A1(n_9236),
.A2(n_5939),
.B1(n_5940),
.B2(n_5935),
.Y(n_9402)
);

NAND2xp5_ASAP7_75t_L g9403 ( 
.A(n_9282),
.B(n_9221),
.Y(n_9403)
);

O2A1O1Ixp33_ASAP7_75t_L g9404 ( 
.A1(n_9238),
.A2(n_6345),
.B(n_6248),
.C(n_6215),
.Y(n_9404)
);

NAND2xp5_ASAP7_75t_L g9405 ( 
.A(n_9224),
.B(n_5976),
.Y(n_9405)
);

NOR2xp33_ASAP7_75t_SL g9406 ( 
.A(n_9206),
.B(n_4231),
.Y(n_9406)
);

A2O1A1Ixp33_ASAP7_75t_L g9407 ( 
.A1(n_9201),
.A2(n_5741),
.B(n_5743),
.C(n_5571),
.Y(n_9407)
);

OAI22xp5_ASAP7_75t_L g9408 ( 
.A1(n_9229),
.A2(n_9219),
.B1(n_9230),
.B2(n_9320),
.Y(n_9408)
);

OR2x2_ASAP7_75t_L g9409 ( 
.A(n_9280),
.B(n_5742),
.Y(n_9409)
);

OAI22xp5_ASAP7_75t_L g9410 ( 
.A1(n_9248),
.A2(n_5982),
.B1(n_6000),
.B2(n_5981),
.Y(n_9410)
);

INVx1_ASAP7_75t_L g9411 ( 
.A(n_9316),
.Y(n_9411)
);

INVx1_ASAP7_75t_SL g9412 ( 
.A(n_9233),
.Y(n_9412)
);

AND2x2_ASAP7_75t_L g9413 ( 
.A(n_9202),
.B(n_5981),
.Y(n_9413)
);

OAI22xp33_ASAP7_75t_L g9414 ( 
.A1(n_9267),
.A2(n_5266),
.B1(n_5298),
.B2(n_5255),
.Y(n_9414)
);

NAND3xp33_ASAP7_75t_SL g9415 ( 
.A(n_9358),
.B(n_4675),
.C(n_4367),
.Y(n_9415)
);

OAI21xp5_ASAP7_75t_L g9416 ( 
.A1(n_9262),
.A2(n_5841),
.B(n_5800),
.Y(n_9416)
);

AOI21xp33_ASAP7_75t_L g9417 ( 
.A1(n_9311),
.A2(n_6220),
.B(n_6215),
.Y(n_9417)
);

AOI22xp5_ASAP7_75t_L g9418 ( 
.A1(n_9275),
.A2(n_5069),
.B1(n_4875),
.B2(n_4898),
.Y(n_9418)
);

AOI221x1_ASAP7_75t_L g9419 ( 
.A1(n_9352),
.A2(n_5756),
.B1(n_5766),
.B2(n_5755),
.C(n_5745),
.Y(n_9419)
);

INVx2_ASAP7_75t_SL g9420 ( 
.A(n_9341),
.Y(n_9420)
);

AOI211xp5_ASAP7_75t_L g9421 ( 
.A1(n_9203),
.A2(n_6054),
.B(n_6075),
.C(n_4626),
.Y(n_9421)
);

INVx1_ASAP7_75t_L g9422 ( 
.A(n_9316),
.Y(n_9422)
);

OAI22xp33_ASAP7_75t_SL g9423 ( 
.A1(n_9226),
.A2(n_5755),
.B1(n_5756),
.B2(n_5745),
.Y(n_9423)
);

INVx1_ASAP7_75t_L g9424 ( 
.A(n_9289),
.Y(n_9424)
);

AND2x2_ASAP7_75t_L g9425 ( 
.A(n_9246),
.B(n_5982),
.Y(n_9425)
);

INVx1_ASAP7_75t_L g9426 ( 
.A(n_9200),
.Y(n_9426)
);

INVx1_ASAP7_75t_L g9427 ( 
.A(n_9204),
.Y(n_9427)
);

INVx1_ASAP7_75t_L g9428 ( 
.A(n_9287),
.Y(n_9428)
);

INVxp67_ASAP7_75t_L g9429 ( 
.A(n_9242),
.Y(n_9429)
);

NAND2xp5_ASAP7_75t_L g9430 ( 
.A(n_9317),
.B(n_6000),
.Y(n_9430)
);

NOR2xp33_ASAP7_75t_L g9431 ( 
.A(n_9268),
.B(n_6012),
.Y(n_9431)
);

INVx1_ASAP7_75t_L g9432 ( 
.A(n_9241),
.Y(n_9432)
);

AOI22xp5_ASAP7_75t_L g9433 ( 
.A1(n_9216),
.A2(n_5001),
.B1(n_5098),
.B2(n_4853),
.Y(n_9433)
);

XOR2xp5_ASAP7_75t_L g9434 ( 
.A(n_9312),
.B(n_4178),
.Y(n_9434)
);

XNOR2x2_ASAP7_75t_L g9435 ( 
.A(n_9241),
.B(n_5741),
.Y(n_9435)
);

OAI21xp5_ASAP7_75t_L g9436 ( 
.A1(n_9196),
.A2(n_6075),
.B(n_6054),
.Y(n_9436)
);

OA21x2_ASAP7_75t_L g9437 ( 
.A1(n_9366),
.A2(n_6016),
.B(n_6012),
.Y(n_9437)
);

INVx1_ASAP7_75t_L g9438 ( 
.A(n_9264),
.Y(n_9438)
);

OAI211xp5_ASAP7_75t_L g9439 ( 
.A1(n_9274),
.A2(n_6215),
.B(n_6220),
.C(n_6248),
.Y(n_9439)
);

NAND2xp5_ASAP7_75t_L g9440 ( 
.A(n_9303),
.B(n_6016),
.Y(n_9440)
);

INVx2_ASAP7_75t_L g9441 ( 
.A(n_9327),
.Y(n_9441)
);

AO21x1_ASAP7_75t_L g9442 ( 
.A1(n_9245),
.A2(n_6038),
.B(n_6020),
.Y(n_9442)
);

OAI321xp33_ASAP7_75t_L g9443 ( 
.A1(n_9207),
.A2(n_4675),
.A3(n_4366),
.B1(n_4573),
.B2(n_4572),
.C(n_4525),
.Y(n_9443)
);

INVx1_ASAP7_75t_L g9444 ( 
.A(n_9374),
.Y(n_9444)
);

AND2x2_ASAP7_75t_L g9445 ( 
.A(n_9209),
.B(n_6020),
.Y(n_9445)
);

OAI22xp33_ASAP7_75t_L g9446 ( 
.A1(n_9222),
.A2(n_5266),
.B1(n_5298),
.B2(n_5255),
.Y(n_9446)
);

AOI22xp33_ASAP7_75t_L g9447 ( 
.A1(n_9235),
.A2(n_6220),
.B1(n_3760),
.B2(n_3755),
.Y(n_9447)
);

INVx1_ASAP7_75t_SL g9448 ( 
.A(n_9315),
.Y(n_9448)
);

INVx1_ASAP7_75t_L g9449 ( 
.A(n_9356),
.Y(n_9449)
);

OAI21xp33_ASAP7_75t_SL g9450 ( 
.A1(n_9277),
.A2(n_5743),
.B(n_5603),
.Y(n_9450)
);

NAND2xp5_ASAP7_75t_L g9451 ( 
.A(n_9250),
.B(n_6038),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_9298),
.Y(n_9452)
);

NAND2xp5_ASAP7_75t_L g9453 ( 
.A(n_9360),
.B(n_6039),
.Y(n_9453)
);

AND2x2_ASAP7_75t_L g9454 ( 
.A(n_9215),
.B(n_6039),
.Y(n_9454)
);

NAND2xp5_ASAP7_75t_L g9455 ( 
.A(n_9285),
.B(n_6049),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_9340),
.Y(n_9456)
);

AND2x2_ASAP7_75t_L g9457 ( 
.A(n_9279),
.B(n_6049),
.Y(n_9457)
);

AOI221xp5_ASAP7_75t_L g9458 ( 
.A1(n_9211),
.A2(n_5771),
.B1(n_5773),
.B2(n_5768),
.C(n_5766),
.Y(n_9458)
);

INVx2_ASAP7_75t_SL g9459 ( 
.A(n_9288),
.Y(n_9459)
);

AOI221xp5_ASAP7_75t_L g9460 ( 
.A1(n_9333),
.A2(n_5773),
.B1(n_5780),
.B2(n_5771),
.C(n_5768),
.Y(n_9460)
);

AND2x2_ASAP7_75t_L g9461 ( 
.A(n_9319),
.B(n_6052),
.Y(n_9461)
);

INVxp67_ASAP7_75t_L g9462 ( 
.A(n_9225),
.Y(n_9462)
);

INVx1_ASAP7_75t_L g9463 ( 
.A(n_9260),
.Y(n_9463)
);

NAND2xp5_ASAP7_75t_L g9464 ( 
.A(n_9197),
.B(n_6052),
.Y(n_9464)
);

INVx1_ASAP7_75t_L g9465 ( 
.A(n_9272),
.Y(n_9465)
);

OAI31xp33_ASAP7_75t_L g9466 ( 
.A1(n_9373),
.A2(n_4573),
.A3(n_4572),
.B(n_3848),
.Y(n_9466)
);

OAI22xp5_ASAP7_75t_L g9467 ( 
.A1(n_9293),
.A2(n_9326),
.B1(n_9301),
.B2(n_9337),
.Y(n_9467)
);

NAND2xp5_ASAP7_75t_SL g9468 ( 
.A(n_9307),
.B(n_4853),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_SL g9469 ( 
.A(n_9214),
.B(n_4898),
.Y(n_9469)
);

AOI21xp5_ASAP7_75t_L g9470 ( 
.A1(n_9278),
.A2(n_9263),
.B(n_9253),
.Y(n_9470)
);

OR2x2_ASAP7_75t_L g9471 ( 
.A(n_9255),
.B(n_5780),
.Y(n_9471)
);

OAI221xp5_ASAP7_75t_L g9472 ( 
.A1(n_9291),
.A2(n_3760),
.B1(n_3755),
.B2(n_4995),
.C(n_4910),
.Y(n_9472)
);

NAND2xp5_ASAP7_75t_L g9473 ( 
.A(n_9252),
.B(n_6070),
.Y(n_9473)
);

INVx2_ASAP7_75t_L g9474 ( 
.A(n_9328),
.Y(n_9474)
);

NAND2x1_ASAP7_75t_L g9475 ( 
.A(n_9331),
.B(n_6070),
.Y(n_9475)
);

INVx2_ASAP7_75t_L g9476 ( 
.A(n_9321),
.Y(n_9476)
);

AOI221xp5_ASAP7_75t_L g9477 ( 
.A1(n_9208),
.A2(n_5804),
.B1(n_5805),
.B2(n_5783),
.C(n_5782),
.Y(n_9477)
);

OAI322xp33_ASAP7_75t_L g9478 ( 
.A1(n_9302),
.A2(n_5804),
.A3(n_5782),
.B1(n_5807),
.B2(n_5809),
.C1(n_5805),
.C2(n_5783),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_9292),
.Y(n_9479)
);

OAI21xp33_ASAP7_75t_L g9480 ( 
.A1(n_9310),
.A2(n_4910),
.B(n_4898),
.Y(n_9480)
);

AOI21xp33_ASAP7_75t_SL g9481 ( 
.A1(n_9322),
.A2(n_9329),
.B(n_9325),
.Y(n_9481)
);

INVx1_ASAP7_75t_L g9482 ( 
.A(n_9339),
.Y(n_9482)
);

INVx1_ASAP7_75t_L g9483 ( 
.A(n_9343),
.Y(n_9483)
);

INVx1_ASAP7_75t_L g9484 ( 
.A(n_9346),
.Y(n_9484)
);

O2A1O1Ixp5_ASAP7_75t_L g9485 ( 
.A1(n_9338),
.A2(n_9269),
.B(n_9251),
.C(n_9306),
.Y(n_9485)
);

INVxp67_ASAP7_75t_L g9486 ( 
.A(n_9349),
.Y(n_9486)
);

INVx2_ASAP7_75t_L g9487 ( 
.A(n_9342),
.Y(n_9487)
);

INVx1_ASAP7_75t_L g9488 ( 
.A(n_9350),
.Y(n_9488)
);

AOI21xp5_ASAP7_75t_L g9489 ( 
.A1(n_9244),
.A2(n_6248),
.B(n_6236),
.Y(n_9489)
);

NAND2xp5_ASAP7_75t_L g9490 ( 
.A(n_9257),
.B(n_5807),
.Y(n_9490)
);

AND2x2_ASAP7_75t_L g9491 ( 
.A(n_9351),
.B(n_5809),
.Y(n_9491)
);

INVx1_ASAP7_75t_SL g9492 ( 
.A(n_9249),
.Y(n_9492)
);

INVxp67_ASAP7_75t_L g9493 ( 
.A(n_9259),
.Y(n_9493)
);

OAI22xp5_ASAP7_75t_L g9494 ( 
.A1(n_9240),
.A2(n_5816),
.B1(n_5819),
.B2(n_5811),
.Y(n_9494)
);

AOI221xp5_ASAP7_75t_L g9495 ( 
.A1(n_9370),
.A2(n_5819),
.B1(n_5821),
.B2(n_5816),
.C(n_5811),
.Y(n_9495)
);

INVx1_ASAP7_75t_L g9496 ( 
.A(n_9270),
.Y(n_9496)
);

AND2x2_ASAP7_75t_L g9497 ( 
.A(n_9299),
.B(n_5821),
.Y(n_9497)
);

NAND2xp5_ASAP7_75t_L g9498 ( 
.A(n_9355),
.B(n_9369),
.Y(n_9498)
);

NAND2xp5_ASAP7_75t_L g9499 ( 
.A(n_9344),
.B(n_5822),
.Y(n_9499)
);

INVx2_ASAP7_75t_L g9500 ( 
.A(n_9286),
.Y(n_9500)
);

NAND2xp33_ASAP7_75t_L g9501 ( 
.A(n_9295),
.B(n_5822),
.Y(n_9501)
);

INVx1_ASAP7_75t_L g9502 ( 
.A(n_9335),
.Y(n_9502)
);

INVx1_ASAP7_75t_L g9503 ( 
.A(n_9336),
.Y(n_9503)
);

OAI22xp5_ASAP7_75t_L g9504 ( 
.A1(n_9247),
.A2(n_5829),
.B1(n_5832),
.B2(n_5825),
.Y(n_9504)
);

AOI21xp5_ASAP7_75t_SL g9505 ( 
.A1(n_9331),
.A2(n_3760),
.B(n_4178),
.Y(n_9505)
);

XOR2x2_ASAP7_75t_L g9506 ( 
.A(n_9345),
.B(n_4629),
.Y(n_9506)
);

OAI22xp5_ASAP7_75t_L g9507 ( 
.A1(n_9348),
.A2(n_5829),
.B1(n_5832),
.B2(n_5825),
.Y(n_9507)
);

OAI31xp33_ASAP7_75t_L g9508 ( 
.A1(n_9281),
.A2(n_4573),
.A3(n_4572),
.B(n_3848),
.Y(n_9508)
);

O2A1O1Ixp33_ASAP7_75t_L g9509 ( 
.A1(n_9273),
.A2(n_9254),
.B(n_9372),
.C(n_9323),
.Y(n_9509)
);

INVx1_ASAP7_75t_L g9510 ( 
.A(n_9330),
.Y(n_9510)
);

AND2x2_ASAP7_75t_L g9511 ( 
.A(n_9364),
.B(n_5844),
.Y(n_9511)
);

AOI222xp33_ASAP7_75t_L g9512 ( 
.A1(n_9371),
.A2(n_5854),
.B1(n_5844),
.B2(n_5861),
.C1(n_5859),
.C2(n_5848),
.Y(n_9512)
);

INVx1_ASAP7_75t_SL g9513 ( 
.A(n_9318),
.Y(n_9513)
);

AND2x2_ASAP7_75t_L g9514 ( 
.A(n_9237),
.B(n_5848),
.Y(n_9514)
);

AOI22xp5_ASAP7_75t_L g9515 ( 
.A1(n_9290),
.A2(n_9258),
.B1(n_9304),
.B2(n_9266),
.Y(n_9515)
);

INVx1_ASAP7_75t_L g9516 ( 
.A(n_9363),
.Y(n_9516)
);

NAND2xp5_ASAP7_75t_L g9517 ( 
.A(n_9309),
.B(n_9300),
.Y(n_9517)
);

INVx1_ASAP7_75t_L g9518 ( 
.A(n_9294),
.Y(n_9518)
);

NAND3x2_ASAP7_75t_L g9519 ( 
.A(n_9332),
.B(n_4225),
.C(n_4220),
.Y(n_9519)
);

AOI221xp5_ASAP7_75t_L g9520 ( 
.A1(n_9365),
.A2(n_5861),
.B1(n_5863),
.B2(n_5859),
.C(n_5854),
.Y(n_9520)
);

AOI21xp33_ASAP7_75t_SL g9521 ( 
.A1(n_9256),
.A2(n_9367),
.B(n_9265),
.Y(n_9521)
);

AOI22x1_ASAP7_75t_L g9522 ( 
.A1(n_9296),
.A2(n_5865),
.B1(n_5869),
.B2(n_5863),
.Y(n_9522)
);

INVx1_ASAP7_75t_L g9523 ( 
.A(n_9313),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_9398),
.Y(n_9524)
);

NAND2xp5_ASAP7_75t_L g9525 ( 
.A(n_9432),
.B(n_9354),
.Y(n_9525)
);

NAND2xp5_ASAP7_75t_SL g9526 ( 
.A(n_9385),
.B(n_9308),
.Y(n_9526)
);

INVx1_ASAP7_75t_L g9527 ( 
.A(n_9377),
.Y(n_9527)
);

INVx1_ASAP7_75t_L g9528 ( 
.A(n_9377),
.Y(n_9528)
);

NAND2xp5_ASAP7_75t_L g9529 ( 
.A(n_9376),
.B(n_9353),
.Y(n_9529)
);

AND2x2_ASAP7_75t_L g9530 ( 
.A(n_9375),
.B(n_9314),
.Y(n_9530)
);

NAND2xp5_ASAP7_75t_L g9531 ( 
.A(n_9411),
.B(n_9243),
.Y(n_9531)
);

NAND2xp5_ASAP7_75t_L g9532 ( 
.A(n_9422),
.B(n_9334),
.Y(n_9532)
);

NAND2xp5_ASAP7_75t_SL g9533 ( 
.A(n_9423),
.B(n_9386),
.Y(n_9533)
);

NAND2xp5_ASAP7_75t_L g9534 ( 
.A(n_9429),
.B(n_9424),
.Y(n_9534)
);

NAND3xp33_ASAP7_75t_L g9535 ( 
.A(n_9391),
.B(n_9361),
.C(n_9357),
.Y(n_9535)
);

INVx1_ASAP7_75t_L g9536 ( 
.A(n_9403),
.Y(n_9536)
);

NAND2xp5_ASAP7_75t_L g9537 ( 
.A(n_9412),
.B(n_9392),
.Y(n_9537)
);

AND2x2_ASAP7_75t_L g9538 ( 
.A(n_9441),
.B(n_9347),
.Y(n_9538)
);

INVx2_ASAP7_75t_L g9539 ( 
.A(n_9389),
.Y(n_9539)
);

NAND2xp5_ASAP7_75t_L g9540 ( 
.A(n_9428),
.B(n_9359),
.Y(n_9540)
);

INVx1_ASAP7_75t_L g9541 ( 
.A(n_9459),
.Y(n_9541)
);

INVxp67_ASAP7_75t_L g9542 ( 
.A(n_9406),
.Y(n_9542)
);

INVxp33_ASAP7_75t_SL g9543 ( 
.A(n_9408),
.Y(n_9543)
);

NAND2xp5_ASAP7_75t_L g9544 ( 
.A(n_9420),
.B(n_9324),
.Y(n_9544)
);

NAND2xp5_ASAP7_75t_L g9545 ( 
.A(n_9448),
.B(n_5865),
.Y(n_9545)
);

NAND2xp5_ASAP7_75t_L g9546 ( 
.A(n_9444),
.B(n_5869),
.Y(n_9546)
);

AOI222xp33_ASAP7_75t_L g9547 ( 
.A1(n_9469),
.A2(n_9368),
.B1(n_5879),
.B2(n_5871),
.C1(n_5882),
.C2(n_5881),
.Y(n_9547)
);

OR2x2_ASAP7_75t_L g9548 ( 
.A(n_9476),
.B(n_6236),
.Y(n_9548)
);

INVx1_ASAP7_75t_SL g9549 ( 
.A(n_9492),
.Y(n_9549)
);

NOR2x1p5_ASAP7_75t_SL g9550 ( 
.A(n_9516),
.B(n_5871),
.Y(n_9550)
);

NAND2xp5_ASAP7_75t_L g9551 ( 
.A(n_9487),
.B(n_5876),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9435),
.Y(n_9552)
);

INVx1_ASAP7_75t_SL g9553 ( 
.A(n_9380),
.Y(n_9553)
);

INVx1_ASAP7_75t_L g9554 ( 
.A(n_9453),
.Y(n_9554)
);

NAND2xp5_ASAP7_75t_L g9555 ( 
.A(n_9426),
.B(n_5876),
.Y(n_9555)
);

INVx1_ASAP7_75t_L g9556 ( 
.A(n_9506),
.Y(n_9556)
);

AOI22xp33_ASAP7_75t_L g9557 ( 
.A1(n_9438),
.A2(n_5746),
.B1(n_5477),
.B2(n_5849),
.Y(n_9557)
);

INVx1_ASAP7_75t_L g9558 ( 
.A(n_9427),
.Y(n_9558)
);

AND2x2_ASAP7_75t_L g9559 ( 
.A(n_9462),
.B(n_5879),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_9452),
.Y(n_9560)
);

OR2x2_ASAP7_75t_L g9561 ( 
.A(n_9474),
.B(n_6236),
.Y(n_9561)
);

INVx1_ASAP7_75t_L g9562 ( 
.A(n_9405),
.Y(n_9562)
);

NAND2xp5_ASAP7_75t_L g9563 ( 
.A(n_9470),
.B(n_5881),
.Y(n_9563)
);

INVx1_ASAP7_75t_L g9564 ( 
.A(n_9409),
.Y(n_9564)
);

INVx1_ASAP7_75t_L g9565 ( 
.A(n_9425),
.Y(n_9565)
);

AOI22xp33_ASAP7_75t_SL g9566 ( 
.A1(n_9519),
.A2(n_4995),
.B1(n_5021),
.B2(n_5001),
.Y(n_9566)
);

NAND2xp5_ASAP7_75t_L g9567 ( 
.A(n_9465),
.B(n_5882),
.Y(n_9567)
);

INVx1_ASAP7_75t_L g9568 ( 
.A(n_9479),
.Y(n_9568)
);

INVx1_ASAP7_75t_L g9569 ( 
.A(n_9482),
.Y(n_9569)
);

INVx2_ASAP7_75t_L g9570 ( 
.A(n_9434),
.Y(n_9570)
);

INVx1_ASAP7_75t_L g9571 ( 
.A(n_9483),
.Y(n_9571)
);

HB1xp67_ASAP7_75t_L g9572 ( 
.A(n_9381),
.Y(n_9572)
);

INVx1_ASAP7_75t_L g9573 ( 
.A(n_9484),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_9488),
.Y(n_9574)
);

INVx2_ASAP7_75t_L g9575 ( 
.A(n_9381),
.Y(n_9575)
);

NAND2xp5_ASAP7_75t_L g9576 ( 
.A(n_9500),
.B(n_5893),
.Y(n_9576)
);

NAND2xp5_ASAP7_75t_L g9577 ( 
.A(n_9481),
.B(n_9413),
.Y(n_9577)
);

AND2x2_ASAP7_75t_L g9578 ( 
.A(n_9449),
.B(n_5893),
.Y(n_9578)
);

INVx1_ASAP7_75t_SL g9579 ( 
.A(n_9390),
.Y(n_9579)
);

INVx1_ASAP7_75t_L g9580 ( 
.A(n_9464),
.Y(n_9580)
);

INVx1_ASAP7_75t_SL g9581 ( 
.A(n_9457),
.Y(n_9581)
);

AND2x2_ASAP7_75t_L g9582 ( 
.A(n_9456),
.B(n_5898),
.Y(n_9582)
);

NOR2xp33_ASAP7_75t_L g9583 ( 
.A(n_9486),
.B(n_5898),
.Y(n_9583)
);

AND2x2_ASAP7_75t_L g9584 ( 
.A(n_9399),
.B(n_5899),
.Y(n_9584)
);

AOI21xp33_ASAP7_75t_L g9585 ( 
.A1(n_9509),
.A2(n_6240),
.B(n_5477),
.Y(n_9585)
);

NOR2xp33_ASAP7_75t_L g9586 ( 
.A(n_9493),
.B(n_5899),
.Y(n_9586)
);

NOR2xp33_ASAP7_75t_L g9587 ( 
.A(n_9513),
.B(n_5906),
.Y(n_9587)
);

NAND2xp5_ASAP7_75t_L g9588 ( 
.A(n_9445),
.B(n_5906),
.Y(n_9588)
);

NAND2xp5_ASAP7_75t_SL g9589 ( 
.A(n_9446),
.B(n_5907),
.Y(n_9589)
);

INVx1_ASAP7_75t_L g9590 ( 
.A(n_9396),
.Y(n_9590)
);

INVx2_ASAP7_75t_L g9591 ( 
.A(n_9522),
.Y(n_9591)
);

NAND2xp5_ASAP7_75t_L g9592 ( 
.A(n_9454),
.B(n_5907),
.Y(n_9592)
);

HB1xp67_ASAP7_75t_L g9593 ( 
.A(n_9437),
.Y(n_9593)
);

INVx1_ASAP7_75t_L g9594 ( 
.A(n_9401),
.Y(n_9594)
);

INVx1_ASAP7_75t_L g9595 ( 
.A(n_9491),
.Y(n_9595)
);

NAND2xp5_ASAP7_75t_SL g9596 ( 
.A(n_9404),
.B(n_5925),
.Y(n_9596)
);

OR2x2_ASAP7_75t_L g9597 ( 
.A(n_9430),
.B(n_6240),
.Y(n_9597)
);

CKINVDCx16_ASAP7_75t_R g9598 ( 
.A(n_9518),
.Y(n_9598)
);

NAND2xp5_ASAP7_75t_L g9599 ( 
.A(n_9461),
.B(n_5925),
.Y(n_9599)
);

NAND2xp5_ASAP7_75t_SL g9600 ( 
.A(n_9402),
.B(n_9458),
.Y(n_9600)
);

OR2x6_ASAP7_75t_L g9601 ( 
.A(n_9498),
.B(n_9463),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_9471),
.Y(n_9602)
);

INVx1_ASAP7_75t_L g9603 ( 
.A(n_9384),
.Y(n_9603)
);

NAND2xp5_ASAP7_75t_L g9604 ( 
.A(n_9431),
.B(n_5927),
.Y(n_9604)
);

NAND2xp5_ASAP7_75t_L g9605 ( 
.A(n_9523),
.B(n_5927),
.Y(n_9605)
);

AND2x2_ASAP7_75t_L g9606 ( 
.A(n_9510),
.B(n_5930),
.Y(n_9606)
);

AND2x2_ASAP7_75t_L g9607 ( 
.A(n_9496),
.B(n_5930),
.Y(n_9607)
);

NAND2xp5_ASAP7_75t_L g9608 ( 
.A(n_9502),
.B(n_5931),
.Y(n_9608)
);

INVx1_ASAP7_75t_L g9609 ( 
.A(n_9440),
.Y(n_9609)
);

BUFx2_ASAP7_75t_SL g9610 ( 
.A(n_9503),
.Y(n_9610)
);

INVx1_ASAP7_75t_SL g9611 ( 
.A(n_9388),
.Y(n_9611)
);

AND2x4_ASAP7_75t_L g9612 ( 
.A(n_9517),
.B(n_5931),
.Y(n_9612)
);

NOR2xp33_ASAP7_75t_L g9613 ( 
.A(n_9393),
.B(n_9467),
.Y(n_9613)
);

INVx1_ASAP7_75t_L g9614 ( 
.A(n_9485),
.Y(n_9614)
);

INVx1_ASAP7_75t_SL g9615 ( 
.A(n_9451),
.Y(n_9615)
);

INVx1_ASAP7_75t_SL g9616 ( 
.A(n_9455),
.Y(n_9616)
);

HB1xp67_ASAP7_75t_L g9617 ( 
.A(n_9437),
.Y(n_9617)
);

NAND2xp5_ASAP7_75t_L g9618 ( 
.A(n_9497),
.B(n_9515),
.Y(n_9618)
);

INVx1_ASAP7_75t_L g9619 ( 
.A(n_9501),
.Y(n_9619)
);

NAND2x1p5_ASAP7_75t_L g9620 ( 
.A(n_9475),
.B(n_4231),
.Y(n_9620)
);

AND2x2_ASAP7_75t_L g9621 ( 
.A(n_9505),
.B(n_5937),
.Y(n_9621)
);

AND2x2_ASAP7_75t_L g9622 ( 
.A(n_9511),
.B(n_9521),
.Y(n_9622)
);

OAI221xp5_ASAP7_75t_L g9623 ( 
.A1(n_9460),
.A2(n_6240),
.B1(n_3848),
.B2(n_3846),
.C(n_5001),
.Y(n_9623)
);

OR2x2_ASAP7_75t_L g9624 ( 
.A(n_9473),
.B(n_5967),
.Y(n_9624)
);

NAND2xp5_ASAP7_75t_L g9625 ( 
.A(n_9490),
.B(n_5937),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_9499),
.Y(n_9626)
);

NAND2xp5_ASAP7_75t_L g9627 ( 
.A(n_9419),
.B(n_5949),
.Y(n_9627)
);

NOR2x1_ASAP7_75t_L g9628 ( 
.A(n_9514),
.B(n_5949),
.Y(n_9628)
);

INVx1_ASAP7_75t_L g9629 ( 
.A(n_9442),
.Y(n_9629)
);

INVx1_ASAP7_75t_L g9630 ( 
.A(n_9504),
.Y(n_9630)
);

AOI22xp33_ASAP7_75t_L g9631 ( 
.A1(n_9415),
.A2(n_5746),
.B1(n_5477),
.B2(n_5849),
.Y(n_9631)
);

AND2x2_ASAP7_75t_L g9632 ( 
.A(n_9433),
.B(n_5952),
.Y(n_9632)
);

NAND2xp5_ASAP7_75t_L g9633 ( 
.A(n_9414),
.B(n_5952),
.Y(n_9633)
);

INVx1_ASAP7_75t_L g9634 ( 
.A(n_9494),
.Y(n_9634)
);

INVxp67_ASAP7_75t_L g9635 ( 
.A(n_9472),
.Y(n_9635)
);

INVx1_ASAP7_75t_SL g9636 ( 
.A(n_9468),
.Y(n_9636)
);

NOR2xp33_ASAP7_75t_L g9637 ( 
.A(n_9400),
.B(n_5955),
.Y(n_9637)
);

INVx1_ASAP7_75t_L g9638 ( 
.A(n_9478),
.Y(n_9638)
);

NAND2xp5_ASAP7_75t_L g9639 ( 
.A(n_9407),
.B(n_5955),
.Y(n_9639)
);

NAND2xp5_ASAP7_75t_L g9640 ( 
.A(n_9447),
.B(n_5957),
.Y(n_9640)
);

INVx1_ASAP7_75t_SL g9641 ( 
.A(n_9383),
.Y(n_9641)
);

NAND2xp5_ASAP7_75t_L g9642 ( 
.A(n_9421),
.B(n_9416),
.Y(n_9642)
);

NAND2xp5_ASAP7_75t_SL g9643 ( 
.A(n_9443),
.B(n_5957),
.Y(n_9643)
);

OR2x2_ASAP7_75t_L g9644 ( 
.A(n_9507),
.B(n_5983),
.Y(n_9644)
);

INVx1_ASAP7_75t_L g9645 ( 
.A(n_9395),
.Y(n_9645)
);

NOR3xp33_ASAP7_75t_L g9646 ( 
.A(n_9598),
.B(n_9534),
.C(n_9536),
.Y(n_9646)
);

NAND2xp5_ASAP7_75t_SL g9647 ( 
.A(n_9543),
.B(n_9379),
.Y(n_9647)
);

NAND4xp75_ASAP7_75t_L g9648 ( 
.A(n_9537),
.B(n_9436),
.C(n_9508),
.D(n_9466),
.Y(n_9648)
);

NAND3xp33_ASAP7_75t_SL g9649 ( 
.A(n_9549),
.B(n_9489),
.C(n_9382),
.Y(n_9649)
);

NOR2x1_ASAP7_75t_L g9650 ( 
.A(n_9527),
.B(n_9439),
.Y(n_9650)
);

INVx1_ASAP7_75t_L g9651 ( 
.A(n_9550),
.Y(n_9651)
);

NOR3xp33_ASAP7_75t_L g9652 ( 
.A(n_9524),
.B(n_9450),
.C(n_9417),
.Y(n_9652)
);

AOI21xp5_ASAP7_75t_L g9653 ( 
.A1(n_9577),
.A2(n_9378),
.B(n_9394),
.Y(n_9653)
);

AOI221xp5_ASAP7_75t_L g9654 ( 
.A1(n_9614),
.A2(n_9541),
.B1(n_9636),
.B2(n_9638),
.C(n_9579),
.Y(n_9654)
);

NAND2xp5_ASAP7_75t_L g9655 ( 
.A(n_9530),
.B(n_9477),
.Y(n_9655)
);

NAND2xp5_ASAP7_75t_L g9656 ( 
.A(n_9539),
.B(n_9480),
.Y(n_9656)
);

NOR2xp33_ASAP7_75t_L g9657 ( 
.A(n_9553),
.B(n_9418),
.Y(n_9657)
);

NOR3x1_ASAP7_75t_L g9658 ( 
.A(n_9544),
.B(n_9410),
.C(n_9394),
.Y(n_9658)
);

NAND2xp5_ASAP7_75t_L g9659 ( 
.A(n_9581),
.B(n_9495),
.Y(n_9659)
);

NAND2xp5_ASAP7_75t_L g9660 ( 
.A(n_9622),
.B(n_9554),
.Y(n_9660)
);

OAI211xp5_ASAP7_75t_SL g9661 ( 
.A1(n_9635),
.A2(n_9387),
.B(n_9520),
.C(n_9397),
.Y(n_9661)
);

NOR2x1_ASAP7_75t_L g9662 ( 
.A(n_9528),
.B(n_5962),
.Y(n_9662)
);

NOR2xp33_ASAP7_75t_SL g9663 ( 
.A(n_9572),
.B(n_4231),
.Y(n_9663)
);

AOI21xp33_ASAP7_75t_L g9664 ( 
.A1(n_9618),
.A2(n_9512),
.B(n_5477),
.Y(n_9664)
);

NAND5xp2_ASAP7_75t_L g9665 ( 
.A(n_9613),
.B(n_4572),
.C(n_4573),
.D(n_4525),
.E(n_4480),
.Y(n_9665)
);

OR2x2_ASAP7_75t_L g9666 ( 
.A(n_9529),
.B(n_5962),
.Y(n_9666)
);

INVx1_ASAP7_75t_L g9667 ( 
.A(n_9593),
.Y(n_9667)
);

NAND4xp25_ASAP7_75t_L g9668 ( 
.A(n_9556),
.B(n_4715),
.C(n_3846),
.D(n_4637),
.Y(n_9668)
);

NOR2xp33_ASAP7_75t_L g9669 ( 
.A(n_9526),
.B(n_5967),
.Y(n_9669)
);

INVx1_ASAP7_75t_L g9670 ( 
.A(n_9617),
.Y(n_9670)
);

INVx1_ASAP7_75t_L g9671 ( 
.A(n_9552),
.Y(n_9671)
);

INVx1_ASAP7_75t_L g9672 ( 
.A(n_9525),
.Y(n_9672)
);

NAND3xp33_ASAP7_75t_L g9673 ( 
.A(n_9535),
.B(n_5969),
.C(n_5968),
.Y(n_9673)
);

NAND2xp5_ASAP7_75t_L g9674 ( 
.A(n_9558),
.B(n_5968),
.Y(n_9674)
);

NOR3xp33_ASAP7_75t_SL g9675 ( 
.A(n_9535),
.B(n_4638),
.C(n_4635),
.Y(n_9675)
);

NOR3xp33_ASAP7_75t_L g9676 ( 
.A(n_9570),
.B(n_4715),
.C(n_4396),
.Y(n_9676)
);

NAND4xp75_ASAP7_75t_L g9677 ( 
.A(n_9538),
.B(n_9531),
.C(n_9560),
.D(n_9568),
.Y(n_9677)
);

NOR3x1_ASAP7_75t_L g9678 ( 
.A(n_9532),
.B(n_5571),
.C(n_5603),
.Y(n_9678)
);

OAI211xp5_ASAP7_75t_SL g9679 ( 
.A1(n_9542),
.A2(n_4316),
.B(n_4404),
.C(n_4396),
.Y(n_9679)
);

NAND2xp5_ASAP7_75t_L g9680 ( 
.A(n_9595),
.B(n_9569),
.Y(n_9680)
);

NAND3xp33_ASAP7_75t_SL g9681 ( 
.A(n_9641),
.B(n_9611),
.C(n_9615),
.Y(n_9681)
);

AND2x2_ASAP7_75t_L g9682 ( 
.A(n_9565),
.B(n_5969),
.Y(n_9682)
);

AOI21xp5_ASAP7_75t_L g9683 ( 
.A1(n_9601),
.A2(n_5972),
.B(n_5970),
.Y(n_9683)
);

NAND2xp5_ASAP7_75t_L g9684 ( 
.A(n_9571),
.B(n_5970),
.Y(n_9684)
);

INVx1_ASAP7_75t_L g9685 ( 
.A(n_9629),
.Y(n_9685)
);

AOI221xp5_ASAP7_75t_SL g9686 ( 
.A1(n_9533),
.A2(n_5972),
.B1(n_5989),
.B2(n_5984),
.C(n_5983),
.Y(n_9686)
);

NOR3xp33_ASAP7_75t_L g9687 ( 
.A(n_9540),
.B(n_4715),
.C(n_4404),
.Y(n_9687)
);

HB1xp67_ASAP7_75t_L g9688 ( 
.A(n_9601),
.Y(n_9688)
);

INVx2_ASAP7_75t_L g9689 ( 
.A(n_9620),
.Y(n_9689)
);

INVx1_ASAP7_75t_L g9690 ( 
.A(n_9573),
.Y(n_9690)
);

OAI22xp5_ASAP7_75t_L g9691 ( 
.A1(n_9566),
.A2(n_5989),
.B1(n_5990),
.B2(n_5984),
.Y(n_9691)
);

OAI21xp33_ASAP7_75t_L g9692 ( 
.A1(n_9642),
.A2(n_5001),
.B(n_4995),
.Y(n_9692)
);

OAI221xp5_ASAP7_75t_L g9693 ( 
.A1(n_9645),
.A2(n_5990),
.B1(n_5993),
.B2(n_5992),
.C(n_5991),
.Y(n_9693)
);

NAND2xp5_ASAP7_75t_L g9694 ( 
.A(n_9574),
.B(n_5992),
.Y(n_9694)
);

INVx1_ASAP7_75t_L g9695 ( 
.A(n_9545),
.Y(n_9695)
);

INVx1_ASAP7_75t_L g9696 ( 
.A(n_9610),
.Y(n_9696)
);

INVx1_ASAP7_75t_L g9697 ( 
.A(n_9564),
.Y(n_9697)
);

NAND2xp5_ASAP7_75t_L g9698 ( 
.A(n_9621),
.B(n_5993),
.Y(n_9698)
);

AND2x2_ASAP7_75t_L g9699 ( 
.A(n_9584),
.B(n_5991),
.Y(n_9699)
);

NOR3xp33_ASAP7_75t_L g9700 ( 
.A(n_9580),
.B(n_4715),
.C(n_4995),
.Y(n_9700)
);

INVx1_ASAP7_75t_L g9701 ( 
.A(n_9551),
.Y(n_9701)
);

INVx1_ASAP7_75t_L g9702 ( 
.A(n_9559),
.Y(n_9702)
);

AOI21xp5_ASAP7_75t_L g9703 ( 
.A1(n_9601),
.A2(n_6003),
.B(n_5997),
.Y(n_9703)
);

NAND4xp25_ASAP7_75t_L g9704 ( 
.A(n_9583),
.B(n_3846),
.C(n_4637),
.D(n_4225),
.Y(n_9704)
);

NOR2xp33_ASAP7_75t_L g9705 ( 
.A(n_9616),
.B(n_5997),
.Y(n_9705)
);

NOR3xp33_ASAP7_75t_L g9706 ( 
.A(n_9562),
.B(n_5069),
.C(n_5021),
.Y(n_9706)
);

AOI21xp5_ASAP7_75t_L g9707 ( 
.A1(n_9600),
.A2(n_9563),
.B(n_9602),
.Y(n_9707)
);

NOR3x1_ASAP7_75t_L g9708 ( 
.A(n_9630),
.B(n_5626),
.C(n_5779),
.Y(n_9708)
);

NAND4xp25_ASAP7_75t_L g9709 ( 
.A(n_9587),
.B(n_4252),
.C(n_4322),
.D(n_4220),
.Y(n_9709)
);

INVx1_ASAP7_75t_L g9710 ( 
.A(n_9576),
.Y(n_9710)
);

NOR4xp25_ASAP7_75t_L g9711 ( 
.A(n_9615),
.B(n_6004),
.C(n_6005),
.D(n_6003),
.Y(n_9711)
);

NOR3x1_ASAP7_75t_L g9712 ( 
.A(n_9634),
.B(n_5779),
.C(n_6004),
.Y(n_9712)
);

NAND3xp33_ASAP7_75t_L g9713 ( 
.A(n_9591),
.B(n_6010),
.C(n_6005),
.Y(n_9713)
);

INVx1_ASAP7_75t_L g9714 ( 
.A(n_9578),
.Y(n_9714)
);

INVx1_ASAP7_75t_L g9715 ( 
.A(n_9582),
.Y(n_9715)
);

NAND2xp5_ASAP7_75t_L g9716 ( 
.A(n_9575),
.B(n_6010),
.Y(n_9716)
);

O2A1O1Ixp5_ASAP7_75t_L g9717 ( 
.A1(n_9596),
.A2(n_6013),
.B(n_6017),
.C(n_6011),
.Y(n_9717)
);

OAI21xp5_ASAP7_75t_SL g9718 ( 
.A1(n_9637),
.A2(n_5069),
.B(n_5021),
.Y(n_9718)
);

OAI221xp5_ASAP7_75t_SL g9719 ( 
.A1(n_9605),
.A2(n_5074),
.B1(n_5021),
.B2(n_5098),
.C(n_5069),
.Y(n_9719)
);

INVx1_ASAP7_75t_L g9720 ( 
.A(n_9546),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_9555),
.Y(n_9721)
);

NAND3xp33_ASAP7_75t_L g9722 ( 
.A(n_9619),
.B(n_6013),
.C(n_6011),
.Y(n_9722)
);

NAND4xp25_ASAP7_75t_L g9723 ( 
.A(n_9590),
.B(n_4638),
.C(n_4635),
.D(n_4322),
.Y(n_9723)
);

NOR2xp67_ASAP7_75t_L g9724 ( 
.A(n_9548),
.B(n_6017),
.Y(n_9724)
);

NOR3xp33_ASAP7_75t_SL g9725 ( 
.A(n_9609),
.B(n_4667),
.C(n_4575),
.Y(n_9725)
);

NOR2x1_ASAP7_75t_L g9726 ( 
.A(n_9603),
.B(n_6018),
.Y(n_9726)
);

NAND2xp5_ASAP7_75t_SL g9727 ( 
.A(n_9612),
.B(n_6018),
.Y(n_9727)
);

NAND2xp5_ASAP7_75t_L g9728 ( 
.A(n_9612),
.B(n_6019),
.Y(n_9728)
);

NAND2xp5_ASAP7_75t_L g9729 ( 
.A(n_9586),
.B(n_6019),
.Y(n_9729)
);

OAI211xp5_ASAP7_75t_SL g9730 ( 
.A1(n_9626),
.A2(n_5098),
.B(n_5175),
.C(n_5074),
.Y(n_9730)
);

INVx1_ASAP7_75t_L g9731 ( 
.A(n_9567),
.Y(n_9731)
);

NAND2xp5_ASAP7_75t_SL g9732 ( 
.A(n_9561),
.B(n_6021),
.Y(n_9732)
);

INVx1_ASAP7_75t_L g9733 ( 
.A(n_9606),
.Y(n_9733)
);

NAND3xp33_ASAP7_75t_L g9734 ( 
.A(n_9594),
.B(n_6022),
.C(n_6021),
.Y(n_9734)
);

NOR3x1_ASAP7_75t_L g9735 ( 
.A(n_9608),
.B(n_6023),
.C(n_6022),
.Y(n_9735)
);

INVx1_ASAP7_75t_L g9736 ( 
.A(n_9607),
.Y(n_9736)
);

AOI21xp5_ASAP7_75t_L g9737 ( 
.A1(n_9627),
.A2(n_6031),
.B(n_6023),
.Y(n_9737)
);

NAND2xp5_ASAP7_75t_L g9738 ( 
.A(n_9599),
.B(n_6031),
.Y(n_9738)
);

NOR2xp33_ASAP7_75t_L g9739 ( 
.A(n_9604),
.B(n_6035),
.Y(n_9739)
);

INVx1_ASAP7_75t_L g9740 ( 
.A(n_9625),
.Y(n_9740)
);

AND4x1_ASAP7_75t_L g9741 ( 
.A(n_9628),
.B(n_4676),
.C(n_4610),
.D(n_4614),
.Y(n_9741)
);

AOI221xp5_ASAP7_75t_L g9742 ( 
.A1(n_9589),
.A2(n_6035),
.B1(n_6050),
.B2(n_6047),
.C(n_6040),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_9624),
.Y(n_9743)
);

INVx1_ASAP7_75t_L g9744 ( 
.A(n_9633),
.Y(n_9744)
);

NOR2xp33_ASAP7_75t_L g9745 ( 
.A(n_9640),
.B(n_9588),
.Y(n_9745)
);

NOR2xp67_ASAP7_75t_L g9746 ( 
.A(n_9597),
.B(n_6040),
.Y(n_9746)
);

NOR3x1_ASAP7_75t_L g9747 ( 
.A(n_9639),
.B(n_6050),
.C(n_6047),
.Y(n_9747)
);

NAND2xp5_ASAP7_75t_L g9748 ( 
.A(n_9592),
.B(n_6055),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_9644),
.Y(n_9749)
);

INVx1_ASAP7_75t_L g9750 ( 
.A(n_9632),
.Y(n_9750)
);

AOI22xp5_ASAP7_75t_L g9751 ( 
.A1(n_9643),
.A2(n_5098),
.B1(n_5175),
.B2(n_5074),
.Y(n_9751)
);

OAI221xp5_ASAP7_75t_L g9752 ( 
.A1(n_9623),
.A2(n_6055),
.B1(n_6059),
.B2(n_6058),
.C(n_6057),
.Y(n_9752)
);

AND3x1_ASAP7_75t_L g9753 ( 
.A(n_9557),
.B(n_5175),
.C(n_5074),
.Y(n_9753)
);

NOR2xp67_ASAP7_75t_L g9754 ( 
.A(n_9631),
.B(n_6057),
.Y(n_9754)
);

NAND2xp5_ASAP7_75t_SL g9755 ( 
.A(n_9585),
.B(n_6058),
.Y(n_9755)
);

NAND4xp25_ASAP7_75t_L g9756 ( 
.A(n_9547),
.B(n_4327),
.C(n_4252),
.D(n_5175),
.Y(n_9756)
);

AOI21xp5_ASAP7_75t_L g9757 ( 
.A1(n_9688),
.A2(n_6060),
.B(n_6059),
.Y(n_9757)
);

INVx1_ASAP7_75t_L g9758 ( 
.A(n_9651),
.Y(n_9758)
);

NOR2x1p5_ASAP7_75t_L g9759 ( 
.A(n_9677),
.B(n_5202),
.Y(n_9759)
);

AOI211xp5_ASAP7_75t_L g9760 ( 
.A1(n_9654),
.A2(n_4382),
.B(n_4315),
.C(n_6060),
.Y(n_9760)
);

NAND2xp5_ASAP7_75t_L g9761 ( 
.A(n_9671),
.B(n_6063),
.Y(n_9761)
);

NAND3xp33_ASAP7_75t_SL g9762 ( 
.A(n_9646),
.B(n_4525),
.C(n_4480),
.Y(n_9762)
);

INVx1_ASAP7_75t_L g9763 ( 
.A(n_9667),
.Y(n_9763)
);

NOR3xp33_ASAP7_75t_L g9764 ( 
.A(n_9681),
.B(n_5210),
.C(n_5202),
.Y(n_9764)
);

NAND3xp33_ASAP7_75t_L g9765 ( 
.A(n_9652),
.B(n_6064),
.C(n_6063),
.Y(n_9765)
);

INVx2_ASAP7_75t_L g9766 ( 
.A(n_9670),
.Y(n_9766)
);

NOR2xp33_ASAP7_75t_L g9767 ( 
.A(n_9696),
.B(n_5202),
.Y(n_9767)
);

INVx1_ASAP7_75t_L g9768 ( 
.A(n_9660),
.Y(n_9768)
);

INVx2_ASAP7_75t_L g9769 ( 
.A(n_9658),
.Y(n_9769)
);

INVx2_ASAP7_75t_L g9770 ( 
.A(n_9697),
.Y(n_9770)
);

INVx1_ASAP7_75t_L g9771 ( 
.A(n_9650),
.Y(n_9771)
);

BUFx2_ASAP7_75t_L g9772 ( 
.A(n_9689),
.Y(n_9772)
);

AOI211xp5_ASAP7_75t_L g9773 ( 
.A1(n_9661),
.A2(n_4382),
.B(n_4315),
.C(n_6064),
.Y(n_9773)
);

NAND2xp5_ASAP7_75t_L g9774 ( 
.A(n_9663),
.B(n_6065),
.Y(n_9774)
);

NAND2xp5_ASAP7_75t_L g9775 ( 
.A(n_9685),
.B(n_6065),
.Y(n_9775)
);

AOI322xp5_ASAP7_75t_L g9776 ( 
.A1(n_9649),
.A2(n_6076),
.A3(n_6072),
.B1(n_6073),
.B2(n_6067),
.C1(n_5210),
.C2(n_5202),
.Y(n_9776)
);

AOI221xp5_ASAP7_75t_SL g9777 ( 
.A1(n_9653),
.A2(n_6072),
.B1(n_6076),
.B2(n_6073),
.C(n_6067),
.Y(n_9777)
);

NAND4xp25_ASAP7_75t_L g9778 ( 
.A(n_9707),
.B(n_4327),
.C(n_4676),
.D(n_4342),
.Y(n_9778)
);

OAI22xp5_ASAP7_75t_L g9779 ( 
.A1(n_9680),
.A2(n_5210),
.B1(n_5302),
.B2(n_5267),
.Y(n_9779)
);

AOI21xp5_ASAP7_75t_L g9780 ( 
.A1(n_9647),
.A2(n_5746),
.B(n_5849),
.Y(n_9780)
);

INVx1_ASAP7_75t_L g9781 ( 
.A(n_9662),
.Y(n_9781)
);

OR2x2_ASAP7_75t_L g9782 ( 
.A(n_9709),
.B(n_5210),
.Y(n_9782)
);

AOI21xp5_ASAP7_75t_L g9783 ( 
.A1(n_9655),
.A2(n_5746),
.B(n_5849),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_9690),
.Y(n_9784)
);

AOI21xp5_ASAP7_75t_L g9785 ( 
.A1(n_9659),
.A2(n_6009),
.B(n_4645),
.Y(n_9785)
);

NOR4xp25_ASAP7_75t_L g9786 ( 
.A(n_9656),
.B(n_5302),
.C(n_5328),
.D(n_5267),
.Y(n_9786)
);

NOR4xp25_ASAP7_75t_L g9787 ( 
.A(n_9749),
.B(n_5302),
.C(n_5328),
.D(n_5267),
.Y(n_9787)
);

NAND2xp5_ASAP7_75t_L g9788 ( 
.A(n_9714),
.B(n_5267),
.Y(n_9788)
);

INVx1_ASAP7_75t_L g9789 ( 
.A(n_9682),
.Y(n_9789)
);

NAND4xp25_ASAP7_75t_L g9790 ( 
.A(n_9657),
.B(n_9669),
.C(n_9745),
.D(n_9664),
.Y(n_9790)
);

NOR3xp33_ASAP7_75t_L g9791 ( 
.A(n_9672),
.B(n_5410),
.C(n_5328),
.Y(n_9791)
);

NAND4xp25_ASAP7_75t_L g9792 ( 
.A(n_9686),
.B(n_4342),
.C(n_4358),
.D(n_4248),
.Y(n_9792)
);

AND2x4_ASAP7_75t_SL g9793 ( 
.A(n_9715),
.B(n_5302),
.Y(n_9793)
);

AND2x2_ASAP7_75t_L g9794 ( 
.A(n_9702),
.B(n_5328),
.Y(n_9794)
);

AND2x2_ASAP7_75t_L g9795 ( 
.A(n_9733),
.B(n_5410),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_9698),
.Y(n_9796)
);

NOR3xp33_ASAP7_75t_L g9797 ( 
.A(n_9744),
.B(n_5387),
.C(n_5410),
.Y(n_9797)
);

NOR2xp33_ASAP7_75t_L g9798 ( 
.A(n_9736),
.B(n_5387),
.Y(n_9798)
);

AOI211x1_ASAP7_75t_L g9799 ( 
.A1(n_9713),
.A2(n_5137),
.B(n_5141),
.C(n_5139),
.Y(n_9799)
);

AOI21xp5_ASAP7_75t_L g9800 ( 
.A1(n_9743),
.A2(n_6009),
.B(n_4650),
.Y(n_9800)
);

NAND2xp5_ASAP7_75t_L g9801 ( 
.A(n_9699),
.B(n_5387),
.Y(n_9801)
);

INVx1_ASAP7_75t_L g9802 ( 
.A(n_9666),
.Y(n_9802)
);

AOI21xp5_ASAP7_75t_L g9803 ( 
.A1(n_9746),
.A2(n_6009),
.B(n_4650),
.Y(n_9803)
);

INVx1_ASAP7_75t_L g9804 ( 
.A(n_9674),
.Y(n_9804)
);

NAND2xp5_ASAP7_75t_L g9805 ( 
.A(n_9750),
.B(n_5387),
.Y(n_9805)
);

NAND2xp5_ASAP7_75t_SL g9806 ( 
.A(n_9692),
.B(n_5410),
.Y(n_9806)
);

NAND2xp33_ASAP7_75t_SL g9807 ( 
.A(n_9675),
.B(n_4240),
.Y(n_9807)
);

AND3x1_ASAP7_75t_L g9808 ( 
.A(n_9695),
.B(n_4620),
.C(n_4591),
.Y(n_9808)
);

INVxp67_ASAP7_75t_SL g9809 ( 
.A(n_9724),
.Y(n_9809)
);

NAND2xp5_ASAP7_75t_L g9810 ( 
.A(n_9705),
.B(n_5232),
.Y(n_9810)
);

NAND4xp25_ASAP7_75t_L g9811 ( 
.A(n_9718),
.B(n_4342),
.C(n_4358),
.D(n_4248),
.Y(n_9811)
);

NAND2xp5_ASAP7_75t_L g9812 ( 
.A(n_9739),
.B(n_5232),
.Y(n_9812)
);

INVx1_ASAP7_75t_L g9813 ( 
.A(n_9684),
.Y(n_9813)
);

AOI221x1_ASAP7_75t_L g9814 ( 
.A1(n_9710),
.A2(n_4666),
.B1(n_4620),
.B2(n_4591),
.C(n_4699),
.Y(n_9814)
);

NOR5xp2_ASAP7_75t_L g9815 ( 
.A(n_9719),
.B(n_4578),
.C(n_4570),
.D(n_4520),
.E(n_5139),
.Y(n_9815)
);

NOR2xp33_ASAP7_75t_L g9816 ( 
.A(n_9648),
.B(n_4240),
.Y(n_9816)
);

INVx2_ASAP7_75t_SL g9817 ( 
.A(n_9726),
.Y(n_9817)
);

INVx1_ASAP7_75t_L g9818 ( 
.A(n_9694),
.Y(n_9818)
);

NAND3xp33_ASAP7_75t_SL g9819 ( 
.A(n_9701),
.B(n_9720),
.C(n_9721),
.Y(n_9819)
);

OAI21xp5_ASAP7_75t_L g9820 ( 
.A1(n_9716),
.A2(n_4465),
.B(n_4474),
.Y(n_9820)
);

INVx1_ASAP7_75t_L g9821 ( 
.A(n_9728),
.Y(n_9821)
);

AND2x2_ASAP7_75t_L g9822 ( 
.A(n_9740),
.B(n_5394),
.Y(n_9822)
);

NOR3xp33_ASAP7_75t_L g9823 ( 
.A(n_9731),
.B(n_4620),
.C(n_4591),
.Y(n_9823)
);

AOI22xp33_ASAP7_75t_L g9824 ( 
.A1(n_9700),
.A2(n_4620),
.B1(n_4666),
.B2(n_4591),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_9729),
.Y(n_9825)
);

NOR4xp25_ASAP7_75t_L g9826 ( 
.A(n_9756),
.B(n_9727),
.C(n_9755),
.D(n_9732),
.Y(n_9826)
);

AOI211xp5_ASAP7_75t_L g9827 ( 
.A1(n_9756),
.A2(n_4081),
.B(n_4240),
.C(n_4280),
.Y(n_9827)
);

NAND2xp5_ASAP7_75t_L g9828 ( 
.A(n_9683),
.B(n_5232),
.Y(n_9828)
);

INVx1_ASAP7_75t_L g9829 ( 
.A(n_9747),
.Y(n_9829)
);

A2O1A1Ixp33_ASAP7_75t_L g9830 ( 
.A1(n_9717),
.A2(n_4666),
.B(n_4406),
.C(n_4461),
.Y(n_9830)
);

NAND2xp5_ASAP7_75t_L g9831 ( 
.A(n_9703),
.B(n_5232),
.Y(n_9831)
);

AOI21xp5_ASAP7_75t_SL g9832 ( 
.A1(n_9673),
.A2(n_4461),
.B(n_4397),
.Y(n_9832)
);

NOR2x1_ASAP7_75t_SL g9833 ( 
.A(n_9722),
.B(n_5312),
.Y(n_9833)
);

OAI32xp33_ASAP7_75t_L g9834 ( 
.A1(n_9706),
.A2(n_9687),
.A3(n_9738),
.B1(n_9748),
.B2(n_9676),
.Y(n_9834)
);

NAND3xp33_ASAP7_75t_L g9835 ( 
.A(n_9753),
.B(n_6009),
.C(n_4317),
.Y(n_9835)
);

NOR4xp75_ASAP7_75t_L g9836 ( 
.A(n_9693),
.B(n_4666),
.C(n_4627),
.D(n_4270),
.Y(n_9836)
);

NAND2xp5_ASAP7_75t_SL g9837 ( 
.A(n_9754),
.B(n_4240),
.Y(n_9837)
);

INVx1_ASAP7_75t_L g9838 ( 
.A(n_9735),
.Y(n_9838)
);

INVx1_ASAP7_75t_L g9839 ( 
.A(n_9712),
.Y(n_9839)
);

AOI21xp5_ASAP7_75t_L g9840 ( 
.A1(n_9737),
.A2(n_4628),
.B(n_5312),
.Y(n_9840)
);

AO21x1_ASAP7_75t_L g9841 ( 
.A1(n_9691),
.A2(n_4525),
.B(n_4480),
.Y(n_9841)
);

NAND2xp5_ASAP7_75t_L g9842 ( 
.A(n_9734),
.B(n_5312),
.Y(n_9842)
);

NAND4xp25_ASAP7_75t_L g9843 ( 
.A(n_9668),
.B(n_4358),
.C(n_4370),
.D(n_4248),
.Y(n_9843)
);

NAND2xp5_ASAP7_75t_L g9844 ( 
.A(n_9711),
.B(n_5312),
.Y(n_9844)
);

INVx1_ASAP7_75t_L g9845 ( 
.A(n_9708),
.Y(n_9845)
);

NAND2xp5_ASAP7_75t_SL g9846 ( 
.A(n_9751),
.B(n_4240),
.Y(n_9846)
);

AOI211xp5_ASAP7_75t_L g9847 ( 
.A1(n_9730),
.A2(n_4280),
.B(n_4317),
.C(n_4240),
.Y(n_9847)
);

INVx1_ASAP7_75t_L g9848 ( 
.A(n_9678),
.Y(n_9848)
);

NAND3xp33_ASAP7_75t_L g9849 ( 
.A(n_9725),
.B(n_4317),
.C(n_4280),
.Y(n_9849)
);

OAI211xp5_ASAP7_75t_L g9850 ( 
.A1(n_9704),
.A2(n_4461),
.B(n_4397),
.C(n_4798),
.Y(n_9850)
);

OR2x2_ASAP7_75t_L g9851 ( 
.A(n_9723),
.B(n_5404),
.Y(n_9851)
);

NAND2xp5_ASAP7_75t_L g9852 ( 
.A(n_9742),
.B(n_5404),
.Y(n_9852)
);

AND2x2_ASAP7_75t_L g9853 ( 
.A(n_9741),
.B(n_4586),
.Y(n_9853)
);

NAND4xp25_ASAP7_75t_L g9854 ( 
.A(n_9723),
.B(n_4386),
.C(n_4370),
.D(n_4429),
.Y(n_9854)
);

NAND3xp33_ASAP7_75t_SL g9855 ( 
.A(n_9752),
.B(n_4480),
.C(n_4640),
.Y(n_9855)
);

AOI211xp5_ASAP7_75t_L g9856 ( 
.A1(n_9665),
.A2(n_4280),
.B(n_4317),
.C(n_4240),
.Y(n_9856)
);

NOR3xp33_ASAP7_75t_L g9857 ( 
.A(n_9679),
.B(n_4267),
.C(n_4699),
.Y(n_9857)
);

NAND2xp5_ASAP7_75t_L g9858 ( 
.A(n_9688),
.B(n_5404),
.Y(n_9858)
);

AND2x2_ASAP7_75t_L g9859 ( 
.A(n_9696),
.B(n_4586),
.Y(n_9859)
);

NAND2xp5_ASAP7_75t_L g9860 ( 
.A(n_9688),
.B(n_5404),
.Y(n_9860)
);

INVx1_ASAP7_75t_L g9861 ( 
.A(n_9651),
.Y(n_9861)
);

NAND3xp33_ASAP7_75t_L g9862 ( 
.A(n_9654),
.B(n_4317),
.C(n_4280),
.Y(n_9862)
);

INVx1_ASAP7_75t_L g9863 ( 
.A(n_9651),
.Y(n_9863)
);

NAND4xp25_ASAP7_75t_L g9864 ( 
.A(n_9654),
.B(n_4386),
.C(n_4370),
.D(n_4429),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_9651),
.Y(n_9865)
);

NAND4xp75_ASAP7_75t_L g9866 ( 
.A(n_9658),
.B(n_4798),
.C(n_4821),
.D(n_4397),
.Y(n_9866)
);

NAND2xp5_ASAP7_75t_L g9867 ( 
.A(n_9688),
.B(n_5413),
.Y(n_9867)
);

AOI22xp33_ASAP7_75t_L g9868 ( 
.A1(n_9772),
.A2(n_4303),
.B1(n_4421),
.B2(n_4308),
.Y(n_9868)
);

NAND2xp5_ASAP7_75t_L g9869 ( 
.A(n_9816),
.B(n_5274),
.Y(n_9869)
);

NAND2xp5_ASAP7_75t_L g9870 ( 
.A(n_9771),
.B(n_5274),
.Y(n_9870)
);

INVx2_ASAP7_75t_L g9871 ( 
.A(n_9759),
.Y(n_9871)
);

AOI321xp33_ASAP7_75t_L g9872 ( 
.A1(n_9760),
.A2(n_4492),
.A3(n_4429),
.B1(n_4386),
.B2(n_4493),
.C(n_4478),
.Y(n_9872)
);

INVx1_ASAP7_75t_L g9873 ( 
.A(n_9859),
.Y(n_9873)
);

NAND2xp5_ASAP7_75t_L g9874 ( 
.A(n_9766),
.B(n_5274),
.Y(n_9874)
);

INVxp67_ASAP7_75t_L g9875 ( 
.A(n_9767),
.Y(n_9875)
);

NAND2xp5_ASAP7_75t_L g9876 ( 
.A(n_9795),
.B(n_5282),
.Y(n_9876)
);

INVx1_ASAP7_75t_L g9877 ( 
.A(n_9817),
.Y(n_9877)
);

XNOR2xp5_ASAP7_75t_L g9878 ( 
.A(n_9862),
.B(n_4429),
.Y(n_9878)
);

NAND4xp75_ASAP7_75t_L g9879 ( 
.A(n_9763),
.B(n_4821),
.C(n_4798),
.D(n_4503),
.Y(n_9879)
);

AOI31xp33_ASAP7_75t_L g9880 ( 
.A1(n_9784),
.A2(n_4640),
.A3(n_4603),
.B(n_4667),
.Y(n_9880)
);

OAI211xp5_ASAP7_75t_L g9881 ( 
.A1(n_9826),
.A2(n_5424),
.B(n_5425),
.C(n_5417),
.Y(n_9881)
);

AOI21xp5_ASAP7_75t_L g9882 ( 
.A1(n_9809),
.A2(n_4628),
.B(n_4269),
.Y(n_9882)
);

INVx1_ASAP7_75t_SL g9883 ( 
.A(n_9770),
.Y(n_9883)
);

INVx1_ASAP7_75t_L g9884 ( 
.A(n_9805),
.Y(n_9884)
);

INVxp67_ASAP7_75t_L g9885 ( 
.A(n_9789),
.Y(n_9885)
);

NOR2xp33_ASAP7_75t_L g9886 ( 
.A(n_9769),
.B(n_4280),
.Y(n_9886)
);

AND2x2_ASAP7_75t_L g9887 ( 
.A(n_9794),
.B(n_4533),
.Y(n_9887)
);

NAND2xp5_ASAP7_75t_L g9888 ( 
.A(n_9793),
.B(n_5282),
.Y(n_9888)
);

AOI21xp33_ASAP7_75t_L g9889 ( 
.A1(n_9768),
.A2(n_4208),
.B(n_4205),
.Y(n_9889)
);

INVxp33_ASAP7_75t_L g9890 ( 
.A(n_9790),
.Y(n_9890)
);

AOI21xp5_ASAP7_75t_L g9891 ( 
.A1(n_9758),
.A2(n_9863),
.B(n_9861),
.Y(n_9891)
);

INVx1_ASAP7_75t_L g9892 ( 
.A(n_9788),
.Y(n_9892)
);

AOI22xp5_ASAP7_75t_L g9893 ( 
.A1(n_9764),
.A2(n_9864),
.B1(n_9822),
.B2(n_9849),
.Y(n_9893)
);

NOR2xp33_ASAP7_75t_L g9894 ( 
.A(n_9798),
.B(n_4280),
.Y(n_9894)
);

INVx1_ASAP7_75t_L g9895 ( 
.A(n_9865),
.Y(n_9895)
);

AOI21x1_ASAP7_75t_L g9896 ( 
.A1(n_9781),
.A2(n_4821),
.B(n_4798),
.Y(n_9896)
);

INVx1_ASAP7_75t_L g9897 ( 
.A(n_9761),
.Y(n_9897)
);

NAND2xp5_ASAP7_75t_L g9898 ( 
.A(n_9773),
.B(n_5282),
.Y(n_9898)
);

O2A1O1Ixp33_ASAP7_75t_L g9899 ( 
.A1(n_9839),
.A2(n_4426),
.B(n_4640),
.C(n_4603),
.Y(n_9899)
);

NAND3xp33_ASAP7_75t_L g9900 ( 
.A(n_9845),
.B(n_9848),
.C(n_9829),
.Y(n_9900)
);

NOR3xp33_ASAP7_75t_L g9901 ( 
.A(n_9819),
.B(n_4267),
.C(n_4699),
.Y(n_9901)
);

OAI22xp5_ASAP7_75t_L g9902 ( 
.A1(n_9782),
.A2(n_4303),
.B1(n_4308),
.B2(n_4270),
.Y(n_9902)
);

INVx2_ASAP7_75t_L g9903 ( 
.A(n_9866),
.Y(n_9903)
);

NAND2xp5_ASAP7_75t_L g9904 ( 
.A(n_9853),
.B(n_9776),
.Y(n_9904)
);

AOI22xp5_ASAP7_75t_L g9905 ( 
.A1(n_9807),
.A2(n_4270),
.B1(n_4308),
.B2(n_4303),
.Y(n_9905)
);

OA22x2_ASAP7_75t_L g9906 ( 
.A1(n_9838),
.A2(n_4308),
.B1(n_4313),
.B2(n_4303),
.Y(n_9906)
);

AOI22xp5_ASAP7_75t_L g9907 ( 
.A1(n_9802),
.A2(n_4313),
.B1(n_4391),
.B2(n_4368),
.Y(n_9907)
);

CKINVDCx20_ASAP7_75t_R g9908 ( 
.A(n_9825),
.Y(n_9908)
);

INVxp33_ASAP7_75t_L g9909 ( 
.A(n_9775),
.Y(n_9909)
);

INVx1_ASAP7_75t_L g9910 ( 
.A(n_9867),
.Y(n_9910)
);

NOR2x1_ASAP7_75t_L g9911 ( 
.A(n_9804),
.B(n_4821),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_9774),
.Y(n_9912)
);

AOI22xp5_ASAP7_75t_L g9913 ( 
.A1(n_9791),
.A2(n_4313),
.B1(n_4391),
.B2(n_4368),
.Y(n_9913)
);

INVx1_ASAP7_75t_L g9914 ( 
.A(n_9837),
.Y(n_9914)
);

NAND2xp5_ASAP7_75t_L g9915 ( 
.A(n_9776),
.B(n_5289),
.Y(n_9915)
);

OAI22xp5_ASAP7_75t_L g9916 ( 
.A1(n_9827),
.A2(n_4368),
.B1(n_4391),
.B2(n_4313),
.Y(n_9916)
);

AOI21xp5_ASAP7_75t_L g9917 ( 
.A1(n_9834),
.A2(n_4269),
.B(n_4610),
.Y(n_9917)
);

NAND2xp5_ASAP7_75t_L g9918 ( 
.A(n_9827),
.B(n_5289),
.Y(n_9918)
);

INVx1_ASAP7_75t_L g9919 ( 
.A(n_9858),
.Y(n_9919)
);

INVx1_ASAP7_75t_L g9920 ( 
.A(n_9860),
.Y(n_9920)
);

OR2x2_ASAP7_75t_L g9921 ( 
.A(n_9801),
.B(n_4368),
.Y(n_9921)
);

CKINVDCx20_ASAP7_75t_R g9922 ( 
.A(n_9796),
.Y(n_9922)
);

NOR2xp33_ASAP7_75t_L g9923 ( 
.A(n_9813),
.B(n_4317),
.Y(n_9923)
);

OAI322xp33_ASAP7_75t_L g9924 ( 
.A1(n_9821),
.A2(n_4391),
.A3(n_4421),
.B1(n_4413),
.B2(n_4459),
.C1(n_4416),
.C2(n_4503),
.Y(n_9924)
);

NAND2xp5_ASAP7_75t_L g9925 ( 
.A(n_9777),
.B(n_5289),
.Y(n_9925)
);

OAI211xp5_ASAP7_75t_L g9926 ( 
.A1(n_9818),
.A2(n_5417),
.B(n_5424),
.C(n_5411),
.Y(n_9926)
);

OR2x2_ASAP7_75t_L g9927 ( 
.A(n_9792),
.B(n_4413),
.Y(n_9927)
);

OAI31xp33_ASAP7_75t_L g9928 ( 
.A1(n_9850),
.A2(n_4603),
.A3(n_4640),
.B(n_4492),
.Y(n_9928)
);

AOI22xp5_ASAP7_75t_L g9929 ( 
.A1(n_9797),
.A2(n_4416),
.B1(n_4421),
.B2(n_4413),
.Y(n_9929)
);

OAI21xp5_ASAP7_75t_L g9930 ( 
.A1(n_9765),
.A2(n_9757),
.B(n_9846),
.Y(n_9930)
);

NAND2xp5_ASAP7_75t_L g9931 ( 
.A(n_9856),
.B(n_5292),
.Y(n_9931)
);

OAI22xp5_ASAP7_75t_L g9932 ( 
.A1(n_9851),
.A2(n_4416),
.B1(n_4421),
.B2(n_4413),
.Y(n_9932)
);

XNOR2xp5_ASAP7_75t_L g9933 ( 
.A(n_9778),
.B(n_4492),
.Y(n_9933)
);

AOI221xp5_ASAP7_75t_L g9934 ( 
.A1(n_9832),
.A2(n_4344),
.B1(n_4464),
.B2(n_4340),
.C(n_4317),
.Y(n_9934)
);

NAND2xp5_ASAP7_75t_L g9935 ( 
.A(n_9799),
.B(n_5292),
.Y(n_9935)
);

XNOR2x1_ASAP7_75t_L g9936 ( 
.A(n_9836),
.B(n_4492),
.Y(n_9936)
);

AOI21xp5_ASAP7_75t_L g9937 ( 
.A1(n_9833),
.A2(n_4614),
.B(n_4246),
.Y(n_9937)
);

AOI211xp5_ASAP7_75t_L g9938 ( 
.A1(n_9806),
.A2(n_4340),
.B(n_4464),
.C(n_4344),
.Y(n_9938)
);

AOI21xp5_ASAP7_75t_L g9939 ( 
.A1(n_9844),
.A2(n_4246),
.B(n_4411),
.Y(n_9939)
);

NAND2xp5_ASAP7_75t_L g9940 ( 
.A(n_9823),
.B(n_5292),
.Y(n_9940)
);

INVx2_ASAP7_75t_SL g9941 ( 
.A(n_9810),
.Y(n_9941)
);

HB1xp67_ASAP7_75t_L g9942 ( 
.A(n_9808),
.Y(n_9942)
);

AOI221xp5_ASAP7_75t_L g9943 ( 
.A1(n_9786),
.A2(n_4464),
.B1(n_4542),
.B2(n_4344),
.C(n_4340),
.Y(n_9943)
);

AOI22xp5_ASAP7_75t_L g9944 ( 
.A1(n_9762),
.A2(n_4459),
.B1(n_4416),
.B2(n_4699),
.Y(n_9944)
);

INVx1_ASAP7_75t_L g9945 ( 
.A(n_9842),
.Y(n_9945)
);

NAND2xp33_ASAP7_75t_L g9946 ( 
.A(n_9857),
.B(n_4340),
.Y(n_9946)
);

AND2x2_ASAP7_75t_L g9947 ( 
.A(n_9787),
.B(n_4533),
.Y(n_9947)
);

XNOR2xp5_ASAP7_75t_L g9948 ( 
.A(n_9847),
.B(n_4603),
.Y(n_9948)
);

O2A1O1Ixp33_ASAP7_75t_L g9949 ( 
.A1(n_9830),
.A2(n_4426),
.B(n_4641),
.C(n_4411),
.Y(n_9949)
);

INVx1_ASAP7_75t_L g9950 ( 
.A(n_9904),
.Y(n_9950)
);

NAND2xp5_ASAP7_75t_L g9951 ( 
.A(n_9883),
.B(n_9852),
.Y(n_9951)
);

AOI22xp5_ASAP7_75t_L g9952 ( 
.A1(n_9922),
.A2(n_9855),
.B1(n_9779),
.B2(n_9854),
.Y(n_9952)
);

INVx1_ASAP7_75t_L g9953 ( 
.A(n_9877),
.Y(n_9953)
);

AOI22xp5_ASAP7_75t_L g9954 ( 
.A1(n_9908),
.A2(n_9843),
.B1(n_9841),
.B2(n_9812),
.Y(n_9954)
);

AOI22xp5_ASAP7_75t_L g9955 ( 
.A1(n_9886),
.A2(n_9811),
.B1(n_9831),
.B2(n_9828),
.Y(n_9955)
);

AOI211xp5_ASAP7_75t_SL g9956 ( 
.A1(n_9885),
.A2(n_9785),
.B(n_9780),
.C(n_9783),
.Y(n_9956)
);

NOR2xp33_ASAP7_75t_L g9957 ( 
.A(n_9873),
.B(n_9835),
.Y(n_9957)
);

OAI22xp33_ASAP7_75t_L g9958 ( 
.A1(n_9890),
.A2(n_9814),
.B1(n_9840),
.B2(n_9800),
.Y(n_9958)
);

NOR2x1_ASAP7_75t_L g9959 ( 
.A(n_9900),
.B(n_9815),
.Y(n_9959)
);

NAND2xp5_ASAP7_75t_SL g9960 ( 
.A(n_9895),
.B(n_9824),
.Y(n_9960)
);

NOR2xp33_ASAP7_75t_L g9961 ( 
.A(n_9909),
.B(n_9803),
.Y(n_9961)
);

INVx1_ASAP7_75t_L g9962 ( 
.A(n_9942),
.Y(n_9962)
);

AOI22xp5_ASAP7_75t_L g9963 ( 
.A1(n_9923),
.A2(n_9893),
.B1(n_9903),
.B2(n_9875),
.Y(n_9963)
);

AOI22xp5_ASAP7_75t_L g9964 ( 
.A1(n_9894),
.A2(n_9820),
.B1(n_4459),
.B2(n_4746),
.Y(n_9964)
);

INVx1_ASAP7_75t_SL g9965 ( 
.A(n_9871),
.Y(n_9965)
);

INVx1_ASAP7_75t_L g9966 ( 
.A(n_9874),
.Y(n_9966)
);

INVx1_ASAP7_75t_L g9967 ( 
.A(n_9870),
.Y(n_9967)
);

INVx1_ASAP7_75t_SL g9968 ( 
.A(n_9891),
.Y(n_9968)
);

INVx1_ASAP7_75t_L g9969 ( 
.A(n_9914),
.Y(n_9969)
);

INVx1_ASAP7_75t_L g9970 ( 
.A(n_9930),
.Y(n_9970)
);

AOI221xp5_ASAP7_75t_L g9971 ( 
.A1(n_9946),
.A2(n_4340),
.B1(n_4551),
.B2(n_4464),
.C(n_4344),
.Y(n_9971)
);

INVx1_ASAP7_75t_L g9972 ( 
.A(n_9910),
.Y(n_9972)
);

INVx1_ASAP7_75t_L g9973 ( 
.A(n_9912),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_9884),
.Y(n_9974)
);

INVx1_ASAP7_75t_L g9975 ( 
.A(n_9892),
.Y(n_9975)
);

AOI22xp5_ASAP7_75t_L g9976 ( 
.A1(n_9936),
.A2(n_4459),
.B1(n_4746),
.B2(n_4340),
.Y(n_9976)
);

AND2x4_ASAP7_75t_L g9977 ( 
.A(n_9897),
.B(n_4340),
.Y(n_9977)
);

INVx1_ASAP7_75t_L g9978 ( 
.A(n_9945),
.Y(n_9978)
);

NOR2x1_ASAP7_75t_L g9979 ( 
.A(n_9919),
.B(n_4049),
.Y(n_9979)
);

NAND2xp5_ASAP7_75t_L g9980 ( 
.A(n_9933),
.B(n_9947),
.Y(n_9980)
);

AOI22xp5_ASAP7_75t_L g9981 ( 
.A1(n_9906),
.A2(n_4746),
.B1(n_4344),
.B2(n_4542),
.Y(n_9981)
);

NOR2x1_ASAP7_75t_SL g9982 ( 
.A(n_9881),
.B(n_4138),
.Y(n_9982)
);

NAND2xp5_ASAP7_75t_L g9983 ( 
.A(n_9941),
.B(n_5406),
.Y(n_9983)
);

AND2x4_ASAP7_75t_L g9984 ( 
.A(n_9920),
.B(n_9898),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_9925),
.Y(n_9985)
);

NOR2x1_ASAP7_75t_L g9986 ( 
.A(n_9911),
.B(n_4049),
.Y(n_9986)
);

AOI22xp5_ASAP7_75t_L g9987 ( 
.A1(n_9932),
.A2(n_4746),
.B1(n_4344),
.B2(n_4542),
.Y(n_9987)
);

NOR2x1_ASAP7_75t_L g9988 ( 
.A(n_9915),
.B(n_4049),
.Y(n_9988)
);

AOI221xp5_ASAP7_75t_SL g9989 ( 
.A1(n_9869),
.A2(n_4542),
.B1(n_4551),
.B2(n_4464),
.C(n_4344),
.Y(n_9989)
);

OR2x2_ASAP7_75t_L g9990 ( 
.A(n_9927),
.B(n_5334),
.Y(n_9990)
);

INVx1_ASAP7_75t_L g9991 ( 
.A(n_9918),
.Y(n_9991)
);

INVx1_ASAP7_75t_L g9992 ( 
.A(n_9921),
.Y(n_9992)
);

AOI22xp5_ASAP7_75t_L g9993 ( 
.A1(n_9878),
.A2(n_9901),
.B1(n_9887),
.B2(n_9948),
.Y(n_9993)
);

AOI221xp5_ASAP7_75t_L g9994 ( 
.A1(n_9939),
.A2(n_4464),
.B1(n_4559),
.B2(n_4551),
.C(n_4542),
.Y(n_9994)
);

AOI22xp5_ASAP7_75t_L g9995 ( 
.A1(n_9931),
.A2(n_4464),
.B1(n_4551),
.B2(n_4542),
.Y(n_9995)
);

AOI22xp5_ASAP7_75t_L g9996 ( 
.A1(n_9902),
.A2(n_4542),
.B1(n_4559),
.B2(n_4551),
.Y(n_9996)
);

INVx1_ASAP7_75t_L g9997 ( 
.A(n_9935),
.Y(n_9997)
);

NAND2xp5_ASAP7_75t_L g9998 ( 
.A(n_9928),
.B(n_5425),
.Y(n_9998)
);

INVxp33_ASAP7_75t_SL g9999 ( 
.A(n_9940),
.Y(n_9999)
);

NOR4xp25_ASAP7_75t_L g10000 ( 
.A(n_9926),
.B(n_5150),
.C(n_5153),
.D(n_5141),
.Y(n_10000)
);

INVx1_ASAP7_75t_L g10001 ( 
.A(n_9888),
.Y(n_10001)
);

INVx1_ASAP7_75t_L g10002 ( 
.A(n_9876),
.Y(n_10002)
);

NOR4xp25_ASAP7_75t_L g10003 ( 
.A(n_9899),
.B(n_5153),
.C(n_5159),
.D(n_5150),
.Y(n_10003)
);

NAND2xp5_ASAP7_75t_L g10004 ( 
.A(n_9938),
.B(n_5428),
.Y(n_10004)
);

AOI22xp5_ASAP7_75t_L g10005 ( 
.A1(n_9934),
.A2(n_4551),
.B1(n_4560),
.B2(n_4559),
.Y(n_10005)
);

INVx2_ASAP7_75t_L g10006 ( 
.A(n_9896),
.Y(n_10006)
);

INVx2_ASAP7_75t_L g10007 ( 
.A(n_9879),
.Y(n_10007)
);

AOI22xp5_ASAP7_75t_L g10008 ( 
.A1(n_9917),
.A2(n_4551),
.B1(n_4560),
.B2(n_4559),
.Y(n_10008)
);

NOR2x1_ASAP7_75t_L g10009 ( 
.A(n_9937),
.B(n_4049),
.Y(n_10009)
);

NOR2x1_ASAP7_75t_L g10010 ( 
.A(n_9882),
.B(n_4063),
.Y(n_10010)
);

INVx1_ASAP7_75t_L g10011 ( 
.A(n_9944),
.Y(n_10011)
);

AOI22xp5_ASAP7_75t_L g10012 ( 
.A1(n_9868),
.A2(n_4560),
.B1(n_4559),
.B2(n_4557),
.Y(n_10012)
);

NAND4xp25_ASAP7_75t_L g10013 ( 
.A(n_9872),
.B(n_4104),
.C(n_4106),
.D(n_4103),
.Y(n_10013)
);

NOR3xp33_ASAP7_75t_L g10014 ( 
.A(n_9949),
.B(n_4267),
.C(n_4111),
.Y(n_10014)
);

NOR2x1_ASAP7_75t_L g10015 ( 
.A(n_9924),
.B(n_4063),
.Y(n_10015)
);

INVx1_ASAP7_75t_L g10016 ( 
.A(n_9905),
.Y(n_10016)
);

AOI31xp33_ASAP7_75t_L g10017 ( 
.A1(n_9943),
.A2(n_4503),
.A3(n_4588),
.B(n_4557),
.Y(n_10017)
);

INVx1_ASAP7_75t_L g10018 ( 
.A(n_9907),
.Y(n_10018)
);

INVx1_ASAP7_75t_L g10019 ( 
.A(n_9982),
.Y(n_10019)
);

INVx1_ASAP7_75t_L g10020 ( 
.A(n_9953),
.Y(n_10020)
);

NOR3xp33_ASAP7_75t_L g10021 ( 
.A(n_9950),
.B(n_9889),
.C(n_9880),
.Y(n_10021)
);

NAND3x1_ASAP7_75t_SL g10022 ( 
.A(n_9959),
.B(n_9907),
.C(n_9916),
.Y(n_10022)
);

INVx1_ASAP7_75t_L g10023 ( 
.A(n_9980),
.Y(n_10023)
);

AOI211x1_ASAP7_75t_SL g10024 ( 
.A1(n_10007),
.A2(n_9929),
.B(n_9913),
.C(n_5337),
.Y(n_10024)
);

NOR4xp25_ASAP7_75t_L g10025 ( 
.A(n_9968),
.B(n_5169),
.C(n_5176),
.D(n_5159),
.Y(n_10025)
);

AOI32xp33_ASAP7_75t_L g10026 ( 
.A1(n_9962),
.A2(n_4642),
.A3(n_4714),
.B1(n_4588),
.B2(n_4557),
.Y(n_10026)
);

NAND2xp5_ASAP7_75t_L g10027 ( 
.A(n_9977),
.B(n_5334),
.Y(n_10027)
);

AND2x4_ASAP7_75t_SL g10028 ( 
.A(n_9969),
.B(n_4559),
.Y(n_10028)
);

NAND2xp5_ASAP7_75t_SL g10029 ( 
.A(n_9965),
.B(n_4559),
.Y(n_10029)
);

NAND2xp5_ASAP7_75t_L g10030 ( 
.A(n_9977),
.B(n_5334),
.Y(n_10030)
);

XNOR2xp5_ASAP7_75t_L g10031 ( 
.A(n_9963),
.B(n_4537),
.Y(n_10031)
);

INVx1_ASAP7_75t_L g10032 ( 
.A(n_9988),
.Y(n_10032)
);

NOR2xp33_ASAP7_75t_L g10033 ( 
.A(n_9970),
.B(n_3936),
.Y(n_10033)
);

AND2x2_ASAP7_75t_L g10034 ( 
.A(n_9973),
.B(n_4537),
.Y(n_10034)
);

NAND2xp5_ASAP7_75t_L g10035 ( 
.A(n_9957),
.B(n_5337),
.Y(n_10035)
);

INVx1_ASAP7_75t_L g10036 ( 
.A(n_9979),
.Y(n_10036)
);

OAI211xp5_ASAP7_75t_L g10037 ( 
.A1(n_9960),
.A2(n_4116),
.B(n_4126),
.C(n_4115),
.Y(n_10037)
);

INVx1_ASAP7_75t_L g10038 ( 
.A(n_10006),
.Y(n_10038)
);

HB1xp67_ASAP7_75t_L g10039 ( 
.A(n_9986),
.Y(n_10039)
);

BUFx3_ASAP7_75t_L g10040 ( 
.A(n_9972),
.Y(n_10040)
);

INVxp67_ASAP7_75t_L g10041 ( 
.A(n_9961),
.Y(n_10041)
);

NOR3xp33_ASAP7_75t_L g10042 ( 
.A(n_9951),
.B(n_4111),
.C(n_4063),
.Y(n_10042)
);

NAND2xp5_ASAP7_75t_SL g10043 ( 
.A(n_9954),
.B(n_4560),
.Y(n_10043)
);

OR2x2_ASAP7_75t_L g10044 ( 
.A(n_10013),
.B(n_5337),
.Y(n_10044)
);

NOR3xp33_ASAP7_75t_L g10045 ( 
.A(n_9974),
.B(n_4111),
.C(n_4063),
.Y(n_10045)
);

INVx1_ASAP7_75t_L g10046 ( 
.A(n_10009),
.Y(n_10046)
);

NOR2xp33_ASAP7_75t_L g10047 ( 
.A(n_9999),
.B(n_3936),
.Y(n_10047)
);

NOR3xp33_ASAP7_75t_L g10048 ( 
.A(n_9975),
.B(n_4111),
.C(n_4245),
.Y(n_10048)
);

HB1xp67_ASAP7_75t_L g10049 ( 
.A(n_9997),
.Y(n_10049)
);

INVx1_ASAP7_75t_L g10050 ( 
.A(n_10018),
.Y(n_10050)
);

INVxp67_ASAP7_75t_L g10051 ( 
.A(n_9985),
.Y(n_10051)
);

OAI22xp5_ASAP7_75t_L g10052 ( 
.A1(n_9976),
.A2(n_4499),
.B1(n_4560),
.B2(n_4588),
.Y(n_10052)
);

NAND3x1_ASAP7_75t_L g10053 ( 
.A(n_9967),
.B(n_5176),
.C(n_5169),
.Y(n_10053)
);

NAND2x1_ASAP7_75t_L g10054 ( 
.A(n_9984),
.B(n_4641),
.Y(n_10054)
);

INVx1_ASAP7_75t_L g10055 ( 
.A(n_9983),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_SL g10056 ( 
.A(n_9952),
.B(n_4560),
.Y(n_10056)
);

INVx1_ASAP7_75t_L g10057 ( 
.A(n_9993),
.Y(n_10057)
);

NAND2xp5_ASAP7_75t_L g10058 ( 
.A(n_9958),
.B(n_5353),
.Y(n_10058)
);

NAND2xp5_ASAP7_75t_SL g10059 ( 
.A(n_9955),
.B(n_4560),
.Y(n_10059)
);

INVx2_ASAP7_75t_L g10060 ( 
.A(n_9990),
.Y(n_10060)
);

AND2x2_ASAP7_75t_L g10061 ( 
.A(n_9992),
.B(n_4537),
.Y(n_10061)
);

NAND3xp33_ASAP7_75t_L g10062 ( 
.A(n_9956),
.B(n_5428),
.C(n_5181),
.Y(n_10062)
);

NAND3xp33_ASAP7_75t_L g10063 ( 
.A(n_9978),
.B(n_5181),
.C(n_5178),
.Y(n_10063)
);

NAND2xp5_ASAP7_75t_L g10064 ( 
.A(n_9966),
.B(n_10002),
.Y(n_10064)
);

INVx1_ASAP7_75t_L g10065 ( 
.A(n_9991),
.Y(n_10065)
);

AOI21xp5_ASAP7_75t_L g10066 ( 
.A1(n_9984),
.A2(n_4426),
.B(n_4411),
.Y(n_10066)
);

INVx1_ASAP7_75t_L g10067 ( 
.A(n_10016),
.Y(n_10067)
);

NAND2xp5_ASAP7_75t_L g10068 ( 
.A(n_10001),
.B(n_5353),
.Y(n_10068)
);

NAND2xp5_ASAP7_75t_L g10069 ( 
.A(n_10011),
.B(n_5353),
.Y(n_10069)
);

NAND2xp5_ASAP7_75t_SL g10070 ( 
.A(n_10015),
.B(n_4642),
.Y(n_10070)
);

INVx1_ASAP7_75t_L g10071 ( 
.A(n_10010),
.Y(n_10071)
);

AOI22xp33_ASAP7_75t_L g10072 ( 
.A1(n_10014),
.A2(n_9994),
.B1(n_9998),
.B2(n_9971),
.Y(n_10072)
);

AND2x2_ASAP7_75t_L g10073 ( 
.A(n_10008),
.B(n_4537),
.Y(n_10073)
);

NAND2xp5_ASAP7_75t_L g10074 ( 
.A(n_10003),
.B(n_5356),
.Y(n_10074)
);

OAI21xp33_ASAP7_75t_L g10075 ( 
.A1(n_10031),
.A2(n_10017),
.B(n_9964),
.Y(n_10075)
);

NOR2x1_ASAP7_75t_L g10076 ( 
.A(n_10040),
.B(n_10004),
.Y(n_10076)
);

NAND5xp2_ASAP7_75t_L g10077 ( 
.A(n_10033),
.B(n_9989),
.C(n_10012),
.D(n_9987),
.E(n_9995),
.Y(n_10077)
);

NOR3xp33_ASAP7_75t_SL g10078 ( 
.A(n_10050),
.B(n_10000),
.C(n_10005),
.Y(n_10078)
);

NAND4xp75_ASAP7_75t_L g10079 ( 
.A(n_10020),
.B(n_9981),
.C(n_9996),
.D(n_4714),
.Y(n_10079)
);

NOR2x1p5_ASAP7_75t_L g10080 ( 
.A(n_10067),
.B(n_10019),
.Y(n_10080)
);

NAND2xp5_ASAP7_75t_L g10081 ( 
.A(n_10034),
.B(n_4205),
.Y(n_10081)
);

NAND5xp2_ASAP7_75t_L g10082 ( 
.A(n_10047),
.B(n_10057),
.C(n_10023),
.D(n_10021),
.E(n_10041),
.Y(n_10082)
);

NAND4xp75_ASAP7_75t_L g10083 ( 
.A(n_10065),
.B(n_4714),
.C(n_4721),
.D(n_4642),
.Y(n_10083)
);

AOI211xp5_ASAP7_75t_SL g10084 ( 
.A1(n_10051),
.A2(n_4597),
.B(n_5182),
.C(n_5178),
.Y(n_10084)
);

NOR2x1_ASAP7_75t_L g10085 ( 
.A(n_10036),
.B(n_4123),
.Y(n_10085)
);

NOR2x1_ASAP7_75t_L g10086 ( 
.A(n_10046),
.B(n_4123),
.Y(n_10086)
);

OR3x1_ASAP7_75t_L g10087 ( 
.A(n_10038),
.B(n_10071),
.C(n_10055),
.Y(n_10087)
);

NOR3xp33_ASAP7_75t_L g10088 ( 
.A(n_10022),
.B(n_4250),
.C(n_4245),
.Y(n_10088)
);

NAND4xp25_ASAP7_75t_SL g10089 ( 
.A(n_10072),
.B(n_5183),
.C(n_5190),
.D(n_5182),
.Y(n_10089)
);

NOR2x1_ASAP7_75t_L g10090 ( 
.A(n_10032),
.B(n_4152),
.Y(n_10090)
);

NOR2x1_ASAP7_75t_L g10091 ( 
.A(n_10060),
.B(n_4152),
.Y(n_10091)
);

NAND2xp5_ASAP7_75t_L g10092 ( 
.A(n_10061),
.B(n_4205),
.Y(n_10092)
);

NOR2xp67_ASAP7_75t_L g10093 ( 
.A(n_10039),
.B(n_3936),
.Y(n_10093)
);

NAND2xp5_ASAP7_75t_L g10094 ( 
.A(n_10049),
.B(n_4205),
.Y(n_10094)
);

NOR3xp33_ASAP7_75t_L g10095 ( 
.A(n_10064),
.B(n_10043),
.C(n_10056),
.Y(n_10095)
);

NOR3xp33_ASAP7_75t_L g10096 ( 
.A(n_10058),
.B(n_4250),
.C(n_4245),
.Y(n_10096)
);

OAI211xp5_ASAP7_75t_SL g10097 ( 
.A1(n_10024),
.A2(n_5190),
.B(n_5194),
.C(n_5183),
.Y(n_10097)
);

NAND3xp33_ASAP7_75t_L g10098 ( 
.A(n_10070),
.B(n_3878),
.C(n_3864),
.Y(n_10098)
);

NAND4xp75_ASAP7_75t_L g10099 ( 
.A(n_10059),
.B(n_4741),
.C(n_4721),
.D(n_5194),
.Y(n_10099)
);

NOR3xp33_ASAP7_75t_SL g10100 ( 
.A(n_10029),
.B(n_4597),
.C(n_4690),
.Y(n_10100)
);

AOI221xp5_ASAP7_75t_L g10101 ( 
.A1(n_10069),
.A2(n_5203),
.B1(n_5205),
.B2(n_5199),
.C(n_5196),
.Y(n_10101)
);

INVx1_ASAP7_75t_L g10102 ( 
.A(n_10035),
.Y(n_10102)
);

NOR3xp33_ASAP7_75t_L g10103 ( 
.A(n_10068),
.B(n_4251),
.C(n_4250),
.Y(n_10103)
);

NOR2x1_ASAP7_75t_L g10104 ( 
.A(n_10062),
.B(n_4164),
.Y(n_10104)
);

NOR3xp33_ASAP7_75t_L g10105 ( 
.A(n_10042),
.B(n_10045),
.C(n_10044),
.Y(n_10105)
);

NOR3xp33_ASAP7_75t_L g10106 ( 
.A(n_10052),
.B(n_4261),
.C(n_4251),
.Y(n_10106)
);

AND2x4_ASAP7_75t_L g10107 ( 
.A(n_10028),
.B(n_3902),
.Y(n_10107)
);

INVx1_ASAP7_75t_L g10108 ( 
.A(n_10024),
.Y(n_10108)
);

NAND4xp25_ASAP7_75t_L g10109 ( 
.A(n_10063),
.B(n_4104),
.C(n_4106),
.D(n_4103),
.Y(n_10109)
);

NAND4xp25_ASAP7_75t_SL g10110 ( 
.A(n_10074),
.B(n_5199),
.C(n_5203),
.D(n_5196),
.Y(n_10110)
);

AND3x4_ASAP7_75t_L g10111 ( 
.A(n_10025),
.B(n_3909),
.C(n_3902),
.Y(n_10111)
);

NOR3xp33_ASAP7_75t_SL g10112 ( 
.A(n_10037),
.B(n_4690),
.C(n_4678),
.Y(n_10112)
);

XOR2x2_ASAP7_75t_L g10113 ( 
.A(n_10053),
.B(n_4010),
.Y(n_10113)
);

NAND3xp33_ASAP7_75t_L g10114 ( 
.A(n_10073),
.B(n_3878),
.C(n_3864),
.Y(n_10114)
);

INVx1_ASAP7_75t_L g10115 ( 
.A(n_10027),
.Y(n_10115)
);

NAND2x1_ASAP7_75t_SL g10116 ( 
.A(n_10054),
.B(n_4081),
.Y(n_10116)
);

NOR3xp33_ASAP7_75t_L g10117 ( 
.A(n_10030),
.B(n_4261),
.C(n_4251),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_10048),
.Y(n_10118)
);

NAND2xp5_ASAP7_75t_SL g10119 ( 
.A(n_10026),
.B(n_4721),
.Y(n_10119)
);

INVx2_ASAP7_75t_L g10120 ( 
.A(n_10066),
.Y(n_10120)
);

AND2x4_ASAP7_75t_L g10121 ( 
.A(n_10034),
.B(n_3902),
.Y(n_10121)
);

NAND2xp5_ASAP7_75t_SL g10122 ( 
.A(n_10050),
.B(n_4741),
.Y(n_10122)
);

NOR4xp25_ASAP7_75t_L g10123 ( 
.A(n_10050),
.B(n_5205),
.C(n_5213),
.D(n_5206),
.Y(n_10123)
);

NOR5xp2_ASAP7_75t_L g10124 ( 
.A(n_10108),
.B(n_4578),
.C(n_4570),
.D(n_4520),
.E(n_5206),
.Y(n_10124)
);

NAND4xp75_ASAP7_75t_L g10125 ( 
.A(n_10076),
.B(n_4741),
.C(n_5221),
.D(n_5213),
.Y(n_10125)
);

NOR2x1_ASAP7_75t_L g10126 ( 
.A(n_10087),
.B(n_4164),
.Y(n_10126)
);

NOR4xp25_ASAP7_75t_L g10127 ( 
.A(n_10115),
.B(n_5221),
.C(n_5226),
.D(n_5222),
.Y(n_10127)
);

XOR2xp5_ASAP7_75t_L g10128 ( 
.A(n_10102),
.B(n_3909),
.Y(n_10128)
);

NAND4xp25_ASAP7_75t_L g10129 ( 
.A(n_10082),
.B(n_4104),
.C(n_4106),
.D(n_4103),
.Y(n_10129)
);

NOR3xp33_ASAP7_75t_L g10130 ( 
.A(n_10095),
.B(n_4261),
.C(n_4237),
.Y(n_10130)
);

HB1xp67_ASAP7_75t_L g10131 ( 
.A(n_10080),
.Y(n_10131)
);

NOR2x1_ASAP7_75t_L g10132 ( 
.A(n_10120),
.B(n_3909),
.Y(n_10132)
);

OAI22xp5_ASAP7_75t_L g10133 ( 
.A1(n_10098),
.A2(n_5226),
.B1(n_5229),
.B2(n_5222),
.Y(n_10133)
);

INVx2_ASAP7_75t_L g10134 ( 
.A(n_10113),
.Y(n_10134)
);

INVx4_ASAP7_75t_L g10135 ( 
.A(n_10118),
.Y(n_10135)
);

AOI311xp33_ASAP7_75t_L g10136 ( 
.A1(n_10105),
.A2(n_5243),
.A3(n_5246),
.B(n_5230),
.C(n_5229),
.Y(n_10136)
);

OAI21xp33_ASAP7_75t_L g10137 ( 
.A1(n_10075),
.A2(n_4056),
.B(n_4037),
.Y(n_10137)
);

NOR3xp33_ASAP7_75t_L g10138 ( 
.A(n_10077),
.B(n_4237),
.C(n_4230),
.Y(n_10138)
);

AND3x4_ASAP7_75t_L g10139 ( 
.A(n_10093),
.B(n_4001),
.C(n_3999),
.Y(n_10139)
);

NOR3xp33_ASAP7_75t_L g10140 ( 
.A(n_10079),
.B(n_4237),
.C(n_4230),
.Y(n_10140)
);

INVxp67_ASAP7_75t_L g10141 ( 
.A(n_10078),
.Y(n_10141)
);

NAND3xp33_ASAP7_75t_SL g10142 ( 
.A(n_10111),
.B(n_4149),
.C(n_4395),
.Y(n_10142)
);

INVx1_ASAP7_75t_L g10143 ( 
.A(n_10116),
.Y(n_10143)
);

NOR2x1_ASAP7_75t_L g10144 ( 
.A(n_10090),
.B(n_4641),
.Y(n_10144)
);

NOR2xp33_ASAP7_75t_L g10145 ( 
.A(n_10121),
.B(n_3958),
.Y(n_10145)
);

INVx2_ASAP7_75t_L g10146 ( 
.A(n_10107),
.Y(n_10146)
);

NAND4xp75_ASAP7_75t_L g10147 ( 
.A(n_10104),
.B(n_5243),
.C(n_5246),
.D(n_5230),
.Y(n_10147)
);

NOR2xp33_ASAP7_75t_L g10148 ( 
.A(n_10121),
.B(n_10122),
.Y(n_10148)
);

AND2x2_ASAP7_75t_L g10149 ( 
.A(n_10107),
.B(n_4641),
.Y(n_10149)
);

INVx2_ASAP7_75t_SL g10150 ( 
.A(n_10086),
.Y(n_10150)
);

OR2x2_ASAP7_75t_L g10151 ( 
.A(n_10109),
.B(n_4426),
.Y(n_10151)
);

NAND5xp2_ASAP7_75t_L g10152 ( 
.A(n_10094),
.B(n_4395),
.C(n_4684),
.D(n_4709),
.E(n_4136),
.Y(n_10152)
);

AND2x4_ASAP7_75t_L g10153 ( 
.A(n_10114),
.B(n_4586),
.Y(n_10153)
);

AND2x4_ASAP7_75t_L g10154 ( 
.A(n_10085),
.B(n_4056),
.Y(n_10154)
);

NOR2x1_ASAP7_75t_L g10155 ( 
.A(n_10091),
.B(n_4641),
.Y(n_10155)
);

INVx2_ASAP7_75t_L g10156 ( 
.A(n_10099),
.Y(n_10156)
);

OR2x2_ASAP7_75t_L g10157 ( 
.A(n_10119),
.B(n_4426),
.Y(n_10157)
);

NOR2x1_ASAP7_75t_L g10158 ( 
.A(n_10110),
.B(n_4411),
.Y(n_10158)
);

NOR2x1_ASAP7_75t_L g10159 ( 
.A(n_10089),
.B(n_4411),
.Y(n_10159)
);

INVx3_ASAP7_75t_L g10160 ( 
.A(n_10154),
.Y(n_10160)
);

AND2x2_ASAP7_75t_L g10161 ( 
.A(n_10126),
.B(n_10112),
.Y(n_10161)
);

NOR4xp25_ASAP7_75t_L g10162 ( 
.A(n_10141),
.B(n_10097),
.C(n_10081),
.D(n_10092),
.Y(n_10162)
);

NAND2x1p5_ASAP7_75t_L g10163 ( 
.A(n_10146),
.B(n_10100),
.Y(n_10163)
);

NAND4xp75_ASAP7_75t_L g10164 ( 
.A(n_10143),
.B(n_10101),
.C(n_10083),
.D(n_10123),
.Y(n_10164)
);

AND2x4_ASAP7_75t_L g10165 ( 
.A(n_10131),
.B(n_10106),
.Y(n_10165)
);

AND4x1_ASAP7_75t_L g10166 ( 
.A(n_10148),
.B(n_10132),
.C(n_10145),
.D(n_10144),
.Y(n_10166)
);

NOR2x1p5_ASAP7_75t_L g10167 ( 
.A(n_10134),
.B(n_10084),
.Y(n_10167)
);

XOR2xp5_ASAP7_75t_L g10168 ( 
.A(n_10128),
.B(n_10088),
.Y(n_10168)
);

OR2x2_ASAP7_75t_L g10169 ( 
.A(n_10129),
.B(n_10096),
.Y(n_10169)
);

NAND3xp33_ASAP7_75t_L g10170 ( 
.A(n_10135),
.B(n_10103),
.C(n_10117),
.Y(n_10170)
);

NOR2x1_ASAP7_75t_L g10171 ( 
.A(n_10156),
.B(n_4166),
.Y(n_10171)
);

INVx2_ASAP7_75t_L g10172 ( 
.A(n_10150),
.Y(n_10172)
);

AOI22xp33_ASAP7_75t_L g10173 ( 
.A1(n_10139),
.A2(n_3986),
.B1(n_3984),
.B2(n_4183),
.Y(n_10173)
);

AND2x2_ASAP7_75t_L g10174 ( 
.A(n_10153),
.B(n_4411),
.Y(n_10174)
);

NOR2xp67_ASAP7_75t_L g10175 ( 
.A(n_10142),
.B(n_3958),
.Y(n_10175)
);

NAND2x1p5_ASAP7_75t_L g10176 ( 
.A(n_10155),
.B(n_10158),
.Y(n_10176)
);

OR2x2_ASAP7_75t_L g10177 ( 
.A(n_10157),
.B(n_4200),
.Y(n_10177)
);

AND2x2_ASAP7_75t_L g10178 ( 
.A(n_10149),
.B(n_4133),
.Y(n_10178)
);

NAND3xp33_ASAP7_75t_SL g10179 ( 
.A(n_10124),
.B(n_4149),
.C(n_4044),
.Y(n_10179)
);

AND2x2_ASAP7_75t_L g10180 ( 
.A(n_10159),
.B(n_4133),
.Y(n_10180)
);

NOR2xp33_ASAP7_75t_L g10181 ( 
.A(n_10137),
.B(n_10151),
.Y(n_10181)
);

INVx1_ASAP7_75t_L g10182 ( 
.A(n_10147),
.Y(n_10182)
);

NOR2xp33_ASAP7_75t_L g10183 ( 
.A(n_10125),
.B(n_3958),
.Y(n_10183)
);

INVx1_ASAP7_75t_L g10184 ( 
.A(n_10140),
.Y(n_10184)
);

INVx1_ASAP7_75t_SL g10185 ( 
.A(n_10133),
.Y(n_10185)
);

NAND2xp5_ASAP7_75t_L g10186 ( 
.A(n_10138),
.B(n_10127),
.Y(n_10186)
);

OR2x2_ASAP7_75t_SL g10187 ( 
.A(n_10152),
.B(n_3788),
.Y(n_10187)
);

NAND5xp2_ASAP7_75t_L g10188 ( 
.A(n_10163),
.B(n_10136),
.C(n_10130),
.D(n_4395),
.E(n_4136),
.Y(n_10188)
);

HB1xp67_ASAP7_75t_L g10189 ( 
.A(n_10176),
.Y(n_10189)
);

INVx2_ASAP7_75t_L g10190 ( 
.A(n_10172),
.Y(n_10190)
);

INVx2_ASAP7_75t_L g10191 ( 
.A(n_10161),
.Y(n_10191)
);

INVxp67_ASAP7_75t_L g10192 ( 
.A(n_10168),
.Y(n_10192)
);

INVx2_ASAP7_75t_L g10193 ( 
.A(n_10160),
.Y(n_10193)
);

INVx1_ASAP7_75t_L g10194 ( 
.A(n_10186),
.Y(n_10194)
);

INVx1_ASAP7_75t_L g10195 ( 
.A(n_10164),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_10182),
.Y(n_10196)
);

AOI222xp33_ASAP7_75t_L g10197 ( 
.A1(n_10175),
.A2(n_5272),
.B1(n_5263),
.B2(n_5275),
.C1(n_5264),
.C2(n_5259),
.Y(n_10197)
);

NAND2xp5_ASAP7_75t_L g10198 ( 
.A(n_10183),
.B(n_4208),
.Y(n_10198)
);

AOI222xp33_ASAP7_75t_L g10199 ( 
.A1(n_10179),
.A2(n_5272),
.B1(n_5263),
.B2(n_5275),
.C1(n_5264),
.C2(n_5259),
.Y(n_10199)
);

OAI221xp5_ASAP7_75t_SL g10200 ( 
.A1(n_10166),
.A2(n_5278),
.B1(n_5295),
.B2(n_5291),
.C(n_5287),
.Y(n_10200)
);

NAND4xp75_ASAP7_75t_L g10201 ( 
.A(n_10184),
.B(n_4168),
.C(n_4170),
.D(n_4167),
.Y(n_10201)
);

INVx2_ASAP7_75t_L g10202 ( 
.A(n_10171),
.Y(n_10202)
);

NAND2xp5_ASAP7_75t_L g10203 ( 
.A(n_10180),
.B(n_4208),
.Y(n_10203)
);

AND2x4_ASAP7_75t_L g10204 ( 
.A(n_10167),
.B(n_4727),
.Y(n_10204)
);

INVx1_ASAP7_75t_L g10205 ( 
.A(n_10169),
.Y(n_10205)
);

INVx2_ASAP7_75t_L g10206 ( 
.A(n_10165),
.Y(n_10206)
);

AOI22xp5_ASAP7_75t_L g10207 ( 
.A1(n_10181),
.A2(n_4138),
.B1(n_3985),
.B2(n_4005),
.Y(n_10207)
);

AOI21xp33_ASAP7_75t_L g10208 ( 
.A1(n_10185),
.A2(n_3985),
.B(n_3965),
.Y(n_10208)
);

AOI222xp33_ASAP7_75t_L g10209 ( 
.A1(n_10170),
.A2(n_5295),
.B1(n_5287),
.B2(n_5300),
.C1(n_5291),
.C2(n_5278),
.Y(n_10209)
);

INVx2_ASAP7_75t_L g10210 ( 
.A(n_10187),
.Y(n_10210)
);

OA22x2_ASAP7_75t_L g10211 ( 
.A1(n_10174),
.A2(n_10178),
.B1(n_10162),
.B2(n_10177),
.Y(n_10211)
);

INVx3_ASAP7_75t_L g10212 ( 
.A(n_10173),
.Y(n_10212)
);

AO22x2_ASAP7_75t_L g10213 ( 
.A1(n_10190),
.A2(n_5358),
.B1(n_5366),
.B2(n_5356),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_10189),
.Y(n_10214)
);

OAI22xp5_ASAP7_75t_L g10215 ( 
.A1(n_10195),
.A2(n_3888),
.B1(n_3912),
.B2(n_3788),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_10193),
.Y(n_10216)
);

INVx2_ASAP7_75t_L g10217 ( 
.A(n_10191),
.Y(n_10217)
);

INVx2_ASAP7_75t_L g10218 ( 
.A(n_10211),
.Y(n_10218)
);

AOI22xp5_ASAP7_75t_L g10219 ( 
.A1(n_10196),
.A2(n_3985),
.B1(n_4005),
.B2(n_3965),
.Y(n_10219)
);

XOR2x1_ASAP7_75t_L g10220 ( 
.A(n_10202),
.B(n_4095),
.Y(n_10220)
);

INVx1_ASAP7_75t_L g10221 ( 
.A(n_10206),
.Y(n_10221)
);

XNOR2xp5_ASAP7_75t_L g10222 ( 
.A(n_10205),
.B(n_4133),
.Y(n_10222)
);

INVx1_ASAP7_75t_L g10223 ( 
.A(n_10194),
.Y(n_10223)
);

AOI22xp5_ASAP7_75t_L g10224 ( 
.A1(n_10192),
.A2(n_4005),
.B1(n_4008),
.B2(n_3965),
.Y(n_10224)
);

AND3x1_ASAP7_75t_L g10225 ( 
.A(n_10210),
.B(n_10212),
.C(n_10188),
.Y(n_10225)
);

INVx1_ASAP7_75t_L g10226 ( 
.A(n_10199),
.Y(n_10226)
);

AOI22x1_ASAP7_75t_L g10227 ( 
.A1(n_10197),
.A2(n_4025),
.B1(n_4061),
.B2(n_4008),
.Y(n_10227)
);

INVx1_ASAP7_75t_L g10228 ( 
.A(n_10198),
.Y(n_10228)
);

INVxp67_ASAP7_75t_L g10229 ( 
.A(n_10208),
.Y(n_10229)
);

INVx1_ASAP7_75t_L g10230 ( 
.A(n_10203),
.Y(n_10230)
);

INVx2_ASAP7_75t_L g10231 ( 
.A(n_10201),
.Y(n_10231)
);

AOI22xp5_ASAP7_75t_L g10232 ( 
.A1(n_10207),
.A2(n_4025),
.B1(n_4061),
.B2(n_4008),
.Y(n_10232)
);

INVx1_ASAP7_75t_L g10233 ( 
.A(n_10200),
.Y(n_10233)
);

INVx2_ASAP7_75t_L g10234 ( 
.A(n_10204),
.Y(n_10234)
);

NOR2x1p5_ASAP7_75t_L g10235 ( 
.A(n_10209),
.B(n_4025),
.Y(n_10235)
);

OA22x2_ASAP7_75t_L g10236 ( 
.A1(n_10214),
.A2(n_5358),
.B1(n_5366),
.B2(n_5356),
.Y(n_10236)
);

INVx1_ASAP7_75t_L g10237 ( 
.A(n_10218),
.Y(n_10237)
);

INVxp67_ASAP7_75t_SL g10238 ( 
.A(n_10221),
.Y(n_10238)
);

HB1xp67_ASAP7_75t_L g10239 ( 
.A(n_10217),
.Y(n_10239)
);

HB1xp67_ASAP7_75t_L g10240 ( 
.A(n_10216),
.Y(n_10240)
);

AOI21xp5_ASAP7_75t_L g10241 ( 
.A1(n_10223),
.A2(n_4246),
.B(n_4500),
.Y(n_10241)
);

CKINVDCx20_ASAP7_75t_R g10242 ( 
.A(n_10229),
.Y(n_10242)
);

AOI22xp5_ASAP7_75t_L g10243 ( 
.A1(n_10225),
.A2(n_4061),
.B1(n_4138),
.B2(n_3888),
.Y(n_10243)
);

INVx1_ASAP7_75t_L g10244 ( 
.A(n_10234),
.Y(n_10244)
);

A2O1A1Ixp33_ASAP7_75t_L g10245 ( 
.A1(n_10231),
.A2(n_5311),
.B(n_5316),
.C(n_5300),
.Y(n_10245)
);

NOR2xp33_ASAP7_75t_SL g10246 ( 
.A(n_10233),
.B(n_4080),
.Y(n_10246)
);

HB1xp67_ASAP7_75t_L g10247 ( 
.A(n_10226),
.Y(n_10247)
);

NAND3x1_ASAP7_75t_L g10248 ( 
.A(n_10230),
.B(n_10228),
.C(n_10224),
.Y(n_10248)
);

OAI22x1_ASAP7_75t_L g10249 ( 
.A1(n_10222),
.A2(n_4081),
.B1(n_3938),
.B2(n_3966),
.Y(n_10249)
);

INVx2_ASAP7_75t_L g10250 ( 
.A(n_10235),
.Y(n_10250)
);

INVx1_ASAP7_75t_L g10251 ( 
.A(n_10240),
.Y(n_10251)
);

INVx1_ASAP7_75t_L g10252 ( 
.A(n_10239),
.Y(n_10252)
);

INVx1_ASAP7_75t_L g10253 ( 
.A(n_10238),
.Y(n_10253)
);

INVx1_ASAP7_75t_L g10254 ( 
.A(n_10237),
.Y(n_10254)
);

INVx1_ASAP7_75t_L g10255 ( 
.A(n_10247),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_10244),
.Y(n_10256)
);

INVx2_ASAP7_75t_L g10257 ( 
.A(n_10242),
.Y(n_10257)
);

INVx1_ASAP7_75t_L g10258 ( 
.A(n_10246),
.Y(n_10258)
);

INVx1_ASAP7_75t_L g10259 ( 
.A(n_10250),
.Y(n_10259)
);

INVx1_ASAP7_75t_L g10260 ( 
.A(n_10248),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_10243),
.Y(n_10261)
);

INVx1_ASAP7_75t_L g10262 ( 
.A(n_10249),
.Y(n_10262)
);

INVx1_ASAP7_75t_L g10263 ( 
.A(n_10255),
.Y(n_10263)
);

BUFx2_ASAP7_75t_L g10264 ( 
.A(n_10251),
.Y(n_10264)
);

INVx2_ASAP7_75t_L g10265 ( 
.A(n_10257),
.Y(n_10265)
);

OAI21xp5_ASAP7_75t_L g10266 ( 
.A1(n_10256),
.A2(n_10215),
.B(n_10227),
.Y(n_10266)
);

AOI221x1_ASAP7_75t_L g10267 ( 
.A1(n_10260),
.A2(n_10241),
.B1(n_10213),
.B2(n_10245),
.C(n_10220),
.Y(n_10267)
);

OR3x2_ASAP7_75t_L g10268 ( 
.A(n_10254),
.B(n_10219),
.C(n_10232),
.Y(n_10268)
);

AOI22xp33_ASAP7_75t_L g10269 ( 
.A1(n_10264),
.A2(n_10252),
.B1(n_10253),
.B2(n_10259),
.Y(n_10269)
);

INVx1_ASAP7_75t_L g10270 ( 
.A(n_10263),
.Y(n_10270)
);

NAND2xp5_ASAP7_75t_SL g10271 ( 
.A(n_10265),
.B(n_10258),
.Y(n_10271)
);

AOI22xp5_ASAP7_75t_L g10272 ( 
.A1(n_10268),
.A2(n_10261),
.B1(n_10262),
.B2(n_10236),
.Y(n_10272)
);

AOI22x1_ASAP7_75t_L g10273 ( 
.A1(n_10270),
.A2(n_10266),
.B1(n_10267),
.B2(n_4087),
.Y(n_10273)
);

OAI22xp5_ASAP7_75t_SL g10274 ( 
.A1(n_10269),
.A2(n_4087),
.B1(n_4113),
.B2(n_4080),
.Y(n_10274)
);

AOI21xp5_ASAP7_75t_L g10275 ( 
.A1(n_10273),
.A2(n_10271),
.B(n_10272),
.Y(n_10275)
);

AOI22xp5_ASAP7_75t_SL g10276 ( 
.A1(n_10275),
.A2(n_10274),
.B1(n_4069),
.B2(n_4056),
.Y(n_10276)
);

INVx1_ASAP7_75t_L g10277 ( 
.A(n_10276),
.Y(n_10277)
);

AO221x2_ASAP7_75t_L g10278 ( 
.A1(n_10277),
.A2(n_5316),
.B1(n_5335),
.B2(n_5329),
.C(n_5311),
.Y(n_10278)
);

AOI221xp5_ASAP7_75t_L g10279 ( 
.A1(n_10278),
.A2(n_5340),
.B1(n_5348),
.B2(n_5335),
.C(n_5329),
.Y(n_10279)
);

AOI21xp33_ASAP7_75t_L g10280 ( 
.A1(n_10279),
.A2(n_3878),
.B(n_3864),
.Y(n_10280)
);

AOI211xp5_ASAP7_75t_L g10281 ( 
.A1(n_10280),
.A2(n_3938),
.B(n_3966),
.C(n_3920),
.Y(n_10281)
);


endmodule