module fake_jpeg_28892_n_478 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_478);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_478;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_47),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_53),
.Y(n_121)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_54),
.B(n_72),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_21),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_55),
.Y(n_141)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_8),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_78),
.Y(n_140)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_76),
.B(n_77),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_82),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_29),
.B(n_8),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_36),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_9),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_17),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_9),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_93),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_30),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_46),
.B1(n_39),
.B2(n_23),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_95),
.A2(n_98),
.B1(n_115),
.B2(n_116),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_55),
.B1(n_47),
.B2(n_46),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_46),
.B1(n_25),
.B2(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_103),
.A2(n_120),
.B1(n_125),
.B2(n_127),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_65),
.A2(n_25),
.B1(n_44),
.B2(n_31),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_47),
.A2(n_94),
.B1(n_85),
.B2(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_52),
.A2(n_18),
.B1(n_44),
.B2(n_34),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_145),
.B1(n_58),
.B2(n_20),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_45),
.B1(n_41),
.B2(n_16),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_59),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_24),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_85),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_50),
.B1(n_92),
.B2(n_91),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_150),
.A2(n_172),
.B1(n_181),
.B2(n_110),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_154),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_93),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_18),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_168),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_64),
.B(n_58),
.C(n_24),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_163),
.B(n_176),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_66),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_169),
.Y(n_207)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_130),
.A2(n_53),
.B1(n_22),
.B2(n_56),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_86),
.C(n_63),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_106),
.C(n_139),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_90),
.B1(n_51),
.B2(n_57),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_69),
.B1(n_71),
.B2(n_87),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_49),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_79),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_183),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_134),
.A2(n_74),
.B1(n_75),
.B2(n_81),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_193),
.B1(n_116),
.B2(n_145),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_24),
.B1(n_60),
.B2(n_37),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_191),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_115),
.A2(n_37),
.B1(n_10),
.B2(n_11),
.Y(n_181)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_104),
.B(n_7),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_37),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_185),
.Y(n_215)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_7),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_37),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_141),
.Y(n_191)
);

BUFx24_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_108),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_198),
.B(n_136),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_114),
.B(n_135),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_206),
.B(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_202),
.A2(n_180),
.B1(n_175),
.B2(n_191),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_138),
.B(n_107),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_160),
.B1(n_151),
.B2(n_192),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_165),
.B1(n_194),
.B2(n_154),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_171),
.B1(n_156),
.B2(n_153),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_143),
.B1(n_146),
.B2(n_148),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_231),
.B1(n_103),
.B2(n_95),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_164),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_114),
.B(n_139),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_172),
.A2(n_181),
.B1(n_150),
.B2(n_176),
.Y(n_231)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_241),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_SL g237 ( 
.A1(n_229),
.A2(n_183),
.B(n_163),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_238),
.B1(n_245),
.B2(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_240),
.A2(n_206),
.B1(n_207),
.B2(n_197),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_177),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_165),
.B(n_157),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_243),
.A2(n_207),
.B(n_215),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_158),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_251),
.Y(n_280)
);

OR2x2_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_180),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_227),
.B1(n_219),
.B2(n_202),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_218),
.B1(n_224),
.B2(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_152),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_180),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_262),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_168),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_219),
.C(n_227),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_123),
.B1(n_117),
.B2(n_111),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_255),
.A2(n_259),
.B1(n_261),
.B2(n_155),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_195),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_260),
.Y(n_299)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_212),
.A2(n_146),
.B1(n_148),
.B2(n_110),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_196),
.A2(n_108),
.B1(n_123),
.B2(n_117),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_201),
.B(n_159),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_201),
.B(n_159),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_266),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_211),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_167),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_198),
.B(n_188),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_210),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_147),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_281),
.B1(n_292),
.B2(n_293),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_273),
.A2(n_278),
.B(n_284),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_208),
.C(n_215),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_277),
.B(n_286),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_200),
.B(n_208),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_227),
.B(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_238),
.B1(n_245),
.B2(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_289),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_227),
.B1(n_205),
.B2(n_204),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_228),
.B1(n_232),
.B2(n_205),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_243),
.A2(n_175),
.B(n_226),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_256),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_265),
.A2(n_232),
.B1(n_210),
.B2(n_226),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_259),
.A2(n_251),
.B1(n_249),
.B2(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_297),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_214),
.C(n_220),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_256),
.C(n_247),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_257),
.Y(n_297)
);

OAI22x1_ASAP7_75t_SL g298 ( 
.A1(n_240),
.A2(n_164),
.B1(n_166),
.B2(n_155),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_298),
.A2(n_261),
.B1(n_242),
.B2(n_248),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_270),
.B(n_241),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_303),
.B(n_308),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_300),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_309),
.C(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_276),
.B(n_257),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_286),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_246),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_294),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_313),
.Y(n_340)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_284),
.B(n_290),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx3_ASAP7_75t_SL g317 ( 
.A(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_318),
.A2(n_289),
.B1(n_271),
.B2(n_285),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_279),
.B(n_263),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_319),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_321),
.C(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_236),
.C(n_262),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_280),
.B(n_258),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_291),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_280),
.B(n_252),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_260),
.C(n_239),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_235),
.Y(n_328)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_234),
.Y(n_329)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_291),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_332),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_275),
.C(n_299),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_339),
.C(n_361),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_345),
.Y(n_382)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_299),
.C(n_287),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_271),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_323),
.B(n_305),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_350),
.A2(n_355),
.B1(n_331),
.B2(n_301),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_302),
.Y(n_354)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_305),
.A2(n_278),
.B1(n_273),
.B2(n_283),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_272),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_312),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_301),
.A2(n_272),
.B1(n_221),
.B2(n_209),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_317),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_214),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_380),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_334),
.A2(n_317),
.B(n_323),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_366),
.B(n_369),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_387),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_340),
.B(n_313),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_308),
.Y(n_370)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_335),
.C(n_357),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_386),
.C(n_339),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_377),
.A2(n_334),
.B1(n_362),
.B2(n_349),
.Y(n_390)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_321),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_379),
.B(n_355),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_314),
.Y(n_380)
);

AOI21x1_ASAP7_75t_SL g383 ( 
.A1(n_347),
.A2(n_318),
.B(n_330),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_384),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_342),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_388),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_333),
.B(n_327),
.C(n_331),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_307),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_306),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_400),
.Y(n_413)
);

XOR2x2_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_345),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_366),
.C(n_347),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_336),
.Y(n_397)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_384),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_364),
.C(n_374),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_407),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_361),
.C(n_337),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_406),
.C(n_408),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_362),
.C(n_350),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_386),
.B(n_349),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_358),
.C(n_352),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_372),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_405),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_401),
.A2(n_365),
.B(n_368),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_412),
.A2(n_423),
.B(n_220),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_422),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_382),
.C(n_367),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_417),
.C(n_419),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_382),
.C(n_380),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_391),
.B(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_424),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_381),
.C(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_420),
.B(n_389),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_SL g421 ( 
.A1(n_392),
.A2(n_371),
.B(n_374),
.C(n_360),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_421),
.A2(n_399),
.B1(n_394),
.B2(n_409),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_376),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_392),
.A2(n_396),
.B(n_398),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_396),
.A2(n_385),
.B1(n_358),
.B2(n_343),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_363),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_413),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_426),
.A2(n_399),
.B1(n_398),
.B2(n_405),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_427),
.A2(n_441),
.B1(n_209),
.B2(n_170),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_363),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_433),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_389),
.C(n_395),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_416),
.C(n_421),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_394),
.Y(n_434)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_435),
.B(n_438),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_437),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_221),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_439),
.B(n_440),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_421),
.A2(n_422),
.B1(n_414),
.B2(n_410),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_421),
.A2(n_221),
.B1(n_209),
.B2(n_233),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_410),
.B(n_185),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_442),
.B(n_6),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_444),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_174),
.C(n_186),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_449),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_187),
.C(n_147),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_182),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_454),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_440),
.A2(n_138),
.B(n_7),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_452),
.A2(n_447),
.B(n_437),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_434),
.A2(n_6),
.B(n_14),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_453),
.A2(n_430),
.B(n_14),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_456),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_443),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_464),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_452),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g460 ( 
.A1(n_455),
.A2(n_432),
.B(n_431),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_463),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_450),
.A2(n_445),
.B(n_446),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_432),
.B(n_138),
.Y(n_464)
);

MAJx2_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_449),
.C(n_462),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_457),
.C(n_10),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_466),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_5),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_470),
.A2(n_14),
.B(n_5),
.Y(n_473)
);

AOI221xp5_ASAP7_75t_L g474 ( 
.A1(n_472),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.C(n_10),
.Y(n_474)
);

OAI321xp33_ASAP7_75t_L g475 ( 
.A1(n_473),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_12),
.C(n_471),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_474),
.A2(n_475),
.B(n_12),
.Y(n_476)
);

OAI211xp5_ASAP7_75t_L g477 ( 
.A1(n_476),
.A2(n_0),
.B(n_1),
.C(n_369),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_1),
.Y(n_478)
);


endmodule