module real_jpeg_31820_n_11 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_107, n_6, n_104, n_106, n_110, n_112, n_7, n_3, n_5, n_4, n_105, n_109, n_1, n_113, n_11);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_107;
input n_6;
input n_104;
input n_106;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_105;
input n_109;
input n_1;
input n_113;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_0),
.B(n_42),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_1),
.B(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_2),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI221xp5_ASAP7_75t_L g56 ( 
.A1(n_4),
.A2(n_9),
.B1(n_57),
.B2(n_63),
.C(n_65),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_5),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_57),
.C(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_10),
.B(n_90),
.Y(n_89)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_10),
.B(n_95),
.CON(n_94),
.SN(n_94)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_20),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_104),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_98),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_24),
.Y(n_54)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B(n_96),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_89),
.B(n_94),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_47),
.B(n_87),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_78),
.C(n_79),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_69),
.B(n_77),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_56),
.B1(n_67),
.B2(n_68),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_110),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_94),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_105),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_106),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_107),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_108),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_109),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_111),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_112),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_113),
.Y(n_91)
);


endmodule