module fake_jpeg_23929_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_0),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_47),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_57),
.B(n_29),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_18),
.B1(n_33),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_62),
.B1(n_29),
.B2(n_26),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_26),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_39),
.C(n_38),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_72),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_32),
.B1(n_30),
.B2(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_13),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_11),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_78),
.Y(n_106)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_45),
.B1(n_39),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_63),
.B1(n_4),
.B2(n_3),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_27),
.B(n_26),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_89),
.B(n_90),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_69),
.B(n_66),
.C(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_2),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_92),
.C(n_102),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_9),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_38),
.B(n_9),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_6),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_15),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_15),
.B1(n_63),
.B2(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_78),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_6),
.B(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_103),
.B(n_109),
.Y(n_146)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_70),
.B(n_46),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_118),
.B1(n_120),
.B2(n_124),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_117),
.Y(n_136)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_119),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_46),
.A3(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_129),
.A2(n_85),
.B1(n_77),
.B2(n_76),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_135),
.B1(n_145),
.B2(n_108),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_83),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_118),
.B(n_123),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_81),
.B1(n_79),
.B2(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_90),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_93),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_84),
.B1(n_75),
.B2(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_108),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_157),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_127),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_158),
.C(n_159),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_113),
.B(n_104),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_170),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_107),
.C(n_125),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_147),
.B(n_132),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_161),
.B(n_162),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_139),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_137),
.B1(n_134),
.B2(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_178),
.B(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_179),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_138),
.B(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_159),
.C(n_160),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.C(n_190),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_155),
.C(n_153),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_174),
.A2(n_165),
.B1(n_166),
.B2(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_178),
.C(n_153),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_158),
.C(n_140),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_181),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_183),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_203),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_174),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

AOI21x1_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_141),
.B(n_142),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_142),
.B1(n_190),
.B2(n_186),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_194),
.B(n_169),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_204),
.B1(n_197),
.B2(n_187),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_207),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_206),
.B(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.C(n_209),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_201),
.C(n_207),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_214),
.A3(n_177),
.B1(n_157),
.B2(n_198),
.C1(n_139),
.C2(n_137),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_218),
.B(n_143),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_146),
.Y(n_222)
);


endmodule