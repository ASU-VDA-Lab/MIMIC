module fake_jpeg_306_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_38),
.B(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_31),
.Y(n_54)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_31),
.B1(n_28),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_49),
.B1(n_48),
.B2(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_29),
.B1(n_26),
.B2(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_20),
.B1(n_28),
.B2(n_17),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_89),
.B1(n_99),
.B2(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_92),
.Y(n_104)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_22),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_23),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_96),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_50),
.C(n_40),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_53),
.C(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_118),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_24),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_43),
.B1(n_61),
.B2(n_45),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_61),
.B1(n_68),
.B2(n_24),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_59),
.B1(n_51),
.B2(n_20),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_51),
.B(n_59),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_93),
.B(n_81),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_18),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_7),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_132),
.B1(n_141),
.B2(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_102),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_129),
.B(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_100),
.B1(n_98),
.B2(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_118),
.B(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_90),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_94),
.B1(n_91),
.B2(n_80),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_155),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_145),
.B1(n_147),
.B2(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_137),
.B1(n_138),
.B2(n_135),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_147),
.B(n_149),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_108),
.B1(n_119),
.B2(n_120),
.C(n_116),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_118),
.B1(n_103),
.B2(n_110),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_153),
.B(n_18),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_105),
.B(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_R g154 ( 
.A(n_126),
.B(n_21),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_146),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_131),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_159),
.C(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_130),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_141),
.B1(n_140),
.B2(n_134),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_164),
.B(n_166),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_136),
.B(n_2),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_21),
.B1(n_18),
.B2(n_3),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_161),
.B1(n_167),
.B2(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_175),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_152),
.C(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_166),
.C(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_162),
.B(n_153),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_181),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_18),
.B(n_10),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_6),
.C(n_13),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_169),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_12),
.B1(n_15),
.B2(n_4),
.Y(n_188)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_10),
.B(n_13),
.C(n_12),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_1),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_186),
.Y(n_191)
);

OAI211xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_185),
.B(n_4),
.C(n_5),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_190),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_2),
.Y(n_194)
);


endmodule