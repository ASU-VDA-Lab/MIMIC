module real_aes_8140_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_140;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g543 ( .A1(n_0), .A2(n_160), .B(n_544), .C(n_547), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_1), .B(n_494), .Y(n_548) );
INVx1_ASAP7_75t_L g420 ( .A(n_2), .Y(n_420) );
INVx1_ASAP7_75t_L g172 ( .A(n_3), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_4), .B(n_132), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_5), .A2(n_467), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_6), .A2(n_152), .B(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_7), .A2(n_38), .B1(n_126), .B2(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_8), .B(n_152), .Y(n_161) );
AND2x6_ASAP7_75t_L g144 ( .A(n_9), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_10), .A2(n_144), .B(n_472), .C(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_11), .B(n_39), .Y(n_421) );
INVx1_ASAP7_75t_L g122 ( .A(n_12), .Y(n_122) );
INVx1_ASAP7_75t_L g165 ( .A(n_13), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_14), .B(n_130), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_15), .B(n_132), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_16), .B(n_118), .Y(n_236) );
AO32x2_ASAP7_75t_L g178 ( .A1(n_17), .A2(n_117), .A3(n_143), .B1(n_152), .B2(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_18), .B(n_126), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_19), .B(n_118), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_20), .A2(n_54), .B1(n_126), .B2(n_181), .Y(n_182) );
AOI22xp33_ASAP7_75t_SL g220 ( .A1(n_21), .A2(n_81), .B1(n_126), .B2(n_130), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_22), .B(n_126), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_23), .A2(n_143), .B(n_472), .C(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_24), .A2(n_60), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_24), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_25), .A2(n_143), .B(n_472), .C(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_26), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_27), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_28), .B(n_426), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_29), .A2(n_467), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_30), .B(n_147), .Y(n_195) );
INVx2_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_32), .A2(n_470), .B(n_480), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_33), .B(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_34), .B(n_147), .Y(n_206) );
XNOR2x2_ASAP7_75t_SL g105 ( .A(n_35), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_36), .B(n_202), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_37), .A2(n_85), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_37), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_40), .B(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_41), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_42), .B(n_132), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_43), .B(n_467), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_44), .A2(n_470), .B(n_474), .C(n_480), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_45), .A2(n_104), .B1(n_429), .B2(n_438), .C(n_441), .Y(n_103) );
OAI321xp33_ASAP7_75t_L g104 ( .A1(n_45), .A2(n_105), .A3(n_414), .B1(n_422), .B2(n_423), .C(n_425), .Y(n_104) );
INVx1_ASAP7_75t_L g422 ( .A(n_45), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_46), .B(n_126), .Y(n_155) );
INVx1_ASAP7_75t_L g545 ( .A(n_47), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_48), .A2(n_90), .B1(n_181), .B2(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g475 ( .A(n_49), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_50), .B(n_126), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_51), .B(n_126), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_52), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_53), .B(n_138), .Y(n_159) );
AOI22xp33_ASAP7_75t_SL g234 ( .A1(n_55), .A2(n_61), .B1(n_126), .B2(n_130), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_56), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_57), .B(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_58), .B(n_126), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_59), .B(n_126), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_60), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_60), .A2(n_109), .B1(n_110), .B2(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g145 ( .A(n_62), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_63), .B(n_467), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_64), .B(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_65), .A2(n_138), .B(n_168), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_66), .B(n_126), .Y(n_173) );
INVx1_ASAP7_75t_L g121 ( .A(n_67), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_68), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_69), .B(n_132), .Y(n_512) );
AO32x2_ASAP7_75t_L g216 ( .A1(n_70), .A2(n_143), .A3(n_152), .B1(n_217), .B2(n_221), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_71), .B(n_133), .Y(n_558) );
INVx1_ASAP7_75t_L g136 ( .A(n_72), .Y(n_136) );
INVx1_ASAP7_75t_L g190 ( .A(n_73), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_74), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_75), .B(n_477), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_76), .A2(n_472), .B(n_480), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_77), .B(n_130), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_78), .Y(n_489) );
INVx1_ASAP7_75t_L g437 ( .A(n_79), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_80), .B(n_476), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_82), .B(n_181), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_83), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_84), .B(n_130), .Y(n_194) );
INVx1_ASAP7_75t_L g449 ( .A(n_85), .Y(n_449) );
INVx2_ASAP7_75t_L g119 ( .A(n_86), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_87), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_88), .B(n_142), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_89), .B(n_130), .Y(n_156) );
OR2x2_ASAP7_75t_L g417 ( .A(n_91), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g453 ( .A(n_91), .B(n_419), .Y(n_453) );
INVx2_ASAP7_75t_L g459 ( .A(n_91), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_92), .A2(n_102), .B1(n_130), .B2(n_131), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_93), .B(n_467), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_94), .Y(n_511) );
INVxp67_ASAP7_75t_L g492 ( .A(n_95), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_96), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_97), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g533 ( .A(n_98), .Y(n_533) );
INVx1_ASAP7_75t_L g554 ( .A(n_99), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_100), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_100), .Y(n_445) );
AND2x2_ASAP7_75t_L g482 ( .A(n_101), .B(n_147), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_105), .B(n_424), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_SL g455 ( .A(n_110), .Y(n_455) );
OR3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_342), .C(n_391), .Y(n_110) );
NAND5xp2_ASAP7_75t_L g111 ( .A(n_112), .B(n_257), .C(n_285), .D(n_315), .E(n_329), .Y(n_111) );
AOI221xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_175), .B1(n_207), .B2(n_212), .C(n_223), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_148), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_114), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g237 ( .A(n_115), .Y(n_237) );
AND2x2_ASAP7_75t_L g245 ( .A(n_115), .B(n_151), .Y(n_245) );
AND2x2_ASAP7_75t_L g268 ( .A(n_115), .B(n_150), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_115), .B(n_162), .Y(n_283) );
OR2x2_ASAP7_75t_L g292 ( .A(n_115), .B(n_230), .Y(n_292) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_115), .Y(n_295) );
AND2x2_ASAP7_75t_L g403 ( .A(n_115), .B(n_230), .Y(n_403) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_123), .B(n_146), .Y(n_115) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_116), .A2(n_163), .B(n_174), .Y(n_162) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_117), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_119), .B(n_120), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_135), .B(n_143), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_132), .Y(n_124) );
INVx3_ASAP7_75t_L g189 ( .A(n_126), .Y(n_189) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_126), .Y(n_535) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
BUFx3_ASAP7_75t_L g219 ( .A(n_127), .Y(n_219) );
AND2x6_ASAP7_75t_L g472 ( .A(n_127), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
INVx1_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
INVx2_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_132), .A2(n_155), .B(n_156), .Y(n_154) );
INVx2_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_SL g188 ( .A1(n_132), .A2(n_189), .B(n_190), .C(n_191), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_132), .B(n_492), .Y(n_491) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g217 ( .A1(n_133), .A2(n_142), .B1(n_218), .B2(n_220), .Y(n_217) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_134), .Y(n_170) );
INVx1_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
AND2x2_ASAP7_75t_L g468 ( .A(n_134), .B(n_139), .Y(n_468) );
INVx1_ASAP7_75t_L g473 ( .A(n_134), .Y(n_473) );
O2A1O1Ixp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_140), .C(n_141), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_137), .A2(n_160), .B(n_172), .C(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_137), .A2(n_522), .B(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_141), .A2(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_142), .A2(n_160), .B1(n_180), .B2(n_182), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_142), .A2(n_160), .B1(n_233), .B2(n_234), .Y(n_232) );
INVx4_ASAP7_75t_L g546 ( .A(n_142), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_143), .B(n_231), .C(n_232), .Y(n_256) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_144), .A2(n_154), .B(n_157), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_144), .A2(n_164), .B(n_171), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_144), .A2(n_188), .B(n_192), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_144), .A2(n_198), .B(n_203), .Y(n_197) );
AND2x4_ASAP7_75t_L g467 ( .A(n_144), .B(n_468), .Y(n_467) );
INVx4_ASAP7_75t_SL g481 ( .A(n_144), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_144), .B(n_468), .Y(n_555) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_147), .A2(n_187), .B(n_195), .Y(n_186) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_147), .A2(n_197), .B(n_206), .Y(n_196) );
INVx2_ASAP7_75t_L g221 ( .A(n_147), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_147), .A2(n_466), .B(n_469), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_147), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g527 ( .A(n_147), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_148), .B(n_295), .Y(n_351) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
OAI311xp33_ASAP7_75t_L g293 ( .A1(n_149), .A2(n_294), .A3(n_295), .B1(n_296), .C1(n_311), .Y(n_293) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_162), .Y(n_149) );
AND2x2_ASAP7_75t_L g254 ( .A(n_150), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g261 ( .A(n_150), .Y(n_261) );
AND2x2_ASAP7_75t_L g382 ( .A(n_150), .B(n_211), .Y(n_382) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_151), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g238 ( .A(n_151), .B(n_162), .Y(n_238) );
AND2x2_ASAP7_75t_L g290 ( .A(n_151), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g304 ( .A(n_151), .B(n_237), .Y(n_304) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_161), .Y(n_151) );
INVx4_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_152), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_152), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_160), .Y(n_157) );
INVx2_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
AND2x2_ASAP7_75t_L g253 ( .A(n_162), .B(n_237), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_168), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_166), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_166), .A2(n_558), .B(n_559), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_168), .A2(n_533), .B(n_534), .C(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_169), .A2(n_193), .B(n_194), .Y(n_192) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g477 ( .A(n_170), .Y(n_477) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_183), .Y(n_175) );
OR2x2_ASAP7_75t_L g348 ( .A(n_176), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_176), .B(n_354), .Y(n_365) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_177), .B(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g222 ( .A(n_178), .Y(n_222) );
AND2x2_ASAP7_75t_L g289 ( .A(n_178), .B(n_216), .Y(n_289) );
AND2x2_ASAP7_75t_L g300 ( .A(n_178), .B(n_196), .Y(n_300) );
AND2x2_ASAP7_75t_L g309 ( .A(n_178), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_183), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_183), .B(n_250), .Y(n_294) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g281 ( .A(n_184), .B(n_240), .Y(n_281) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_196), .Y(n_184) );
INVx2_ASAP7_75t_L g214 ( .A(n_185), .Y(n_214) );
AND2x2_ASAP7_75t_L g308 ( .A(n_185), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g226 ( .A(n_186), .Y(n_226) );
OR2x2_ASAP7_75t_L g325 ( .A(n_186), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_186), .Y(n_388) );
AND2x2_ASAP7_75t_L g227 ( .A(n_196), .B(n_222), .Y(n_227) );
INVx1_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
AND2x2_ASAP7_75t_L g269 ( .A(n_196), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g310 ( .A(n_196), .Y(n_310) );
INVx1_ASAP7_75t_L g326 ( .A(n_196), .Y(n_326) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_196), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVxp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_209), .B(n_314), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_209), .A2(n_299), .B1(n_348), .B2(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_210), .A2(n_392), .B(n_394), .C(n_412), .Y(n_391) );
INVx2_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
AND2x2_ASAP7_75t_L g302 ( .A(n_211), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g313 ( .A(n_211), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_212), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_250), .Y(n_286) );
BUFx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g318 ( .A(n_214), .B(n_309), .Y(n_318) );
AND2x2_ASAP7_75t_L g337 ( .A(n_214), .B(n_251), .Y(n_337) );
AND2x4_ASAP7_75t_L g273 ( .A(n_215), .B(n_247), .Y(n_273) );
AND2x2_ASAP7_75t_L g411 ( .A(n_215), .B(n_387), .Y(n_411) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVx1_ASAP7_75t_L g251 ( .A(n_216), .Y(n_251) );
INVx1_ASAP7_75t_L g350 ( .A(n_216), .Y(n_350) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_219), .Y(n_479) );
INVx2_ASAP7_75t_L g547 ( .A(n_219), .Y(n_547) );
INVx1_ASAP7_75t_L g524 ( .A(n_221), .Y(n_524) );
OR2x2_ASAP7_75t_L g241 ( .A(n_222), .B(n_226), .Y(n_241) );
AND2x2_ASAP7_75t_L g250 ( .A(n_222), .B(n_251), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g270 ( .A(n_222), .B(n_271), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_228), .B1(n_239), .B2(n_242), .C(n_246), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_225), .A2(n_247), .B(n_249), .C(n_252), .Y(n_246) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g271 ( .A(n_226), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_226), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_226), .B(n_248), .Y(n_354) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_226), .Y(n_361) );
AND2x2_ASAP7_75t_L g279 ( .A(n_227), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g316 ( .A(n_227), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_238), .Y(n_228) );
INVx2_ASAP7_75t_L g307 ( .A(n_229), .Y(n_307) );
AOI222xp33_ASAP7_75t_L g356 ( .A1(n_229), .A2(n_240), .B1(n_357), .B2(n_359), .C1(n_360), .C2(n_362), .Y(n_356) );
AND2x2_ASAP7_75t_L g413 ( .A(n_229), .B(n_382), .Y(n_413) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_237), .Y(n_229) );
INVx1_ASAP7_75t_L g303 ( .A(n_230), .Y(n_303) );
AO21x1_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_235), .Y(n_230) );
INVx3_ASAP7_75t_L g494 ( .A(n_231), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_231), .B(n_514), .Y(n_513) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_231), .A2(n_530), .B(n_537), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_231), .B(n_538), .Y(n_537) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_231), .A2(n_553), .B(n_560), .Y(n_552) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g255 ( .A(n_236), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g341 ( .A(n_238), .B(n_275), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g352 ( .A1(n_239), .A2(n_353), .B(n_355), .Y(n_352) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g280 ( .A(n_240), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_240), .B(n_247), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_240), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx3_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
OR2x2_ASAP7_75t_L g358 ( .A(n_244), .B(n_280), .Y(n_358) );
AND2x2_ASAP7_75t_L g274 ( .A(n_245), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g312 ( .A(n_245), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_245), .B(n_306), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_245), .B(n_302), .Y(n_328) );
AND2x2_ASAP7_75t_L g332 ( .A(n_245), .B(n_314), .Y(n_332) );
INVxp67_ASAP7_75t_L g264 ( .A(n_247), .Y(n_264) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_249), .A2(n_322), .B1(n_327), .B2(n_328), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_249), .B(n_354), .Y(n_384) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g370 ( .A(n_250), .B(n_361), .Y(n_370) );
AND2x2_ASAP7_75t_L g399 ( .A(n_250), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g404 ( .A(n_250), .B(n_354), .Y(n_404) );
INVx1_ASAP7_75t_L g317 ( .A(n_251), .Y(n_317) );
BUFx2_ASAP7_75t_L g323 ( .A(n_251), .Y(n_323) );
INVx1_ASAP7_75t_L g408 ( .A(n_252), .Y(n_408) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_253), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_255), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g267 ( .A(n_255), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
INVx3_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
OR2x2_ASAP7_75t_L g380 ( .A(n_255), .B(n_381), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B(n_265), .C(n_277), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_258), .A2(n_395), .B1(n_402), .B2(n_404), .C(n_405), .Y(n_394) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_266), .B(n_272), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_268), .B(n_306), .Y(n_320) );
AND2x2_ASAP7_75t_L g362 ( .A(n_268), .B(n_302), .Y(n_362) );
INVx1_ASAP7_75t_SL g375 ( .A(n_269), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_269), .B(n_323), .Y(n_378) );
INVx1_ASAP7_75t_L g396 ( .A(n_270), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_274), .A2(n_364), .B1(n_366), .B2(n_370), .C(n_371), .Y(n_363) );
AND2x2_ASAP7_75t_L g390 ( .A(n_275), .B(n_382), .Y(n_390) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g374 ( .A(n_276), .Y(n_374) );
AOI21xp33_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_281), .B(n_282), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g345 ( .A(n_280), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g331 ( .A(n_281), .Y(n_331) );
INVx1_ASAP7_75t_L g359 ( .A(n_282), .Y(n_359) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_290), .C(n_293), .Y(n_285) );
OAI31xp33_ASAP7_75t_L g412 ( .A1(n_286), .A2(n_324), .A3(n_411), .B(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g386 ( .A(n_289), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g407 ( .A(n_289), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_291), .B(n_306), .Y(n_334) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g409 ( .A(n_292), .B(n_306), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_301), .B1(n_305), .B2(n_308), .Y(n_296) );
NAND2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_300), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g336 ( .A(n_300), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g339 ( .A(n_300), .B(n_323), .Y(n_339) );
AND2x2_ASAP7_75t_L g393 ( .A(n_300), .B(n_388), .Y(n_393) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g368 ( .A(n_304), .Y(n_368) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OAI32xp33_ASAP7_75t_L g371 ( .A1(n_306), .A2(n_340), .A3(n_372), .B1(n_374), .B2(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_309), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B(n_319), .C(n_321), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_317), .B(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_318), .A2(n_330), .B1(n_331), .B2(n_332), .C(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g330 ( .A(n_328), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_338), .B2(n_340), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND4xp25_ASAP7_75t_SL g395 ( .A(n_338), .B(n_396), .C(n_397), .D(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NAND4xp25_ASAP7_75t_SL g342 ( .A(n_343), .B(n_356), .C(n_363), .D(n_376), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_351), .C(n_352), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g373 ( .A(n_349), .Y(n_373) );
INVx2_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
OR2x2_ASAP7_75t_L g406 ( .A(n_361), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_383), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_382), .B(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g424 ( .A(n_416), .Y(n_424) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g428 ( .A(n_417), .Y(n_428) );
BUFx2_ASAP7_75t_L g440 ( .A(n_417), .Y(n_440) );
INVx1_ASAP7_75t_SL g770 ( .A(n_417), .Y(n_770) );
NOR2x2_ASAP7_75t_L g766 ( .A(n_418), .B(n_459), .Y(n_766) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g458 ( .A(n_419), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_434), .A2(n_435), .B(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g768 ( .A(n_434), .B(n_436), .Y(n_768) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_763), .B(n_767), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_450), .B2(n_758), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B1(n_456), .B2(n_460), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g759 ( .A(n_452), .Y(n_759) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g760 ( .A(n_454), .Y(n_760) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g761 ( .A(n_457), .Y(n_761) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx4_ASAP7_75t_L g762 ( .A(n_460), .Y(n_762) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR5x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_631), .C(n_709), .D(n_733), .E(n_750), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_503), .B(n_549), .C(n_608), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_483), .Y(n_463) );
AND2x2_ASAP7_75t_L g562 ( .A(n_464), .B(n_485), .Y(n_562) );
INVx5_ASAP7_75t_SL g590 ( .A(n_464), .Y(n_590) );
AND2x2_ASAP7_75t_L g626 ( .A(n_464), .B(n_611), .Y(n_626) );
OR2x2_ASAP7_75t_L g665 ( .A(n_464), .B(n_484), .Y(n_665) );
OR2x2_ASAP7_75t_L g696 ( .A(n_464), .B(n_587), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_464), .B(n_600), .Y(n_732) );
AND2x2_ASAP7_75t_L g744 ( .A(n_464), .B(n_587), .Y(n_744) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_482), .Y(n_464) );
BUFx2_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_471), .A2(n_481), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g541 ( .A1(n_471), .A2(n_481), .B(n_542), .C(n_543), .Y(n_541) );
INVx5_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_478), .C(n_479), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_476), .A2(n_479), .B(n_511), .C(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g743 ( .A(n_483), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g606 ( .A(n_484), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_485), .B(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_485), .Y(n_599) );
INVx3_ASAP7_75t_L g614 ( .A(n_485), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_485), .B(n_495), .Y(n_638) );
OR2x2_ASAP7_75t_L g647 ( .A(n_485), .B(n_590), .Y(n_647) );
AND2x2_ASAP7_75t_L g651 ( .A(n_485), .B(n_611), .Y(n_651) );
AND2x2_ASAP7_75t_L g657 ( .A(n_485), .B(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g694 ( .A(n_485), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_485), .B(n_552), .Y(n_708) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_493), .Y(n_485) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_494), .A2(n_540), .B(n_548), .Y(n_539) );
OR2x2_ASAP7_75t_L g600 ( .A(n_495), .B(n_552), .Y(n_600) );
AND2x2_ASAP7_75t_L g611 ( .A(n_495), .B(n_587), .Y(n_611) );
AND2x2_ASAP7_75t_L g623 ( .A(n_495), .B(n_614), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_495), .B(n_552), .Y(n_646) );
INVx1_ASAP7_75t_SL g658 ( .A(n_495), .Y(n_658) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g551 ( .A(n_496), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_496), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_515), .Y(n_504) );
AND2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_505), .B(n_528), .Y(n_575) );
AND2x2_ASAP7_75t_L g578 ( .A(n_505), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_505), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g603 ( .A(n_505), .B(n_594), .Y(n_603) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_505), .Y(n_622) );
AND2x2_ASAP7_75t_L g643 ( .A(n_505), .B(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g653 ( .A(n_505), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g699 ( .A(n_505), .B(n_582), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_505), .B(n_605), .Y(n_726) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g596 ( .A(n_506), .Y(n_596) );
AND2x2_ASAP7_75t_L g662 ( .A(n_506), .B(n_594), .Y(n_662) );
AND2x2_ASAP7_75t_L g746 ( .A(n_506), .B(n_614), .Y(n_746) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_515), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_515), .Y(n_735) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_528), .Y(n_515) );
AND2x2_ASAP7_75t_L g565 ( .A(n_516), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g574 ( .A(n_516), .B(n_572), .Y(n_574) );
INVx5_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
AND2x2_ASAP7_75t_L g605 ( .A(n_516), .B(n_539), .Y(n_605) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_516), .Y(n_642) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
AOI21xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_520), .B(n_524), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g683 ( .A(n_528), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_528), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g716 ( .A(n_528), .B(n_582), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g745 ( .A1(n_528), .A2(n_639), .B(n_746), .C(n_747), .Y(n_745) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
BUFx2_ASAP7_75t_L g566 ( .A(n_529), .Y(n_566) );
INVx2_ASAP7_75t_L g570 ( .A(n_529), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
INVx2_ASAP7_75t_L g572 ( .A(n_539), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_539), .B(n_570), .Y(n_579) );
AND2x2_ASAP7_75t_L g670 ( .A(n_539), .B(n_582), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AOI211x1_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_563), .B(n_576), .C(n_601), .Y(n_549) );
INVx1_ASAP7_75t_L g667 ( .A(n_550), .Y(n_667) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_562), .Y(n_550) );
INVx5_ASAP7_75t_SL g587 ( .A(n_552), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_552), .B(n_657), .Y(n_656) );
AOI311xp33_ASAP7_75t_L g675 ( .A1(n_552), .A2(n_676), .A3(n_678), .B(n_679), .C(n_685), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_552), .A2(n_623), .B(n_711), .C(n_714), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_556), .Y(n_553) );
INVxp67_ASAP7_75t_L g630 ( .A(n_562), .Y(n_630) );
NAND4xp25_ASAP7_75t_SL g563 ( .A(n_564), .B(n_567), .C(n_573), .D(n_575), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_564), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g621 ( .A(n_565), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_568), .B(n_574), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_568), .B(n_581), .Y(n_701) );
BUFx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_569), .B(n_582), .Y(n_719) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g594 ( .A(n_570), .Y(n_594) );
INVxp67_ASAP7_75t_L g629 ( .A(n_571), .Y(n_629) );
AND2x4_ASAP7_75t_L g581 ( .A(n_572), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g655 ( .A(n_572), .B(n_594), .Y(n_655) );
INVx1_ASAP7_75t_L g682 ( .A(n_572), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_572), .B(n_669), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_573), .B(n_643), .Y(n_663) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_574), .B(n_596), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_574), .B(n_643), .Y(n_742) );
INVx1_ASAP7_75t_L g753 ( .A(n_575), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B(n_583), .C(n_591), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g595 ( .A(n_579), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g633 ( .A(n_579), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g615 ( .A(n_580), .Y(n_615) );
AND2x2_ASAP7_75t_L g592 ( .A(n_581), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_581), .B(n_643), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_581), .B(n_662), .Y(n_686) );
OR2x2_ASAP7_75t_L g602 ( .A(n_582), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g634 ( .A(n_582), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_582), .B(n_594), .Y(n_649) );
AND2x2_ASAP7_75t_L g706 ( .A(n_582), .B(n_662), .Y(n_706) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_582), .Y(n_713) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_584), .A2(n_596), .B1(n_718), .B2(n_720), .C(n_723), .Y(n_717) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g607 ( .A(n_587), .B(n_590), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_587), .B(n_657), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_587), .B(n_614), .Y(n_722) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g707 ( .A(n_589), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g721 ( .A(n_589), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_590), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_590), .B(n_611), .Y(n_618) );
AND2x2_ASAP7_75t_L g688 ( .A(n_590), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_590), .B(n_637), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_590), .B(n_738), .Y(n_737) );
OAI21xp5_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_595), .B(n_597), .Y(n_591) );
INVx2_ASAP7_75t_L g624 ( .A(n_592), .Y(n_624) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g644 ( .A(n_594), .Y(n_644) );
OR2x2_ASAP7_75t_L g648 ( .A(n_596), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g751 ( .A(n_596), .B(n_719), .Y(n_751) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_604), .B(n_606), .Y(n_601) );
INVx1_ASAP7_75t_L g755 ( .A(n_602), .Y(n_755) );
INVx2_ASAP7_75t_SL g669 ( .A(n_603), .Y(n_669) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g750 ( .A1(n_606), .A2(n_687), .B(n_751), .C(n_752), .Y(n_750) );
OAI322xp33_ASAP7_75t_SL g619 ( .A1(n_607), .A2(n_620), .A3(n_623), .B1(n_624), .B2(n_625), .C1(n_627), .C2(n_630), .Y(n_619) );
INVx2_ASAP7_75t_L g639 ( .A(n_607), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_615), .B1(n_616), .B2(n_618), .C(n_619), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI22xp33_ASAP7_75t_SL g685 ( .A1(n_610), .A2(n_686), .B1(n_687), .B2(n_690), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_611), .B(n_614), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_611), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g684 ( .A(n_613), .B(n_646), .Y(n_684) );
INVx1_ASAP7_75t_L g674 ( .A(n_614), .Y(n_674) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_618), .A2(n_728), .B(n_730), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_620), .A2(n_653), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2xp67_ASAP7_75t_SL g681 ( .A(n_622), .B(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_622), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g738 ( .A(n_623), .Y(n_738) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_659), .C(n_675), .D(n_691), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_640), .C(n_652), .Y(n_632) );
INVx1_ASAP7_75t_L g724 ( .A(n_633), .Y(n_724) );
AND2x2_ASAP7_75t_L g672 ( .A(n_634), .B(n_655), .Y(n_672) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_639), .B(n_674), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_645), .B1(n_648), .B2(n_650), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_642), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g690 ( .A(n_643), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_643), .A2(n_682), .B(n_705), .C(n_707), .Y(n_704) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g689 ( .A(n_646), .Y(n_689) );
INVx1_ASAP7_75t_L g749 ( .A(n_647), .Y(n_749) );
NAND2xp33_ASAP7_75t_SL g739 ( .A(n_648), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g678 ( .A(n_657), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_664), .C(n_666), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_671), .B2(n_673), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_669), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_674), .B(n_695), .Y(n_757) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI21xp33_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_683), .B(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_697), .B1(n_700), .B2(n_702), .C(n_704), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_707), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_717), .C(n_727), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx16_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_736), .C(n_745), .Y(n_733) );
INVx1_ASAP7_75t_L g754 ( .A(n_734), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B1(n_741), .B2(n_743), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI22x1_ASAP7_75t_SL g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_758) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
NAND2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
endmodule