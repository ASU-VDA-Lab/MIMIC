module fake_jpeg_28065_n_304 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_300;
wire n_294;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_25),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_29),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_13),
.B1(n_26),
.B2(n_24),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_47),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_20),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_13),
.B1(n_26),
.B2(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_27),
.C(n_33),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_70),
.C(n_38),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_48),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_35),
.B1(n_28),
.B2(n_13),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_71),
.Y(n_93)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_26),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_40),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_73),
.B(n_79),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_28),
.B1(n_25),
.B2(n_35),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_89),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_63),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_29),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_90),
.B(n_56),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_92),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_33),
.B1(n_35),
.B2(n_28),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_88),
.B1(n_34),
.B2(n_66),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_45),
.B(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_69),
.B1(n_60),
.B2(n_58),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_122),
.B1(n_34),
.B2(n_25),
.Y(n_149)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_104),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_57),
.C(n_60),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_121),
.C(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_107),
.B(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_115),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_41),
.B(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_109),
.B(n_110),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_41),
.B(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_118),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_19),
.B(n_23),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_93),
.B(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_30),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_83),
.B1(n_78),
.B2(n_85),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_30),
.C(n_29),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_16),
.B1(n_25),
.B2(n_34),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_88),
.B1(n_73),
.B2(n_94),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_126),
.B1(n_132),
.B2(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_124),
.B(n_129),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_87),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_134),
.C(n_139),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_78),
.B(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_42),
.B1(n_85),
.B2(n_68),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_21),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_29),
.C(n_30),
.Y(n_134)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_141),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_149),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_21),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_29),
.C(n_30),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_67),
.C(n_18),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_148),
.B(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_65),
.B1(n_50),
.B2(n_16),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_0),
.B(n_1),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_117),
.B(n_101),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_140),
.B1(n_146),
.B2(n_142),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_102),
.B1(n_121),
.B2(n_104),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_169),
.B1(n_175),
.B2(n_183),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_172),
.B(n_174),
.Y(n_197)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_98),
.B1(n_117),
.B2(n_16),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_164),
.A2(n_166),
.B1(n_185),
.B2(n_154),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_84),
.B1(n_34),
.B2(n_14),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_139),
.C(n_31),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_150),
.B1(n_152),
.B2(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_181),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_R g171 ( 
.A1(n_124),
.A2(n_18),
.B(n_14),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_22),
.B(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_84),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_130),
.A2(n_134),
.B1(n_145),
.B2(n_131),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_21),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_131),
.A2(n_84),
.B1(n_19),
.B2(n_23),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_18),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_84),
.B1(n_14),
.B2(n_23),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_137),
.A2(n_19),
.B1(n_22),
.B2(n_48),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_135),
.B1(n_22),
.B2(n_18),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_205),
.B1(n_208),
.B2(n_187),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_196),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_125),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_195),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_157),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_183),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_133),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_204),
.C(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_206),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_159),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_161),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_31),
.C(n_12),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_211),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_31),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_31),
.C(n_12),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_11),
.C(n_10),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_218),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_161),
.B1(n_180),
.B2(n_155),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_209),
.B1(n_190),
.B2(n_163),
.Y(n_246)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_233),
.B1(n_181),
.B2(n_177),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_191),
.B1(n_177),
.B2(n_158),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_179),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_189),
.C(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_246),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_162),
.B(n_172),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_178),
.B(n_169),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_227),
.B(n_219),
.C(n_230),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_193),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_226),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_233),
.B1(n_221),
.B2(n_225),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_253),
.B(n_260),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_220),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_258),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_216),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_238),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_223),
.C(n_195),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_242),
.C(n_168),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_215),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_263),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_243),
.B1(n_248),
.B2(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_231),
.C(n_204),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_271),
.Y(n_278)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_219),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_252),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_237),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_228),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_249),
.C(n_238),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_275),
.A2(n_262),
.B1(n_173),
.B2(n_185),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_267),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_9),
.B(n_11),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_4),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_268),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_284),
.B(n_4),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_9),
.B(n_2),
.C(n_3),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_268),
.C(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_288),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_0),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_0),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_4),
.B(n_5),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_6),
.B(n_7),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_4),
.B(n_5),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_6),
.B(n_7),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_289),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_301),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_302),
.A2(n_294),
.B(n_287),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_6),
.B1(n_299),
.B2(n_266),
.Y(n_304)
);


endmodule