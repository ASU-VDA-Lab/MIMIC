module fake_jpeg_9249_n_81 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_7),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_67)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_43),
.B1(n_40),
.B2(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_57),
.B1(n_5),
.B2(n_6),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_0),
.B1(n_32),
.B2(n_4),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_1),
.Y(n_65)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_8),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_64),
.B1(n_71),
.B2(n_12),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_70),
.C(n_68),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_67),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_66),
.B(n_11),
.Y(n_76)
);

OAI21x1_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_10),
.B(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_14),
.B(n_16),
.Y(n_79)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_17),
.B(n_19),
.C(n_21),
.D(n_22),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_23),
.Y(n_81)
);


endmodule