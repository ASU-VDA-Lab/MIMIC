module real_jpeg_13281_n_17 (n_5, n_4, n_8, n_0, n_12, n_309, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_309;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx2_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_43),
.B1(n_47),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_52),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_4),
.A2(n_43),
.B1(n_47),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_4),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_139),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_139),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_139),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_5),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_43),
.B1(n_47),
.B2(n_134),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_134),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_134),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_7),
.A2(n_35),
.B1(n_43),
.B2(n_47),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_10),
.A2(n_38),
.B1(n_43),
.B2(n_47),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_43),
.B1(n_47),
.B2(n_65),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_65),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_12),
.B(n_27),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_13),
.A2(n_43),
.B1(n_47),
.B2(n_59),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_14),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_93),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_14),
.A2(n_43),
.B1(n_47),
.B2(n_93),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_93),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_15),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_43),
.C(n_46),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_15),
.B(n_30),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_15),
.A2(n_137),
.B(n_140),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_15),
.A2(n_28),
.B(n_29),
.C(n_168),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_15),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_15),
.B(n_57),
.Y(n_214)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_107),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_20),
.B(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.C(n_75),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_21),
.B(n_67),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_54),
.B1(n_55),
.B2(n_66),
.Y(n_21)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_39),
.B1(n_40),
.B2(n_53),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_23),
.B(n_40),
.C(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_24),
.B(n_175),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_26),
.A2(n_31),
.B(n_122),
.Y(n_168)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g226 ( 
.A1(n_29),
.A2(n_58),
.A3(n_62),
.B1(n_214),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_30),
.B(n_175),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_49)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_32),
.B(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_37),
.A2(n_69),
.B1(n_71),
.B2(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_39),
.A2(n_40),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_48),
.B(n_50),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_41),
.A2(n_48),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_41),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_41),
.A2(n_48),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_41),
.A2(n_48),
.B1(n_220),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_41),
.A2(n_48),
.B1(n_86),
.B2(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_51),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_42),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_42),
.B(n_122),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_42),
.A2(n_135),
.B(n_219),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_47),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_48),
.B(n_124),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_55),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_61),
.B(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_58),
.A2(n_60),
.B(n_122),
.C(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_60),
.A2(n_61),
.B1(n_241),
.B2(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_60),
.A2(n_261),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_61),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_61),
.B(n_92),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_61),
.A2(n_89),
.B(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_67),
.A2(n_68),
.B(n_72),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_69),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_69),
.A2(n_71),
.B1(n_188),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_69),
.A2(n_174),
.B(n_217),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_263),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_71),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_71),
.A2(n_189),
.B(n_263),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_121),
.B(n_123),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_73),
.A2(n_123),
.B(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_75),
.B(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B(n_88),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_76),
.A2(n_77),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_78),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_78),
.A2(n_79),
.B1(n_88),
.B2(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_81),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_80),
.A2(n_81),
.B1(n_231),
.B2(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_81),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_81),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_83),
.A2(n_137),
.B1(n_154),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_88),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_303),
.B(n_307),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_290),
.B(n_302),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_273),
.B(n_289),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_233),
.A3(n_266),
.B1(n_271),
.B2(n_272),
.C(n_309),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_205),
.B(n_232),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_182),
.B(n_204),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_163),
.B(n_181),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_142),
.B(n_162),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_127),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_125),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_120),
.B1(n_125),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_154),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_132),
.C(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_137),
.A2(n_154),
.B1(n_170),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_137),
.A2(n_154),
.B1(n_196),
.B2(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_150),
.B(n_161),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_148),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_156),
.B(n_160),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_155),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_165),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_176),
.C(n_180),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_197),
.B2(n_198),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_200),
.C(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_191),
.C(n_195),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_207),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_222),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_208),
.B(n_223),
.C(n_224),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_221),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_216),
.C(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_250),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_244),
.C(n_249),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_236),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_247),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_265),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_258),
.C(n_265),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_256),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_262),
.C(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_288),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_288),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_284),
.C(n_287),
.Y(n_301)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.C(n_301),
.Y(n_306)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_306),
.Y(n_307)
);


endmodule