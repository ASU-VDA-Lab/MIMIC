module real_jpeg_27451_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_50;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx11_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_3),
.A2(n_12),
.B1(n_13),
.B2(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_5),
.B(n_13),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_4),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_4),
.A2(n_15),
.B1(n_41),
.B2(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_12),
.B1(n_13),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_23),
.B1(n_41),
.B2(n_45),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_34),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_28),
.B(n_33),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_24),
.Y(n_8)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_11),
.B(n_16),
.Y(n_9)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_10),
.A2(n_11),
.B1(n_18),
.B2(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_19),
.Y(n_18)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_21),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_23),
.A2(n_31),
.B(n_40),
.C(n_41),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_32),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_50),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_41),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_53),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_52),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_47),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);


endmodule