module fake_aes_2739_n_706 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_706);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_706;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_8), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_2), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_70), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_49), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_24), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_31), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_9), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_51), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_63), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_46), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_76), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_8), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_21), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_72), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_69), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_0), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_56), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_34), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_35), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_37), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_14), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_29), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_33), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_64), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_30), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_44), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_3), .Y(n_114) );
NOR2xp33_ASAP7_75t_R g115 ( .A(n_10), .B(n_78), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_58), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_61), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_42), .Y(n_122) );
CKINVDCx14_ASAP7_75t_R g123 ( .A(n_68), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_17), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_25), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_45), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_84), .B(n_27), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
XOR2xp5_ASAP7_75t_L g132 ( .A(n_86), .B(n_1), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_93), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_103), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_96), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_97), .Y(n_142) );
NOR2xp33_ASAP7_75t_SL g143 ( .A(n_84), .B(n_28), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_104), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_80), .B(n_2), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_101), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_103), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_94), .B(n_110), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_104), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_111), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_122), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_91), .B(n_3), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_105), .Y(n_163) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_126), .A2(n_32), .B(n_74), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_79), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_92), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_99), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_106), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_112), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_91), .B(n_116), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_170), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_154), .B(n_116), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
OR2x2_ASAP7_75t_SL g176 ( .A(n_132), .B(n_117), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_127), .B(n_109), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_167), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_165), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
OAI221xp5_ASAP7_75t_L g183 ( .A1(n_167), .A2(n_119), .B1(n_113), .B2(n_114), .C(n_83), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_127), .B(n_108), .Y(n_185) );
INVx4_ASAP7_75t_SL g186 ( .A(n_128), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_165), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_146), .B(n_123), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_131), .B(n_108), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_128), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_163), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_168), .B(n_123), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_139), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
OR2x6_ASAP7_75t_L g199 ( .A(n_164), .B(n_125), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
OR2x6_ASAP7_75t_L g201 ( .A(n_164), .B(n_125), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_131), .A2(n_109), .B1(n_107), .B2(n_121), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_133), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_134), .B(n_107), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_156), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_134), .B(n_100), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_136), .B(n_85), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_136), .B(n_121), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_153), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_137), .B(n_4), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_137), .B(n_105), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_128), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_140), .B(n_4), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_169), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_133), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_140), .B(n_115), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_157), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_169), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_169), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_157), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_133), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_169), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_128), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_142), .B(n_5), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_217), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_220), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_220), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_194), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_194), .B(n_149), .Y(n_238) );
BUFx4f_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_189), .B(n_149), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_189), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_171), .B(n_150), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_185), .B(n_150), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_220), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_217), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_178), .B(n_143), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_215), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_193), .B(n_160), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_193), .B(n_160), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_211), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_199), .B(n_142), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_181), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_196), .B(n_158), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_197), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_187), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_172), .B(n_158), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_179), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_222), .B(n_143), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_177), .B(n_152), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_212), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_210), .A2(n_152), .B1(n_157), .B2(n_129), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_224), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_198), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_174), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_175), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_175), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_200), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_187), .Y(n_275) );
CKINVDCx11_ASAP7_75t_R g276 ( .A(n_197), .Y(n_276) );
BUFx12f_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_188), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_227), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_209), .B(n_162), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_190), .B(n_162), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_202), .B(n_132), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_192), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_206), .B(n_162), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_204), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_221), .B(n_159), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_199), .B(n_159), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_183), .A2(n_159), .B1(n_151), .B2(n_133), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_228), .B(n_151), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_199), .Y(n_293) );
CKINVDCx11_ASAP7_75t_R g294 ( .A(n_201), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_188), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_231), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_205), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_239), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_245), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_245), .Y(n_300) );
CKINVDCx6p67_ASAP7_75t_R g301 ( .A(n_276), .Y(n_301) );
O2A1O1Ixp5_ASAP7_75t_SL g302 ( .A1(n_247), .A2(n_141), .B(n_151), .C(n_208), .Y(n_302) );
OAI22x1_ASAP7_75t_L g303 ( .A1(n_259), .A2(n_176), .B1(n_201), .B2(n_151), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_236), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_285), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_248), .A2(n_201), .B(n_173), .C(n_141), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_242), .B(n_201), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_265), .A2(n_141), .B(n_195), .C(n_180), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_255), .B(n_176), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_250), .A2(n_141), .B1(n_224), .B2(n_226), .C(n_225), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_239), .A2(n_218), .B1(n_205), .B2(n_208), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_277), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_255), .B(n_6), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_245), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_262), .B(n_7), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_252), .B(n_214), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_254), .B(n_214), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_262), .A2(n_214), .B1(n_229), .B2(n_226), .C(n_225), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_238), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_234), .B(n_225), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_241), .B(n_9), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_239), .A2(n_296), .B(n_261), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_270), .Y(n_327) );
AOI221x1_ASAP7_75t_L g328 ( .A1(n_289), .A2(n_218), .B1(n_130), .B2(n_135), .C(n_138), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_240), .A2(n_184), .B(n_195), .C(n_207), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_244), .A2(n_229), .B(n_226), .Y(n_330) );
INVx4_ASAP7_75t_L g331 ( .A(n_234), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_241), .Y(n_332) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_266), .B(n_144), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_282), .A2(n_184), .B(n_207), .C(n_180), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_237), .B(n_10), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_233), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_264), .B(n_229), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_256), .A2(n_144), .B1(n_130), .B2(n_135), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_258), .A2(n_144), .B(n_138), .C(n_135), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_235), .A2(n_230), .B(n_216), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_235), .A2(n_230), .B(n_216), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_270), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_259), .Y(n_345) );
INVx4_ASAP7_75t_L g346 ( .A(n_234), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_246), .A2(n_130), .B(n_138), .C(n_128), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_234), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
CKINVDCx6p67_ASAP7_75t_R g351 ( .A(n_301), .Y(n_351) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_323), .A2(n_276), .B1(n_243), .B2(n_294), .C1(n_277), .C2(n_289), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_326), .A2(n_247), .B(n_263), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_302), .A2(n_263), .B(n_293), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_331), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_312), .B(n_284), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_350), .B(n_256), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_347), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_329), .A2(n_289), .B(n_267), .Y(n_360) );
NOR2xp67_ASAP7_75t_L g361 ( .A(n_331), .B(n_234), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_307), .A2(n_286), .B(n_283), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_336), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_307), .A2(n_288), .B(n_274), .Y(n_365) );
AOI22x1_ASAP7_75t_L g366 ( .A1(n_319), .A2(n_147), .B1(n_148), .B2(n_145), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_299), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_329), .A2(n_273), .B(n_269), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_334), .A2(n_278), .B(n_279), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_321), .Y(n_372) );
OAI21x1_ASAP7_75t_SL g373 ( .A1(n_308), .A2(n_256), .B(n_294), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_299), .Y(n_374) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_346), .B(n_256), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_299), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_334), .A2(n_339), .B(n_328), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_299), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_310), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_341), .B(n_290), .Y(n_381) );
OAI21x1_ASAP7_75t_SL g382 ( .A1(n_311), .A2(n_281), .B(n_297), .Y(n_382) );
AOI21x1_ASAP7_75t_L g383 ( .A1(n_338), .A2(n_249), .B(n_251), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_356), .A2(n_312), .B1(n_303), .B2(n_316), .C(n_332), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_371), .A2(n_339), .B(n_311), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_363), .A2(n_316), .B(n_325), .C(n_335), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_358), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_363), .A2(n_335), .B1(n_315), .B2(n_318), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_381), .A2(n_343), .B1(n_284), .B2(n_309), .C(n_304), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_352), .A2(n_345), .B1(n_315), .B2(n_298), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_298), .B1(n_322), .B2(n_313), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_368), .A2(n_348), .B(n_349), .C(n_330), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_381), .B(n_348), .C(n_349), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_357), .A2(n_232), .B1(n_272), .B2(n_271), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_357), .B(n_300), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_353), .A2(n_342), .B(n_340), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_306), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_373), .A2(n_333), .B1(n_300), .B2(n_306), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_364), .A2(n_337), .B1(n_314), .B2(n_272), .C(n_232), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_371), .A2(n_344), .B(n_327), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_369), .A2(n_317), .B1(n_271), .B2(n_324), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_351), .A2(n_270), .B1(n_324), .B2(n_268), .Y(n_404) );
OA21x2_ASAP7_75t_L g405 ( .A1(n_371), .A2(n_297), .B(n_295), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_369), .B(n_268), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_360), .A2(n_295), .B(n_280), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_372), .B(n_268), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_359), .B(n_268), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g411 ( .A1(n_360), .A2(n_145), .B(n_147), .C(n_148), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_380), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_390), .A2(n_373), .B1(n_382), .B2(n_355), .Y(n_413) );
OAI31xp33_ASAP7_75t_L g414 ( .A1(n_388), .A2(n_386), .A3(n_407), .B(n_391), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_399), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_397), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_400), .A2(n_375), .B1(n_355), .B2(n_377), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_397), .B(n_380), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_412), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_412), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_405), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_395), .B(n_374), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_406), .B(n_377), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_405), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_406), .B(n_377), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_393), .B(n_365), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_395), .B(n_377), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_389), .B(n_365), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_398), .B(n_365), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_384), .B(n_370), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_402), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_402), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_392), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_362), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_385), .B(n_362), .Y(n_446) );
BUFx2_ASAP7_75t_SL g447 ( .A(n_408), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_423), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_420), .B(n_385), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_422), .B(n_351), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_423), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_420), .B(n_370), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_420), .B(n_370), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_431), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_440), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_414), .A2(n_401), .B1(n_382), .B2(n_375), .Y(n_458) );
AOI21xp5_ASAP7_75t_SL g459 ( .A1(n_418), .A2(n_411), .B(n_404), .Y(n_459) );
NOR2x1_ASAP7_75t_SL g460 ( .A(n_418), .B(n_374), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_424), .B(n_362), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_424), .B(n_394), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_421), .B(n_378), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_434), .B(n_396), .C(n_361), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_419), .B(n_379), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_436), .B(n_374), .Y(n_468) );
AO31x2_ASAP7_75t_L g469 ( .A1(n_437), .A2(n_379), .A3(n_367), .B(n_378), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_440), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_414), .A2(n_376), .B1(n_367), .B2(n_379), .C(n_14), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_415), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_434), .A2(n_145), .B1(n_147), .B2(n_148), .C(n_376), .Y(n_474) );
OAI321xp33_ASAP7_75t_L g475 ( .A1(n_413), .A2(n_383), .A3(n_148), .B1(n_147), .B2(n_145), .C(n_367), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_444), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_436), .B(n_354), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_435), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_415), .B(n_378), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_438), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_415), .B(n_354), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_417), .B(n_354), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_429), .A2(n_361), .B1(n_366), .B2(n_145), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_429), .A2(n_366), .B1(n_145), .B2(n_148), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_432), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_419), .B(n_11), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_417), .B(n_12), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_417), .B(n_13), .Y(n_492) );
OAI211xp5_ASAP7_75t_SL g493 ( .A1(n_430), .A2(n_249), .B(n_251), .C(n_280), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_438), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_430), .A2(n_383), .B1(n_147), .B2(n_148), .C(n_260), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_476), .B(n_446), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_456), .B(n_429), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_488), .B(n_442), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_459), .B(n_439), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_448), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_470), .B(n_442), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_455), .B(n_426), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_463), .B(n_426), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_489), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_476), .B(n_446), .Y(n_507) );
INVxp67_ASAP7_75t_L g508 ( .A(n_489), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g509 ( .A(n_491), .B(n_425), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_468), .B(n_439), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_491), .B(n_425), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_463), .B(n_428), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_468), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_459), .B(n_439), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_462), .A2(n_429), .B1(n_433), .B2(n_428), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_451), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_492), .B(n_433), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_492), .B(n_437), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_468), .B(n_425), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_468), .B(n_425), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_473), .B(n_427), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_473), .B(n_427), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_466), .B(n_445), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_472), .B(n_443), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_496), .B(n_441), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_484), .B(n_439), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_484), .B(n_443), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_496), .B(n_445), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_457), .B(n_15), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_457), .B(n_15), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_471), .B(n_16), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_464), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_471), .B(n_447), .Y(n_534) );
OAI31xp33_ASAP7_75t_SL g535 ( .A1(n_493), .A2(n_447), .A3(n_19), .B(n_20), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_448), .B(n_147), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_448), .B(n_18), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_490), .B(n_22), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_464), .B(n_23), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_449), .B(n_26), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_458), .A2(n_182), .B1(n_191), .B2(n_216), .C(n_257), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_449), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_38), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_453), .B(n_39), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_453), .B(n_40), .Y(n_546) );
NOR3xp33_ASAP7_75t_SL g547 ( .A(n_475), .B(n_43), .C(n_47), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_477), .B(n_48), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_452), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_477), .B(n_50), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_452), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_452), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_454), .B(n_53), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_467), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_528), .B(n_479), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_497), .B(n_450), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_497), .B(n_477), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_516), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_507), .B(n_450), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_507), .B(n_454), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_499), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_506), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_523), .B(n_480), .Y(n_563) );
NAND4xp25_ASAP7_75t_L g564 ( .A(n_524), .B(n_465), .C(n_474), .D(n_495), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_500), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_549), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_526), .B(n_480), .Y(n_567) );
AOI211xp5_ASAP7_75t_SL g568 ( .A1(n_524), .A2(n_475), .B(n_481), .C(n_479), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_533), .B(n_494), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_506), .B(n_494), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_526), .B(n_494), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_504), .B(n_481), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_503), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_512), .B(n_481), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_549), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_510), .B(n_479), .Y(n_578) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_552), .Y(n_579) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_513), .B(n_467), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_531), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_529), .B(n_467), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_501), .B(n_478), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g584 ( .A1(n_514), .A2(n_485), .B(n_478), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_510), .B(n_485), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_510), .B(n_485), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_525), .B(n_478), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_498), .B(n_483), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_517), .B(n_483), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_515), .B(n_482), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_527), .B(n_482), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_552), .B(n_469), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_530), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_542), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_551), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_532), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_469), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_554), .B(n_469), .Y(n_599) );
NOR2xp33_ASAP7_75t_SL g600 ( .A(n_548), .B(n_460), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_508), .B(n_469), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_518), .B(n_469), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_519), .B(n_469), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_520), .B(n_460), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_538), .B(n_54), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_502), .B(n_486), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_502), .B(n_487), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_557), .B(n_534), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_581), .A2(n_548), .B1(n_550), .B2(n_543), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_565), .Y(n_610) );
AOI322xp5_ASAP7_75t_L g611 ( .A1(n_558), .A2(n_539), .A3(n_547), .B1(n_548), .B2(n_541), .C1(n_545), .C2(n_546), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_580), .B(n_540), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_557), .B(n_509), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_561), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_597), .A2(n_539), .B1(n_511), .B2(n_509), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_573), .Y(n_616) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_574), .B(n_583), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_593), .B(n_553), .Y(n_618) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_604), .A2(n_511), .B1(n_521), .B2(n_522), .C1(n_537), .C2(n_536), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_600), .A2(n_535), .B(n_541), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_568), .A2(n_547), .B1(n_230), .B2(n_62), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_602), .B(n_55), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_602), .B(n_59), .Y(n_625) );
AOI32xp33_ASAP7_75t_L g626 ( .A1(n_562), .A2(n_65), .A3(n_66), .B1(n_71), .B2(n_73), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_559), .B(n_77), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_559), .B(n_182), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_595), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_562), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_582), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_563), .B(n_182), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_572), .Y(n_634) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_601), .A2(n_182), .B(n_191), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_556), .B(n_182), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_555), .Y(n_639) );
AOI21xp5_ASAP7_75t_SL g640 ( .A1(n_566), .A2(n_191), .B(n_216), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_555), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_603), .B(n_191), .Y(n_642) );
AOI32xp33_ASAP7_75t_L g643 ( .A1(n_603), .A2(n_253), .A3(n_260), .B1(n_257), .B2(n_275), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_570), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_632), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_634), .B(n_563), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_622), .A2(n_564), .B(n_583), .C(n_584), .Y(n_648) );
NOR3x1_ASAP7_75t_L g649 ( .A(n_631), .B(n_590), .C(n_579), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_611), .A2(n_580), .B(n_604), .C(n_605), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_628), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_640), .A2(n_592), .B(n_601), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_608), .B(n_567), .Y(n_653) );
BUFx3_ASAP7_75t_L g654 ( .A(n_633), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_636), .B(n_567), .Y(n_655) );
AO21x1_ASAP7_75t_L g656 ( .A1(n_621), .A2(n_587), .B(n_577), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
OAI222xp33_ASAP7_75t_L g658 ( .A1(n_609), .A2(n_560), .B1(n_589), .B2(n_588), .C1(n_578), .C2(n_586), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_642), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_618), .A2(n_578), .B1(n_586), .B2(n_585), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_627), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_613), .B(n_585), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_642), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_628), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_630), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_610), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_644), .A2(n_591), .B(n_592), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_615), .A2(n_571), .B1(n_599), .B2(n_598), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_648), .A2(n_625), .B(n_624), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_659), .B(n_620), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_650), .A2(n_626), .B(n_643), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_646), .Y(n_673) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_650), .A2(n_614), .B(n_616), .C(n_624), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_657), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_654), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_659), .B(n_645), .Y(n_677) );
OAI321xp33_ASAP7_75t_L g678 ( .A1(n_664), .A2(n_612), .A3(n_625), .B1(n_638), .B2(n_639), .C(n_641), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_669), .A2(n_617), .B1(n_637), .B2(n_571), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_654), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_668), .A2(n_612), .B(n_599), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_664), .B(n_598), .Y(n_682) );
NOR4xp25_ASAP7_75t_L g683 ( .A(n_658), .B(n_635), .C(n_619), .D(n_606), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_652), .B1(n_661), .B2(n_660), .C(n_665), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_676), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_672), .A2(n_649), .B(n_656), .C(n_647), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_674), .B(n_665), .C(n_651), .Y(n_687) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_676), .A2(n_651), .B(n_635), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_670), .A2(n_667), .B(n_666), .C(n_663), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_681), .A2(n_655), .B1(n_653), .B2(n_569), .C(n_662), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_679), .A2(n_577), .B1(n_587), .B2(n_607), .Y(n_691) );
NOR3x1_ASAP7_75t_L g692 ( .A(n_684), .B(n_671), .C(n_677), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_685), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_687), .B(n_682), .Y(n_694) );
NAND4xp75_ASAP7_75t_L g695 ( .A(n_691), .B(n_680), .C(n_673), .D(n_675), .Y(n_695) );
AND4x1_ASAP7_75t_L g696 ( .A(n_686), .B(n_678), .C(n_186), .D(n_230), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g697 ( .A(n_696), .B(n_688), .C(n_689), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_693), .B(n_690), .Y(n_698) );
OAI211xp5_ASAP7_75t_SL g699 ( .A1(n_694), .A2(n_253), .B(n_275), .C(n_230), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_698), .A2(n_695), .B1(n_692), .B2(n_216), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_697), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_701), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_700), .B1(n_699), .B2(n_191), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_703), .Y(n_704) );
NOR3x1_ASAP7_75t_L g705 ( .A(n_704), .B(n_186), .C(n_268), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_186), .B(n_701), .Y(n_706) );
endmodule