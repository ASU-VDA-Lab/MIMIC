module fake_jpeg_14488_n_375 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_23),
.A2(n_40),
.B(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_58),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_9),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_34),
.Y(n_62)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_21),
.B(n_10),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_86),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_16),
.B(n_22),
.C(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

NOR2xp67_ASAP7_75t_L g82 ( 
.A(n_17),
.B(n_7),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_32),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_94),
.B(n_101),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_25),
.B1(n_32),
.B2(n_39),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_95),
.A2(n_120),
.B(n_115),
.C(n_140),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_113),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_103),
.B(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_117),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_69),
.B(n_0),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_61),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_29),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_25),
.B1(n_42),
.B2(n_17),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_39),
.B1(n_33),
.B2(n_22),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_44),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_129),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_45),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_51),
.B(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_133),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_28),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_54),
.A2(n_33),
.B1(n_20),
.B2(n_38),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_127),
.B1(n_123),
.B2(n_131),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx2_ASAP7_75t_SL g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_164),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_20),
.B1(n_38),
.B2(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_150),
.B(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_73),
.B1(n_68),
.B2(n_75),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_169),
.B(n_162),
.Y(n_225)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_155),
.B1(n_161),
.B2(n_167),
.Y(n_200)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_88),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_134),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_162),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_165),
.B1(n_175),
.B2(n_180),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_102),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_11),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_168),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_90),
.A2(n_14),
.B1(n_15),
.B2(n_92),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_125),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_168),
.B1(n_154),
.B2(n_156),
.Y(n_214)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_172),
.Y(n_208)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_174),
.Y(n_217)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_177),
.B(n_181),
.Y(n_223)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_95),
.B1(n_109),
.B2(n_122),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_184),
.B(n_186),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_108),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_120),
.A2(n_139),
.B1(n_87),
.B2(n_128),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_111),
.B1(n_138),
.B2(n_115),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_135),
.B1(n_105),
.B2(n_97),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_199),
.B1(n_201),
.B2(n_219),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_97),
.B1(n_87),
.B2(n_128),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_204),
.B1(n_224),
.B2(n_225),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_130),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_206),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_105),
.B1(n_135),
.B2(n_111),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_138),
.B1(n_130),
.B2(n_107),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_175),
.A2(n_146),
.B1(n_155),
.B2(n_144),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_143),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_164),
.B1(n_173),
.B2(n_181),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_196),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_143),
.A2(n_175),
.B1(n_182),
.B2(n_145),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_142),
.B(n_159),
.C(n_175),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_194),
.C(n_204),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_160),
.A2(n_165),
.B1(n_178),
.B2(n_157),
.Y(n_224)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_233),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_149),
.B1(n_202),
.B2(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_248),
.B1(n_252),
.B2(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_203),
.Y(n_234)
);

BUFx24_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_242),
.C(n_251),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_192),
.B(n_223),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_234),
.B(n_232),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_196),
.B(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_209),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_250),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_201),
.B1(n_224),
.B2(n_214),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_215),
.B(n_198),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_251),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_218),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_200),
.B(n_197),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_218),
.B(n_198),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_254),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_209),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_228),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_190),
.B1(n_207),
.B2(n_222),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_259),
.A2(n_237),
.B1(n_235),
.B2(n_254),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_260),
.A2(n_242),
.B1(n_238),
.B2(n_243),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_273),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_230),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_271),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_255),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_239),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_241),
.C(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_240),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_227),
.B(n_252),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_299),
.C(n_276),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_257),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_293),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_253),
.B(n_238),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_287),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_297),
.B1(n_298),
.B2(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_235),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_235),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_260),
.A2(n_261),
.B1(n_278),
.B2(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_258),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_252),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_227),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_301),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_261),
.A2(n_226),
.B1(n_262),
.B2(n_263),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_273),
.C(n_256),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_302),
.B(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_310),
.A2(n_267),
.B(n_286),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_268),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_268),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_319),
.C(n_296),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_280),
.C(n_269),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_289),
.B1(n_284),
.B2(n_264),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_324),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_308),
.A2(n_287),
.B1(n_267),
.B2(n_272),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_331),
.Y(n_336)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_306),
.B(n_312),
.Y(n_337)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_265),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_332),
.A2(n_333),
.B1(n_334),
.B2(n_304),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_318),
.B1(n_314),
.B2(n_316),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_309),
.C(n_314),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_311),
.C(n_315),
.Y(n_339)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_339),
.B(n_340),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_306),
.C(n_310),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_324),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_333),
.A2(n_283),
.B1(n_285),
.B2(n_295),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_344),
.B(n_345),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_325),
.C(n_329),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_323),
.C(n_322),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_343),
.Y(n_361)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_336),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_353),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_346),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_328),
.C(n_327),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_347),
.Y(n_362)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_352),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_357),
.B(n_359),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_337),
.B(n_342),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_358),
.A2(n_360),
.B(n_362),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_348),
.A2(n_340),
.B(n_339),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_274),
.C(n_275),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_363),
.A2(n_364),
.B1(n_274),
.B2(n_275),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g364 ( 
.A1(n_358),
.A2(n_344),
.A3(n_338),
.B1(n_321),
.B2(n_283),
.C1(n_350),
.C2(n_341),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_356),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_367),
.B(n_368),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_366),
.A2(n_361),
.B(n_277),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_270),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_371),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_372),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_370),
.C(n_270),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_270),
.Y(n_375)
);


endmodule