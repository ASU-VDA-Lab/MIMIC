module fake_jpeg_23107_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_9),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_19),
.B1(n_15),
.B2(n_13),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_27),
.B(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_11),
.B1(n_19),
.B2(n_20),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_35),
.B1(n_28),
.B2(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_22),
.B(n_17),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_45),
.B(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_47),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_48),
.B1(n_49),
.B2(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_23),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_27),
.C(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_12),
.B1(n_18),
.B2(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_21),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_27),
.B1(n_26),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_23),
.B1(n_10),
.B2(n_15),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_10),
.B1(n_15),
.B2(n_4),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_61),
.C(n_45),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_3),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_40),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_75),
.B1(n_73),
.B2(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_42),
.C(n_50),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_65),
.C(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_54),
.B1(n_72),
.B2(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_65),
.B(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_54),
.B1(n_75),
.B2(n_78),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_92),
.B(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_62),
.B1(n_67),
.B2(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_62),
.B1(n_56),
.B2(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_63),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_83),
.B2(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_91),
.C(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_89),
.A3(n_85),
.B1(n_83),
.B2(n_59),
.C1(n_55),
.C2(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_8),
.B(n_6),
.Y(n_104)
);

NAND4xp25_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_105),
.C(n_8),
.D(n_106),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_7),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_8),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule