module fake_jpeg_18563_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_3),
.Y(n_13)
);

BUFx2_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_24),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_2),
.C(n_4),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_19),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_25),
.B(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_31),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_19),
.B1(n_10),
.B2(n_18),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_42),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_16),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_25),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_34),
.C(n_33),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_30),
.B1(n_33),
.B2(n_18),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_21),
.B(n_22),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_44),
.B1(n_46),
.B2(n_2),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_11),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_13),
.B(n_26),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_10),
.B1(n_15),
.B2(n_17),
.Y(n_44)
);

OAI31xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_9),
.A3(n_16),
.B(n_11),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_10),
.B1(n_15),
.B2(n_17),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_50),
.C(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_51),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_50),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_38),
.C(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_37),
.C(n_51),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI221xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_46),
.B2(n_56),
.C(n_52),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_2),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_6),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_67),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_71)
);


endmodule