module fake_jpeg_26192_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_4),
.B(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_22),
.B1(n_17),
.B2(n_14),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_16),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_22),
.B1(n_14),
.B2(n_18),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_42),
.B1(n_35),
.B2(n_24),
.Y(n_68)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_53),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_31),
.C(n_12),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_37),
.C(n_12),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_51),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_14),
.B1(n_37),
.B2(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_52),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_77),
.B1(n_59),
.B2(n_58),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_55),
.B1(n_61),
.B2(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_91),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_77),
.B1(n_65),
.B2(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_65),
.B(n_74),
.C(n_66),
.D(n_69),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_19),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_71),
.C(n_57),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_99),
.C(n_87),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_30),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_37),
.C(n_46),
.Y(n_99)
);

HAxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_46),
.CON(n_101),
.SN(n_101)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_108),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_89),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_106),
.B1(n_112),
.B2(n_107),
.Y(n_118)
);

FAx1_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_86),
.CI(n_84),
.CON(n_106),
.SN(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_102),
.C(n_93),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_115),
.B(n_117),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_101),
.A3(n_92),
.B1(n_95),
.B2(n_96),
.C1(n_12),
.C2(n_25),
.Y(n_116)
);

AOI31xp67_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_119),
.A3(n_6),
.B(n_72),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_25),
.C(n_13),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_13),
.B(n_15),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_18),
.A3(n_7),
.B1(n_6),
.B2(n_10),
.C1(n_11),
.C2(n_75),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_118),
.B(n_15),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_123),
.B1(n_44),
.B2(n_3),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_2),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_72),
.C(n_29),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_5),
.C(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_128),
.B(n_124),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_127),
.Y(n_131)
);


endmodule