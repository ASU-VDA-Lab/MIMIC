module fake_aes_12691_n_57 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_57);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_57;
wire n_53;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_54;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_48;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_33;
wire n_50;
wire n_52;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_55;
wire n_17;
wire n_56;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_51;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_6), .B1(n_14), .B2(n_9), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_1), .A2(n_10), .B1(n_13), .B2(n_3), .Y(n_18) );
INVx5_ASAP7_75t_L g19 ( .A(n_3), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_4), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_10), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_7), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_7), .B(n_8), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_22), .B(n_0), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_22), .Y(n_28) );
O2A1O1Ixp33_ASAP7_75t_L g29 ( .A1(n_20), .A2(n_0), .B(n_1), .C(n_2), .Y(n_29) );
NAND2x1_ASAP7_75t_L g30 ( .A(n_21), .B(n_2), .Y(n_30) );
OAI21x1_ASAP7_75t_L g31 ( .A1(n_26), .A2(n_25), .B(n_24), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_28), .B(n_23), .Y(n_32) );
OAI21x1_ASAP7_75t_L g33 ( .A1(n_26), .A2(n_18), .B(n_17), .Y(n_33) );
AND2x4_ASAP7_75t_L g34 ( .A(n_31), .B(n_27), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_31), .A2(n_27), .B1(n_30), .B2(n_19), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_34), .B(n_32), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
OA21x2_ASAP7_75t_L g38 ( .A1(n_34), .A2(n_31), .B(n_33), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_36), .B(n_34), .Y(n_39) );
NOR2xp33_ASAP7_75t_L g40 ( .A(n_37), .B(n_34), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_37), .Y(n_41) );
AND4x1_ASAP7_75t_SL g42 ( .A(n_39), .B(n_41), .C(n_33), .D(n_30), .Y(n_42) );
OAI21xp33_ASAP7_75t_SL g43 ( .A1(n_40), .A2(n_35), .B(n_38), .Y(n_43) );
NOR3xp33_ASAP7_75t_L g44 ( .A(n_39), .B(n_29), .C(n_35), .Y(n_44) );
NAND2xp5_ASAP7_75t_SL g45 ( .A(n_39), .B(n_19), .Y(n_45) );
NOR3x1_ASAP7_75t_SL g46 ( .A(n_42), .B(n_4), .C(n_5), .Y(n_46) );
NAND4xp25_ASAP7_75t_SL g47 ( .A(n_44), .B(n_5), .C(n_6), .D(n_8), .Y(n_47) );
AOI22xp5_ASAP7_75t_L g48 ( .A1(n_43), .A2(n_38), .B1(n_19), .B2(n_12), .Y(n_48) );
AOI221xp5_ASAP7_75t_L g49 ( .A1(n_45), .A2(n_19), .B1(n_38), .B2(n_13), .C(n_14), .Y(n_49) );
XOR2xp5_ASAP7_75t_L g50 ( .A(n_47), .B(n_9), .Y(n_50) );
INVx2_ASAP7_75t_L g51 ( .A(n_48), .Y(n_51) );
BUFx3_ASAP7_75t_L g52 ( .A(n_46), .Y(n_52) );
OR2x2_ASAP7_75t_L g53 ( .A(n_49), .B(n_11), .Y(n_53) );
HB1xp67_ASAP7_75t_L g54 ( .A(n_51), .Y(n_54) );
OAI22xp5_ASAP7_75t_L g55 ( .A1(n_50), .A2(n_42), .B1(n_15), .B2(n_16), .Y(n_55) );
AOI22xp5_ASAP7_75t_L g56 ( .A1(n_55), .A2(n_52), .B1(n_51), .B2(n_53), .Y(n_56) );
OAI21x1_ASAP7_75t_L g57 ( .A1(n_56), .A2(n_54), .B(n_53), .Y(n_57) );
endmodule