module real_aes_16765_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g498 ( .A(n_0), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_1), .A2(n_84), .B1(n_580), .B2(n_581), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_1), .A2(n_271), .B1(n_598), .B2(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g503 ( .A(n_2), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_2), .A2(n_160), .B1(n_552), .B2(n_556), .C(n_558), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_3), .A2(n_221), .B1(n_1291), .B2(n_1295), .Y(n_1318) );
INVx1_ASAP7_75t_L g1145 ( .A(n_4), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_4), .A2(n_121), .B1(n_600), .B2(n_666), .Y(n_1159) );
INVx1_ASAP7_75t_L g592 ( .A(n_5), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_6), .A2(n_39), .B1(n_483), .B2(n_521), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g533 ( .A1(n_6), .A2(n_279), .B1(n_399), .B2(n_534), .C(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_7), .A2(n_140), .B1(n_625), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_7), .A2(n_150), .B1(n_598), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_8), .A2(n_58), .B1(n_1291), .B2(n_1295), .Y(n_1327) );
INVx1_ASAP7_75t_L g1183 ( .A(n_9), .Y(n_1183) );
AO22x1_ASAP7_75t_L g1208 ( .A1(n_9), .A2(n_170), .B1(n_431), .B2(n_754), .Y(n_1208) );
AND2x2_ASAP7_75t_L g358 ( .A(n_10), .B(n_246), .Y(n_358) );
AND2x2_ASAP7_75t_L g377 ( .A(n_10), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g403 ( .A(n_10), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_10), .B(n_402), .Y(n_1074) );
INVx1_ASAP7_75t_L g1191 ( .A(n_11), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_11), .A2(n_250), .B1(n_379), .B2(n_395), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_12), .A2(n_172), .B1(n_483), .B2(n_521), .C(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_12), .A2(n_74), .B1(n_600), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_13), .A2(n_188), .B1(n_367), .B2(n_632), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_13), .A2(n_18), .B1(n_400), .B2(n_708), .C(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g871 ( .A(n_14), .Y(n_871) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_14), .A2(n_163), .B1(n_421), .B2(n_607), .C(n_653), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_15), .A2(n_180), .B1(n_660), .B2(n_666), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_15), .A2(n_280), .B1(n_784), .B2(n_935), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_16), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_17), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_18), .A2(n_43), .B1(n_576), .B2(n_631), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_19), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_20), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_21), .A2(n_171), .B1(n_629), .B2(n_632), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_21), .A2(n_286), .B1(n_535), .B2(n_653), .C(n_656), .Y(n_652) );
INVx2_ASAP7_75t_L g1294 ( .A(n_22), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_22), .B(n_126), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_22), .B(n_1300), .Y(n_1302) );
INVx1_ASAP7_75t_L g685 ( .A(n_23), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_24), .A2(n_231), .B1(n_486), .B2(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g717 ( .A(n_24), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g1312 ( .A1(n_25), .A2(n_42), .B1(n_1298), .B2(n_1301), .Y(n_1312) );
XNOR2xp5_ASAP7_75t_L g1230 ( .A(n_26), .B(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g820 ( .A(n_27), .Y(n_820) );
INVx1_ASAP7_75t_L g1162 ( .A(n_28), .Y(n_1162) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_29), .A2(n_86), .B1(n_507), .B2(n_935), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_29), .A2(n_292), .B1(n_400), .B2(n_596), .C(n_828), .Y(n_1158) );
INVx1_ASAP7_75t_L g386 ( .A(n_30), .Y(n_386) );
INVx1_ASAP7_75t_L g747 ( .A(n_31), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g771 ( .A1(n_31), .A2(n_200), .B1(n_696), .B2(n_772), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_32), .A2(n_67), .B1(n_756), .B2(n_757), .C(n_759), .Y(n_755) );
INVx1_ASAP7_75t_L g786 ( .A(n_32), .Y(n_786) );
INVx1_ASAP7_75t_L g909 ( .A(n_33), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_33), .A2(n_263), .B1(n_439), .B2(n_742), .Y(n_927) );
INVx1_ASAP7_75t_L g1161 ( .A(n_34), .Y(n_1161) );
AOI22xp5_ASAP7_75t_L g1317 ( .A1(n_35), .A2(n_142), .B1(n_1298), .B2(n_1301), .Y(n_1317) );
INVx1_ASAP7_75t_L g417 ( .A(n_36), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_37), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_38), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_38), .A2(n_100), .B1(n_672), .B2(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g550 ( .A(n_39), .Y(n_550) );
NAND2xp33_ASAP7_75t_SL g508 ( .A(n_40), .B(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_40), .A2(n_94), .B1(n_537), .B2(n_540), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_41), .A2(n_292), .B1(n_507), .B2(n_935), .Y(n_1153) );
AOI22xp33_ASAP7_75t_SL g1167 ( .A1(n_41), .A2(n_86), .B1(n_659), .B2(n_667), .Y(n_1167) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_43), .A2(n_721), .B(n_722), .C(n_728), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g1014 ( .A(n_44), .B(n_399), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_44), .A2(n_191), .B1(n_506), .B2(n_805), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_45), .A2(n_137), .B1(n_336), .B2(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_46), .A2(n_191), .B1(n_431), .B2(n_539), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_46), .A2(n_264), .B1(n_631), .B2(n_805), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_47), .A2(n_112), .B1(n_1291), .B2(n_1377), .Y(n_1376) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_48), .A2(n_105), .B1(n_1291), .B2(n_1305), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_49), .A2(n_68), .B1(n_336), .B2(n_439), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_49), .A2(n_429), .B(n_706), .C(n_713), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_50), .Y(n_649) );
INVx1_ASAP7_75t_L g1128 ( .A(n_51), .Y(n_1128) );
XNOR2x2_ASAP7_75t_L g679 ( .A(n_52), .B(n_680), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g1245 ( .A1(n_53), .A2(n_828), .B(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1253 ( .A(n_53), .Y(n_1253) );
INVx1_ASAP7_75t_L g875 ( .A(n_54), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_54), .A2(n_129), .B1(n_421), .B2(n_724), .C(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g328 ( .A(n_55), .Y(n_328) );
INVx1_ASAP7_75t_L g342 ( .A(n_55), .Y(n_342) );
INVx1_ASAP7_75t_L g966 ( .A(n_56), .Y(n_966) );
AO22x1_ASAP7_75t_L g623 ( .A1(n_57), .A2(n_212), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_57), .A2(n_215), .B1(n_659), .B2(n_660), .Y(n_658) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_58), .Y(n_737) );
AND4x1_ASAP7_75t_L g788 ( .A(n_58), .B(n_739), .C(n_743), .D(n_769), .Y(n_788) );
INVx1_ASAP7_75t_L g994 ( .A(n_59), .Y(n_994) );
INVx1_ASAP7_75t_L g1135 ( .A(n_60), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_61), .A2(n_220), .B1(n_540), .B2(n_598), .Y(n_1238) );
INVx1_ASAP7_75t_L g1254 ( .A(n_61), .Y(n_1254) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_62), .A2(n_151), .B1(n_1291), .B2(n_1305), .Y(n_1323) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_63), .A2(n_75), .B1(n_523), .B2(n_525), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_63), .A2(n_75), .B1(n_375), .B2(n_411), .C(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_64), .A2(n_245), .B1(n_1298), .B2(n_1301), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_65), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_65), .A2(n_153), .B1(n_779), .B2(n_807), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_66), .A2(n_150), .B1(n_625), .B2(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_66), .A2(n_140), .B1(n_558), .B2(n_656), .C(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g787 ( .A(n_67), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g1235 ( .A1(n_69), .A2(n_255), .B1(n_400), .B2(n_606), .C(n_1236), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_69), .A2(n_294), .B1(n_331), .B2(n_935), .Y(n_1255) );
INVx2_ASAP7_75t_L g318 ( .A(n_70), .Y(n_318) );
INVx1_ASAP7_75t_L g1226 ( .A(n_71), .Y(n_1226) );
INVx1_ASAP7_75t_L g1274 ( .A(n_72), .Y(n_1274) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_73), .A2(n_279), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g547 ( .A(n_73), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_74), .A2(n_82), .B1(n_483), .B2(n_576), .C(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_76), .B(n_835), .Y(n_922) );
INVx1_ASAP7_75t_L g932 ( .A(n_76), .Y(n_932) );
XNOR2x1_ASAP7_75t_L g491 ( .A(n_77), .B(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_78), .A2(n_95), .B1(n_957), .B2(n_959), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_78), .A2(n_249), .B1(n_531), .B2(n_666), .Y(n_972) );
INVx1_ASAP7_75t_L g568 ( .A(n_79), .Y(n_568) );
INVx1_ASAP7_75t_L g874 ( .A(n_80), .Y(n_874) );
INVx1_ASAP7_75t_L g566 ( .A(n_81), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_82), .A2(n_172), .B1(n_535), .B2(n_556), .C(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g1037 ( .A(n_83), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_84), .A2(n_89), .B1(n_556), .B2(n_606), .C(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_85), .A2(n_208), .B1(n_629), .B2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_85), .A2(n_256), .B1(n_598), .B2(n_667), .Y(n_845) );
INVx1_ASAP7_75t_L g1520 ( .A(n_87), .Y(n_1520) );
AOI221xp5_ASAP7_75t_L g1531 ( .A1(n_87), .A2(n_156), .B1(n_606), .B2(n_828), .C(n_1532), .Y(n_1531) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_88), .A2(n_136), .B1(n_696), .B2(n_772), .Y(n_857) );
INVx1_ASAP7_75t_L g890 ( .A(n_88), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_89), .A2(n_271), .B1(n_580), .B2(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g872 ( .A(n_90), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_90), .A2(n_233), .B1(n_886), .B2(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g867 ( .A(n_91), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_92), .A2(n_229), .B1(n_439), .B2(n_742), .Y(n_741) );
OAI211xp5_ASAP7_75t_L g744 ( .A1(n_92), .A2(n_429), .B(n_745), .C(n_748), .Y(n_744) );
OAI222xp33_ASAP7_75t_L g1197 ( .A1(n_93), .A2(n_227), .B1(n_1111), .B2(n_1113), .C1(n_1198), .C2(n_1201), .Y(n_1197) );
INVx1_ASAP7_75t_L g1211 ( .A(n_93), .Y(n_1211) );
INVx1_ASAP7_75t_L g519 ( .A(n_94), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g982 ( .A1(n_95), .A2(n_422), .B(n_655), .Y(n_982) );
OAI22xp5_ASAP7_75t_SL g1007 ( .A1(n_96), .A2(n_119), .B1(n_1008), .B2(n_1010), .Y(n_1007) );
OAI21xp33_ASAP7_75t_L g1020 ( .A1(n_96), .A2(n_1021), .B(n_1022), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_97), .A2(n_124), .B1(n_1291), .B2(n_1295), .Y(n_1290) );
AOI22xp5_ASAP7_75t_L g1343 ( .A1(n_98), .A2(n_145), .B1(n_1298), .B2(n_1301), .Y(n_1343) );
INVx1_ASAP7_75t_L g307 ( .A(n_99), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_99), .A2(n_268), .B1(n_407), .B2(n_411), .C(n_416), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_100), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_101), .A2(n_103), .B1(n_486), .B2(n_822), .Y(n_967) );
INVx1_ASAP7_75t_L g974 ( .A(n_101), .Y(n_974) );
AOI22xp33_ASAP7_75t_SL g963 ( .A1(n_102), .A2(n_283), .B1(n_576), .B2(n_955), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g983 ( .A1(n_102), .A2(n_202), .B1(n_830), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g975 ( .A(n_103), .Y(n_975) );
CKINVDCx5p33_ASAP7_75t_R g1187 ( .A(n_104), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_106), .A2(n_285), .B1(n_667), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_106), .A2(n_132), .B1(n_777), .B2(n_779), .Y(n_780) );
INVx1_ASAP7_75t_L g334 ( .A(n_107), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_107), .A2(n_148), .B1(n_426), .B2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g1072 ( .A(n_108), .Y(n_1072) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_108), .A2(n_239), .B1(n_521), .B2(n_1096), .C(n_1098), .Y(n_1095) );
INVx1_ASAP7_75t_L g543 ( .A(n_109), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_110), .A2(n_296), .B1(n_807), .B2(n_809), .Y(n_806) );
AOI21xp33_ASAP7_75t_L g842 ( .A1(n_110), .A2(n_607), .B(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g1276 ( .A(n_111), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_111), .B(n_1274), .Y(n_1292) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_113), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_114), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_115), .Y(n_1244) );
OAI211xp5_ASAP7_75t_L g997 ( .A1(n_116), .A2(n_998), .B(n_1000), .C(n_1001), .Y(n_997) );
INVxp33_ASAP7_75t_SL g1023 ( .A(n_116), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_117), .A2(n_278), .B1(n_486), .B2(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g832 ( .A(n_117), .Y(n_832) );
INVx1_ASAP7_75t_L g489 ( .A(n_118), .Y(n_489) );
INVxp67_ASAP7_75t_SL g1043 ( .A(n_119), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g1150 ( .A(n_120), .Y(n_1150) );
INVx1_ASAP7_75t_L g1152 ( .A(n_121), .Y(n_1152) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_122), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_122), .A2(n_230), .B1(n_782), .B2(n_784), .Y(n_781) );
INVx1_ASAP7_75t_L g321 ( .A(n_123), .Y(n_321) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_123), .A2(n_373), .B(n_381), .C(n_404), .Y(n_372) );
INVxp67_ASAP7_75t_L g619 ( .A(n_124), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g1118 ( .A1(n_125), .A2(n_252), .B1(n_1119), .B2(n_1122), .Y(n_1118) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_125), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_126), .B(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1300 ( .A(n_126), .Y(n_1300) );
AOI22xp5_ASAP7_75t_L g1322 ( .A1(n_127), .A2(n_196), .B1(n_1298), .B2(n_1301), .Y(n_1322) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_128), .Y(n_740) );
INVx1_ASAP7_75t_L g863 ( .A(n_129), .Y(n_863) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_130), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_130), .A2(n_275), .B1(n_937), .B2(n_938), .Y(n_936) );
OAI211xp5_ASAP7_75t_SL g910 ( .A1(n_131), .A2(n_411), .B(n_911), .C(n_916), .Y(n_910) );
INVx1_ASAP7_75t_L g931 ( .A(n_131), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_132), .A2(n_238), .B1(n_395), .B2(n_607), .C(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g1141 ( .A(n_133), .Y(n_1141) );
AOI21xp33_ASAP7_75t_L g1166 ( .A1(n_133), .A2(n_607), .B(n_828), .Y(n_1166) );
INVx2_ASAP7_75t_L g320 ( .A(n_134), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_134), .B(n_318), .Y(n_355) );
INVx1_ASAP7_75t_L g474 ( .A(n_134), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g1522 ( .A1(n_135), .A2(n_181), .B1(n_511), .B2(n_783), .Y(n_1522) );
INVx1_ASAP7_75t_L g1533 ( .A(n_135), .Y(n_1533) );
INVx1_ASAP7_75t_L g891 ( .A(n_136), .Y(n_891) );
OAI211xp5_ASAP7_75t_L g881 ( .A1(n_137), .A2(n_825), .B(n_882), .C(n_889), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_138), .A2(n_175), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_138), .A2(n_225), .B1(n_580), .B2(n_782), .Y(n_1099) );
INVx1_ASAP7_75t_L g1083 ( .A(n_139), .Y(n_1083) );
INVx1_ASAP7_75t_L g1195 ( .A(n_141), .Y(n_1195) );
NAND2xp33_ASAP7_75t_SL g1220 ( .A(n_141), .B(n_379), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_143), .A2(n_248), .B1(n_497), .B2(n_742), .Y(n_1136) );
OAI211xp5_ASAP7_75t_L g1156 ( .A1(n_143), .A2(n_825), .B(n_1157), .C(n_1160), .Y(n_1156) );
INVx1_ASAP7_75t_L g908 ( .A(n_144), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_144), .A2(n_288), .B1(n_772), .B2(n_822), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_146), .A2(n_157), .B1(n_395), .B2(n_421), .C(n_422), .Y(n_420) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_146), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_147), .A2(n_259), .B1(n_1298), .B2(n_1301), .Y(n_1297) );
INVx1_ASAP7_75t_L g365 ( .A(n_148), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_149), .A2(n_155), .B1(n_395), .B2(n_399), .C(n_400), .Y(n_394) );
INVx1_ASAP7_75t_L g466 ( .A(n_149), .Y(n_466) );
XNOR2xp5_ASAP7_75t_L g1496 ( .A(n_151), .B(n_1497), .Y(n_1496) );
AOI22xp33_ASAP7_75t_SL g1550 ( .A1(n_151), .A2(n_1551), .B1(n_1556), .B2(n_1561), .Y(n_1550) );
AOI22xp5_ASAP7_75t_L g1342 ( .A1(n_152), .A2(n_154), .B1(n_1291), .B2(n_1295), .Y(n_1342) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_153), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_155), .A2(n_189), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_156), .A2(n_266), .B1(n_332), .B2(n_1514), .C(n_1515), .Y(n_1513) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_157), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g1557 ( .A1(n_158), .A2(n_1558), .B1(n_1559), .B2(n_1560), .Y(n_1557) );
CKINVDCx5p33_ASAP7_75t_R g1560 ( .A(n_158), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_159), .A2(n_249), .B1(n_959), .B2(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g978 ( .A(n_159), .Y(n_978) );
INVx1_ASAP7_75t_L g518 ( .A(n_160), .Y(n_518) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_161), .Y(n_801) );
OAI211xp5_ASAP7_75t_L g824 ( .A1(n_161), .A2(n_825), .B(n_826), .C(n_831), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_162), .A2(n_272), .B1(n_807), .B2(n_809), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_162), .A2(n_296), .B1(n_600), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g868 ( .A(n_163), .Y(n_868) );
INVx1_ASAP7_75t_L g393 ( .A(n_164), .Y(n_393) );
INVx1_ASAP7_75t_L g1241 ( .A(n_165), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_166), .A2(n_169), .B1(n_1298), .B2(n_1301), .Y(n_1326) );
CKINVDCx16_ASAP7_75t_R g1199 ( .A(n_167), .Y(n_1199) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_168), .A2(n_290), .B1(n_1119), .B2(n_1122), .Y(n_1504) );
INVxp33_ASAP7_75t_SL g1542 ( .A(n_168), .Y(n_1542) );
AOI21xp5_ASAP7_75t_L g1196 ( .A1(n_170), .A2(n_578), .B(n_783), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_171), .A2(n_262), .B1(n_666), .B2(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g1222 ( .A(n_173), .Y(n_1222) );
AOI22xp33_ASAP7_75t_SL g1247 ( .A1(n_174), .A2(n_294), .B1(n_431), .B2(n_659), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_174), .A2(n_255), .B1(n_521), .B2(n_935), .Y(n_1259) );
AOI22xp33_ASAP7_75t_SL g1092 ( .A1(n_175), .A2(n_273), .B1(n_809), .B2(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1240 ( .A(n_176), .Y(n_1240) );
INVx1_ASAP7_75t_L g796 ( .A(n_177), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g834 ( .A1(n_177), .A2(n_179), .B1(n_758), .B2(n_835), .C(n_836), .Y(n_834) );
BUFx3_ASAP7_75t_L g312 ( .A(n_178), .Y(n_312) );
INVx1_ASAP7_75t_L g799 ( .A(n_179), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_180), .A2(n_204), .B1(n_775), .B2(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1527 ( .A(n_181), .Y(n_1527) );
CKINVDCx5p33_ASAP7_75t_R g1507 ( .A(n_182), .Y(n_1507) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_183), .A2(n_256), .B1(n_805), .B2(n_812), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_183), .A2(n_208), .B1(n_400), .B2(n_596), .C(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1306 ( .A1(n_184), .A2(n_187), .B1(n_1298), .B2(n_1301), .Y(n_1306) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_185), .A2(n_348), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g1511 ( .A(n_186), .Y(n_1511) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_186), .A2(n_219), .B1(n_606), .B2(n_828), .C(n_1526), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_188), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_189), .Y(n_419) );
INVxp67_ASAP7_75t_L g944 ( .A(n_190), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_190), .A2(n_247), .B1(n_1291), .B2(n_1295), .Y(n_1313) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_192), .A2(n_202), .B1(n_635), .B2(n_955), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g971 ( .A1(n_192), .A2(n_283), .B1(n_395), .B2(n_400), .C(n_921), .Y(n_971) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_193), .Y(n_363) );
INVx1_ASAP7_75t_L g1499 ( .A(n_194), .Y(n_1499) );
INVx1_ASAP7_75t_L g593 ( .A(n_195), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g1508 ( .A(n_197), .Y(n_1508) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_198), .A2(n_209), .B1(n_798), .B2(n_855), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g878 ( .A1(n_198), .A2(n_209), .B1(n_756), .B2(n_757), .C(n_879), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_199), .A2(n_225), .B1(n_1051), .B2(n_1069), .C(n_1070), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1094 ( .A1(n_199), .A2(n_232), .B1(n_578), .B2(n_805), .C(n_935), .Y(n_1094) );
INVx1_ASAP7_75t_L g746 ( .A(n_200), .Y(n_746) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_201), .A2(n_497), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g1518 ( .A(n_203), .Y(n_1518) );
AOI221xp5_ASAP7_75t_L g920 ( .A1(n_204), .A2(n_280), .B1(n_400), .B2(n_750), .C(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g949 ( .A(n_205), .Y(n_949) );
OAI221xp5_ASAP7_75t_SL g976 ( .A1(n_205), .A2(n_281), .B1(n_756), .B2(n_757), .C(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g1178 ( .A(n_206), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_206), .B(n_1119), .Y(n_1180) );
XOR2x2_ASAP7_75t_L g901 ( .A(n_207), .B(n_902), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g1242 ( .A1(n_210), .A2(n_257), .B1(n_758), .B2(n_835), .C(n_1243), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1260 ( .A1(n_210), .A2(n_257), .B1(n_525), .B2(n_798), .Y(n_1260) );
INVx1_ASAP7_75t_L g542 ( .A(n_211), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_212), .B(n_663), .Y(n_662) );
AOI21xp33_ASAP7_75t_L g1017 ( .A1(n_213), .A2(n_422), .B(n_828), .Y(n_1017) );
INVx1_ASAP7_75t_L g1029 ( .A(n_213), .Y(n_1029) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_214), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_215), .A2(n_228), .B1(n_624), .B2(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_216), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_216), .A2(n_237), .B1(n_631), .B2(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_217), .A2(n_851), .B1(n_852), .B2(n_897), .Y(n_850) );
INVx1_ASAP7_75t_L g897 ( .A(n_217), .Y(n_897) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_218), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g1521 ( .A1(n_219), .A2(n_478), .B(n_1098), .Y(n_1521) );
INVx1_ASAP7_75t_L g1258 ( .A(n_220), .Y(n_1258) );
XOR2x2_ASAP7_75t_L g989 ( .A(n_221), .B(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g926 ( .A(n_222), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g702 ( .A(n_223), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_224), .A2(n_276), .B1(n_431), .B2(n_604), .Y(n_1013) );
INVx1_ASAP7_75t_L g1030 ( .A(n_224), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_226), .B(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_226), .A2(n_817), .B1(n_818), .B2(n_846), .Y(n_816) );
INVx1_ASAP7_75t_L g848 ( .A(n_226), .Y(n_848) );
NOR2xp33_ASAP7_75t_R g1213 ( .A(n_227), .B(n_1214), .Y(n_1213) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_228), .A2(n_607), .B(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_230), .A2(n_237), .B1(n_669), .B2(n_750), .C(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g714 ( .A(n_231), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_232), .A2(n_239), .B1(n_1053), .B2(n_1055), .C(n_1057), .Y(n_1052) );
INVx1_ASAP7_75t_L g862 ( .A(n_233), .Y(n_862) );
INVx1_ASAP7_75t_L g684 ( .A(n_234), .Y(n_684) );
INVx1_ASAP7_75t_L g1173 ( .A(n_235), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_236), .A2(n_293), .B1(n_497), .B2(n_742), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_238), .A2(n_285), .B1(n_777), .B2(n_779), .Y(n_776) );
INVxp67_ASAP7_75t_SL g1086 ( .A(n_240), .Y(n_1086) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_240), .A2(n_243), .B1(n_1111), .B2(n_1113), .C(n_1115), .Y(n_1110) );
INVx1_ASAP7_75t_L g1262 ( .A(n_241), .Y(n_1262) );
OAI211xp5_ASAP7_75t_SL g1505 ( .A1(n_242), .A2(n_1108), .B(n_1115), .C(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1538 ( .A(n_242), .Y(n_1538) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_243), .A2(n_254), .B1(n_1060), .B2(n_1065), .C(n_1066), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_244), .Y(n_1003) );
INVx1_ASAP7_75t_L g378 ( .A(n_246), .Y(n_378) );
BUFx3_ASAP7_75t_L g402 ( .A(n_246), .Y(n_402) );
INVx1_ASAP7_75t_L g1188 ( .A(n_250), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_251), .Y(n_642) );
INVxp67_ASAP7_75t_SL g1079 ( .A(n_252), .Y(n_1079) );
OAI21xp5_ASAP7_75t_SL g675 ( .A1(n_253), .A2(n_439), .B(n_676), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_254), .A2(n_258), .B1(n_1101), .B2(n_1104), .Y(n_1100) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_258), .Y(n_1088) );
INVx1_ASAP7_75t_L g315 ( .A(n_260), .Y(n_315) );
INVx1_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
INVx2_ASAP7_75t_L g436 ( .A(n_260), .Y(n_436) );
XNOR2x1_ASAP7_75t_L g563 ( .A(n_261), .B(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_262), .A2(n_286), .B1(n_631), .B2(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g1012 ( .A(n_264), .B(n_828), .Y(n_1012) );
INVx1_ASAP7_75t_L g1185 ( .A(n_265), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_265), .A2(n_295), .B1(n_540), .B2(n_754), .Y(n_1219) );
INVx1_ASAP7_75t_L g1528 ( .A(n_266), .Y(n_1528) );
OR2x2_ASAP7_75t_L g347 ( .A(n_267), .B(n_348), .Y(n_347) );
OAI322xp33_ASAP7_75t_L g449 ( .A1(n_268), .A2(n_450), .A3(n_458), .B1(n_461), .B2(n_469), .C1(n_475), .C2(n_486), .Y(n_449) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_269), .Y(n_952) );
OAI211xp5_ASAP7_75t_SL g969 ( .A1(n_269), .A2(n_429), .B(n_970), .C(n_973), .Y(n_969) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_270), .Y(n_894) );
INVx1_ASAP7_75t_L g837 ( .A(n_272), .Y(n_837) );
INVx1_ASAP7_75t_L g1071 ( .A(n_273), .Y(n_1071) );
INVx1_ASAP7_75t_L g495 ( .A(n_274), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_275), .A2(n_422), .B(n_653), .Y(n_915) );
INVxp67_ASAP7_75t_SL g1034 ( .A(n_276), .Y(n_1034) );
OAI22xp33_ASAP7_75t_SL g1154 ( .A1(n_277), .A2(n_287), .B1(n_525), .B2(n_798), .Y(n_1154) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_277), .A2(n_287), .B1(n_756), .B2(n_758), .C(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g833 ( .A(n_278), .Y(n_833) );
INVx1_ASAP7_75t_L g950 ( .A(n_281), .Y(n_950) );
XNOR2xp5_ASAP7_75t_L g1132 ( .A(n_282), .B(n_1133), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_284), .Y(n_1512) );
INVx1_ASAP7_75t_L g906 ( .A(n_288), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_289), .Y(n_1002) );
INVxp67_ASAP7_75t_SL g1502 ( .A(n_290), .Y(n_1502) );
INVx1_ASAP7_75t_L g1016 ( .A(n_291), .Y(n_1016) );
OAI211xp5_ASAP7_75t_L g1233 ( .A1(n_293), .A2(n_825), .B(n_1234), .C(n_1239), .Y(n_1233) );
INVx1_ASAP7_75t_L g1192 ( .A(n_295), .Y(n_1192) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_1268), .B(n_1284), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_898), .B1(n_1266), .B2(n_1267), .Y(n_298) );
INVxp67_ASAP7_75t_SL g1266 ( .A(n_299), .Y(n_1266) );
XOR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_734), .Y(n_299) );
XOR2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_616), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_490), .B2(n_615), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
XNOR2x1_ASAP7_75t_L g303 ( .A(n_304), .B(n_489), .Y(n_303) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_305), .B(n_370), .Y(n_304) );
NAND5xp2_ASAP7_75t_L g305 ( .A(n_306), .B(n_329), .C(n_333), .D(n_347), .E(n_364), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_321), .B2(n_322), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_308), .A2(n_322), .B1(n_644), .B2(n_645), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_308), .A2(n_322), .B1(n_684), .B2(n_685), .Y(n_683) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .Y(n_308) );
AND2x2_ASAP7_75t_L g524 ( .A(n_309), .B(n_313), .Y(n_524) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_309), .B(n_313), .Y(n_572) );
NAND2x1_ASAP7_75t_L g798 ( .A(n_309), .B(n_313), .Y(n_798) );
AND2x6_ASAP7_75t_L g1112 ( .A(n_309), .B(n_316), .Y(n_1112) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_311), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g511 ( .A(n_311), .B(n_326), .Y(n_511) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g332 ( .A(n_312), .B(n_327), .Y(n_332) );
INVx2_ASAP7_75t_L g339 ( .A(n_312), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_312), .B(n_328), .Y(n_352) );
OR2x2_ASAP7_75t_L g465 ( .A(n_312), .B(n_341), .Y(n_465) );
AND2x4_ASAP7_75t_L g322 ( .A(n_313), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g330 ( .A(n_313), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_SL g526 ( .A(n_313), .B(n_323), .Y(n_526) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
OR2x2_ASAP7_75t_L g356 ( .A(n_314), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g1077 ( .A(n_314), .Y(n_1077) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g473 ( .A(n_315), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_315), .B(n_377), .Y(n_1082) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_316), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_316), .B(n_325), .Y(n_1114) );
INVx1_ASAP7_75t_L g1117 ( .A(n_316), .Y(n_1117) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
NAND3x1_ASAP7_75t_L g472 ( .A(n_317), .B(n_473), .C(n_474), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_317), .B(n_474), .Y(n_578) );
INVx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp33_ASAP7_75t_SL g460 ( .A(n_318), .B(n_320), .Y(n_460) );
BUFx3_ASAP7_75t_L g585 ( .A(n_318), .Y(n_585) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND3x4_ASAP7_75t_L g584 ( .A(n_320), .B(n_585), .C(n_586), .Y(n_584) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_320), .B(n_585), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_322), .A2(n_524), .B1(n_786), .B2(n_787), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_322), .A2(n_796), .B1(n_797), .B2(n_799), .Y(n_795) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_322), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_322), .A2(n_524), .B1(n_931), .B2(n_932), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_322), .A2(n_524), .B1(n_949), .B2(n_950), .Y(n_948) );
AOI221x1_ASAP7_75t_L g1026 ( .A1(n_322), .A2(n_797), .B1(n_994), .B2(n_1002), .C(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g447 ( .A(n_328), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g569 ( .A(n_329), .B(n_570), .C(n_574), .Y(n_569) );
AND4x1_ASAP7_75t_L g769 ( .A(n_329), .B(n_770), .C(n_773), .D(n_785), .Y(n_769) );
INVx2_ASAP7_75t_SL g876 ( .A(n_329), .Y(n_876) );
AND5x1_ASAP7_75t_L g990 ( .A(n_329), .B(n_991), .C(n_1026), .D(n_1036), .E(n_1042), .Y(n_990) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR3xp33_ASAP7_75t_SL g499 ( .A(n_330), .B(n_500), .C(n_522), .Y(n_499) );
INVx3_ASAP7_75t_L g640 ( .A(n_330), .Y(n_640) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_330), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g1249 ( .A(n_330), .B(n_1250), .C(n_1260), .Y(n_1249) );
BUFx2_ASAP7_75t_L g632 ( .A(n_331), .Y(n_632) );
BUFx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g485 ( .A(n_332), .Y(n_485) );
BUFx2_ASAP7_75t_L g507 ( .A(n_332), .Y(n_507) );
BUFx2_ASAP7_75t_L g576 ( .A(n_332), .Y(n_576) );
BUFx2_ASAP7_75t_L g775 ( .A(n_332), .Y(n_775) );
BUFx3_ASAP7_75t_L g805 ( .A(n_332), .Y(n_805) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_332), .B(n_1103), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_335), .A2(n_495), .B1(n_496), .B2(n_498), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_335), .A2(n_566), .B1(n_567), .B2(n_568), .C(n_569), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_335), .B(n_642), .Y(n_641) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx5_ASAP7_75t_L g802 ( .A(n_336), .Y(n_802) );
OR2x6_ASAP7_75t_L g336 ( .A(n_337), .B(n_343), .Y(n_336) );
OR2x2_ASAP7_75t_L g742 ( .A(n_337), .B(n_343), .Y(n_742) );
INVx2_ASAP7_75t_L g1109 ( .A(n_337), .Y(n_1109) );
INVx8_ASAP7_75t_L g368 ( .A(n_338), .Y(n_368) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_338), .Y(n_506) );
BUFx3_ASAP7_75t_L g631 ( .A(n_338), .Y(n_631) );
BUFx3_ASAP7_75t_L g783 ( .A(n_338), .Y(n_783) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_338), .B(n_1103), .Y(n_1102) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x4_ASAP7_75t_L g454 ( .A(n_339), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g455 ( .A(n_342), .Y(n_455) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g440 ( .A(n_344), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g1041 ( .A(n_344), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_344), .B(n_441), .Y(n_1065) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g354 ( .A(n_345), .Y(n_354) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx8_ASAP7_75t_L g567 ( .A(n_348), .Y(n_567) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_356), .Y(n_348) );
INVx1_ASAP7_75t_L g1024 ( .A(n_349), .Y(n_1024) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
BUFx3_ASAP7_75t_L g1033 ( .A(n_350), .Y(n_1033) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_351), .Y(n_457) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g481 ( .A(n_352), .Y(n_481) );
INVx1_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
OR2x2_ASAP7_75t_L g444 ( .A(n_353), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g614 ( .A(n_353), .Y(n_614) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g459 ( .A(n_354), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_SL g1058 ( .A(n_354), .B(n_401), .Y(n_1058) );
INVx1_ASAP7_75t_L g1536 ( .A(n_354), .Y(n_1536) );
INVx1_ASAP7_75t_L g1103 ( .A(n_355), .Y(n_1103) );
INVx1_ASAP7_75t_L g1121 ( .A(n_355), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_356), .B(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1078 ( .A(n_357), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x6_ASAP7_75t_L g405 ( .A(n_358), .B(n_379), .Y(n_405) );
INVx1_ASAP7_75t_L g415 ( .A(n_358), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_358), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g608 ( .A(n_358), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_358), .B(n_436), .Y(n_1062) );
AND2x2_ASAP7_75t_L g428 ( .A(n_359), .B(n_377), .Y(n_428) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_359), .Y(n_539) );
INVx3_ASAP7_75t_L g599 ( .A(n_359), .Y(n_599) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_360), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_360), .B(n_363), .Y(n_1009) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g380 ( .A(n_361), .B(n_363), .Y(n_380) );
OR2x2_ASAP7_75t_L g385 ( .A(n_361), .B(n_363), .Y(n_385) );
INVx2_ASAP7_75t_L g392 ( .A(n_361), .Y(n_392) );
AND2x2_ASAP7_75t_L g397 ( .A(n_361), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g443 ( .A(n_361), .Y(n_443) );
NAND2x1_ASAP7_75t_L g841 ( .A(n_361), .B(n_363), .Y(n_841) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_363), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
BUFx2_ASAP7_75t_L g414 ( .A(n_363), .Y(n_414) );
AND2x2_ASAP7_75t_L g432 ( .A(n_363), .B(n_392), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_366), .A2(n_542), .B1(n_543), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_366), .A2(n_487), .B1(n_649), .B2(n_650), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_366), .A2(n_487), .B1(n_1161), .B2(n_1162), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_366), .A2(n_487), .B1(n_1240), .B2(n_1241), .Y(n_1264) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
AND2x4_ASAP7_75t_L g612 ( .A(n_367), .B(n_369), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_367), .A2(n_1177), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g483 ( .A(n_368), .Y(n_483) );
INVx3_ASAP7_75t_L g812 ( .A(n_368), .Y(n_812) );
INVx8_ASAP7_75t_L g935 ( .A(n_368), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_368), .Y(n_1514) );
AND2x4_ASAP7_75t_L g487 ( .A(n_369), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_437), .Y(n_370) );
OAI31xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_406), .A3(n_425), .B(n_433), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_374), .A2(n_412), .B1(n_684), .B2(n_685), .Y(n_728) );
INVx2_ASAP7_75t_L g756 ( .A(n_374), .Y(n_756) );
INVx2_ASAP7_75t_L g835 ( .A(n_374), .Y(n_835) );
INVx4_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g602 ( .A(n_376), .Y(n_602) );
AND2x4_ASAP7_75t_SL g376 ( .A(n_377), .B(n_379), .Y(n_376) );
AND2x4_ASAP7_75t_L g409 ( .A(n_377), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g430 ( .A(n_377), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g530 ( .A(n_377), .B(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_377), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_377), .B(n_410), .Y(n_1127) );
BUFx3_ASAP7_75t_L g399 ( .A(n_379), .Y(n_399) );
BUFx3_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_379), .Y(n_596) );
BUFx3_ASAP7_75t_L g606 ( .A(n_379), .Y(n_606) );
INVx1_ASAP7_75t_L g670 ( .A(n_379), .Y(n_670) );
BUFx3_ASAP7_75t_L g921 ( .A(n_379), .Y(n_921) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g555 ( .A(n_380), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_386), .B1(n_387), .B2(n_393), .C(n_394), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_382), .A2(n_417), .B1(n_418), .B2(n_419), .C(n_420), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g879 ( .A1(n_382), .A2(n_763), .B1(n_867), .B2(n_874), .C(n_880), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_382), .A2(n_917), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_916) );
INVx1_ASAP7_75t_L g1051 ( .A(n_382), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g546 ( .A(n_383), .Y(n_546) );
INVx2_ASAP7_75t_SL g761 ( .A(n_383), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_383), .A2(n_1527), .B1(n_1528), .B2(n_1529), .Y(n_1526) );
OAI22x1_ASAP7_75t_SL g1532 ( .A1(n_383), .A2(n_1512), .B1(n_1529), .B2(n_1533), .Y(n_1532) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g727 ( .A(n_384), .Y(n_727) );
BUFx4f_ASAP7_75t_L g999 ( .A(n_384), .Y(n_999) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_386), .A2(n_451), .B1(n_452), .B2(n_456), .Y(n_450) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_388), .Y(n_918) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g549 ( .A(n_389), .Y(n_549) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_389), .Y(n_721) );
INVx2_ASAP7_75t_L g765 ( .A(n_389), .Y(n_765) );
INVx4_ASAP7_75t_L g1010 ( .A(n_389), .Y(n_1010) );
INVx2_ASAP7_75t_L g1529 ( .A(n_389), .Y(n_1529) );
INVx8_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g418 ( .A(n_390), .Y(n_418) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g475 ( .A1(n_393), .A2(n_476), .B1(n_479), .B2(n_480), .C(n_482), .Y(n_475) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g655 ( .A(n_396), .Y(n_655) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_397), .Y(n_410) );
BUFx3_ASAP7_75t_L g828 ( .A(n_397), .Y(n_828) );
HB1xp67_ASAP7_75t_SL g884 ( .A(n_400), .Y(n_884) );
INVx4_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx4_ASAP7_75t_L g535 ( .A(n_401), .Y(n_535) );
INVx1_ASAP7_75t_SL g752 ( .A(n_401), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g1011 ( .A(n_401), .B(n_1012), .C(n_1013), .D(n_1014), .Y(n_1011) );
AND2x4_ASAP7_75t_L g1534 ( .A(n_401), .B(n_1535), .Y(n_1534) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
AND2x4_ASAP7_75t_L g423 ( .A(n_403), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g1280 ( .A(n_403), .Y(n_1280) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_405), .A2(n_498), .B1(n_530), .B2(n_533), .C(n_536), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_405), .A2(n_530), .B1(n_566), .B2(n_595), .C(n_597), .Y(n_594) );
AOI221xp5_ASAP7_75t_SL g651 ( .A1(n_405), .A2(n_430), .B1(n_642), .B2(n_652), .C(n_658), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_405), .A2(n_707), .B(n_711), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_405), .A2(n_749), .B(n_753), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_405), .A2(n_827), .B(n_829), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_405), .A2(n_883), .B(n_885), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_405), .A2(n_408), .B(n_906), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g970 ( .A1(n_405), .A2(n_971), .B(n_972), .Y(n_970) );
AOI21xp5_ASAP7_75t_L g1157 ( .A1(n_405), .A2(n_1158), .B(n_1159), .Y(n_1157) );
AOI21xp5_ASAP7_75t_L g1234 ( .A1(n_405), .A2(n_1235), .B(n_1238), .Y(n_1234) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_408), .A2(n_427), .B1(n_746), .B2(n_747), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_408), .A2(n_427), .B1(n_974), .B2(n_975), .Y(n_973) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_409), .A2(n_427), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_409), .A2(n_427), .B1(n_592), .B2(n_593), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_409), .A2(n_427), .B1(n_649), .B2(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g719 ( .A(n_409), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_409), .A2(n_427), .B1(n_832), .B2(n_833), .Y(n_831) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_409), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_409), .A2(n_427), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_409), .A2(n_428), .B1(n_1240), .B2(n_1241), .Y(n_1239) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_410), .Y(n_534) );
INVx2_ASAP7_75t_L g557 ( .A(n_410), .Y(n_557) );
INVx1_ASAP7_75t_L g1237 ( .A(n_410), .Y(n_1237) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g758 ( .A(n_412), .Y(n_758) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g609 ( .A(n_414), .Y(n_609) );
INVx1_ASAP7_75t_L g1064 ( .A(n_414), .Y(n_1064) );
INVx1_ASAP7_75t_L g996 ( .A(n_415), .Y(n_996) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_417), .A2(n_462), .B1(n_466), .B2(n_467), .Y(n_461) );
INVx1_ASAP7_75t_L g1069 ( .A(n_418), .Y(n_1069) );
INVx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g558 ( .A(n_423), .Y(n_558) );
INVx2_ASAP7_75t_L g607 ( .A(n_423), .Y(n_607) );
INVx1_ASAP7_75t_L g1246 ( .A(n_423), .Y(n_1246) );
INVxp67_ASAP7_75t_L g1283 ( .A(n_424), .Y(n_1283) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_427), .A2(n_430), .B1(n_908), .B2(n_909), .Y(n_907) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g716 ( .A(n_428), .Y(n_716) );
AND2x4_ASAP7_75t_L g1040 ( .A(n_428), .B(n_1041), .Y(n_1040) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g825 ( .A(n_430), .Y(n_825) );
BUFx2_ASAP7_75t_L g660 ( .A(n_431), .Y(n_660) );
INVx1_ASAP7_75t_L g985 ( .A(n_431), .Y(n_985) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g532 ( .A(n_432), .Y(n_532) );
BUFx3_ASAP7_75t_L g540 ( .A(n_432), .Y(n_540) );
BUFx3_ASAP7_75t_L g600 ( .A(n_432), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g743 ( .A1(n_433), .A2(n_744), .B(n_755), .Y(n_743) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g560 ( .A(n_434), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_434), .B(n_1123), .Y(n_1228) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g577 ( .A(n_435), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g1073 ( .A(n_435), .B(n_1074), .Y(n_1073) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g586 ( .A(n_436), .Y(n_586) );
AOI21xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_448), .B(n_449), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_438), .A2(n_820), .B(n_821), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_438), .A2(n_966), .B(n_967), .Y(n_965) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_439), .Y(n_896) );
AND2x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_444), .Y(n_439) );
AND2x4_ASAP7_75t_L g497 ( .A(n_440), .B(n_444), .Y(n_497) );
INVx2_ASAP7_75t_SL g1540 ( .A(n_440), .Y(n_1540) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g1025 ( .A(n_444), .Y(n_1025) );
INVx3_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_446), .Y(n_1116) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_453), .Y(n_581) );
INVx2_ASAP7_75t_L g778 ( .A(n_453), .Y(n_778) );
INVx2_ASAP7_75t_L g1149 ( .A(n_453), .Y(n_1149) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_454), .Y(n_478) );
BUFx8_ASAP7_75t_L g488 ( .A(n_454), .Y(n_488) );
INVx2_ASAP7_75t_L g517 ( .A(n_454), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g1028 ( .A1(n_456), .A2(n_504), .B1(n_1029), .B2(n_1030), .C(n_1031), .Y(n_1028) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g861 ( .A(n_457), .Y(n_861) );
CKINVDCx8_ASAP7_75t_R g1151 ( .A(n_457), .Y(n_1151) );
INVx3_ASAP7_75t_L g1184 ( .A(n_457), .Y(n_1184) );
OAI22xp5_ASAP7_75t_SL g1027 ( .A1(n_458), .A2(n_512), .B1(n_1028), .B2(n_1032), .Y(n_1027) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx4f_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
BUFx8_ASAP7_75t_L g859 ( .A(n_459), .Y(n_859) );
BUFx4f_ASAP7_75t_L g1139 ( .A(n_459), .Y(n_1139) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_460), .Y(n_1098) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_464), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1182) );
BUFx4f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g698 ( .A(n_465), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g860 ( .A1(n_467), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_467), .A2(n_865), .B1(n_874), .B2(n_875), .Y(n_873) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g1194 ( .A(n_468), .Y(n_1194) );
OAI33xp33_ASAP7_75t_L g858 ( .A1(n_469), .A2(n_859), .A3(n_860), .B1(n_864), .B2(n_869), .B3(n_873), .Y(n_858) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_470), .B(n_634), .C(n_637), .Y(n_633) );
AOI33xp33_ASAP7_75t_L g773 ( .A1(n_470), .A2(n_584), .A3(n_774), .B1(n_776), .B2(n_780), .B3(n_781), .Y(n_773) );
BUFx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g693 ( .A(n_471), .Y(n_693) );
BUFx2_ASAP7_75t_L g813 ( .A(n_471), .Y(n_813) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g513 ( .A(n_472), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_476), .A2(n_865), .B1(n_867), .B2(n_868), .Y(n_864) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx8_ASAP7_75t_L g692 ( .A(n_477), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g1032 ( .A1(n_477), .A2(n_1016), .B1(n_1033), .B2(n_1034), .C(n_1035), .Y(n_1032) );
INVx5_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g504 ( .A(n_478), .Y(n_504) );
INVx2_ASAP7_75t_SL g808 ( .A(n_478), .Y(n_808) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_478), .Y(n_937) );
INVx3_ASAP7_75t_L g1097 ( .A(n_478), .Y(n_1097) );
OAI221xp5_ASAP7_75t_L g514 ( .A1(n_480), .A2(n_515), .B1(n_518), .B2(n_519), .C(n_520), .Y(n_514) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g1144 ( .A(n_481), .Y(n_1144) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
INVx1_ASAP7_75t_L g784 ( .A(n_485), .Y(n_784) );
INVx2_ASAP7_75t_L g1200 ( .A(n_485), .Y(n_1200) );
INVxp67_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g772 ( .A(n_487), .Y(n_772) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_488), .Y(n_624) );
INVx2_ASAP7_75t_SL g870 ( .A(n_488), .Y(n_870) );
INVx3_ASAP7_75t_L g962 ( .A(n_488), .Y(n_962) );
INVx2_ASAP7_75t_SL g1252 ( .A(n_488), .Y(n_1252) );
INVx1_ASAP7_75t_L g615 ( .A(n_490), .Y(n_615) );
XNOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_563), .Y(n_490) );
NAND4xp75_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .C(n_527), .D(n_561), .Y(n_492) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_512), .B2(n_514), .Y(n_500) );
OAI211xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_505), .C(n_508), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_504), .A2(n_861), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_R g938 ( .A(n_510), .Y(n_938) );
INVx1_ASAP7_75t_L g959 ( .A(n_510), .Y(n_959) );
INVx5_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx12f_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
BUFx3_ASAP7_75t_L g625 ( .A(n_511), .Y(n_625) );
BUFx3_ASAP7_75t_L g779 ( .A(n_511), .Y(n_779) );
BUFx2_ASAP7_75t_L g809 ( .A(n_511), .Y(n_809) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_511), .B(n_1121), .Y(n_1123) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI33xp33_ASAP7_75t_L g953 ( .A1(n_513), .A2(n_627), .A3(n_954), .B1(n_956), .B2(n_960), .B3(n_963), .Y(n_953) );
INVx2_ASAP7_75t_L g1147 ( .A(n_513), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g1256 ( .A(n_513), .Y(n_1256) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g613 ( .A(n_516), .B(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g690 ( .A(n_517), .Y(n_690) );
BUFx2_ASAP7_75t_L g958 ( .A(n_517), .Y(n_958) );
INVx1_ASAP7_75t_L g1093 ( .A(n_517), .Y(n_1093) );
OR2x6_ASAP7_75t_SL g1119 ( .A(n_517), .B(n_1120), .Y(n_1119) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_517), .A2(n_1141), .B1(n_1142), .B2(n_1145), .C(n_1146), .Y(n_1140) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_526), .A2(n_571), .B1(n_572), .B2(n_573), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_544), .B(n_559), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_541), .Y(n_528) );
AND2x4_ASAP7_75t_L g1080 ( .A(n_531), .B(n_1081), .Y(n_1080) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g667 ( .A(n_532), .Y(n_667) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g666 ( .A(n_538), .Y(n_666) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g830 ( .A(n_539), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_548), .B2(n_550), .C(n_551), .Y(n_545) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g657 ( .A(n_555), .Y(n_657) );
INVx1_ASAP7_75t_L g710 ( .A(n_556), .Y(n_710) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g664 ( .A(n_557), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g968 ( .A1(n_559), .A2(n_969), .B(n_976), .Y(n_968) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g589 ( .A(n_560), .Y(n_589) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_588), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_567), .B(n_678), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_567), .A2(n_702), .B(n_703), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g739 ( .A1(n_567), .A2(n_740), .B(n_741), .Y(n_739) );
NAND2xp33_ASAP7_75t_L g814 ( .A(n_567), .B(n_815), .Y(n_814) );
AOI21xp33_ASAP7_75t_L g893 ( .A1(n_567), .A2(n_894), .B(n_895), .Y(n_893) );
AOI21xp33_ASAP7_75t_SL g925 ( .A1(n_567), .A2(n_926), .B(n_927), .Y(n_925) );
AOI211x1_ASAP7_75t_L g945 ( .A1(n_567), .A2(n_946), .B(n_947), .C(n_964), .Y(n_945) );
AOI21xp5_ASAP7_75t_L g1134 ( .A1(n_567), .A2(n_1135), .B(n_1136), .Y(n_1134) );
AOI21xp5_ASAP7_75t_L g1261 ( .A1(n_567), .A2(n_1262), .B(n_1263), .Y(n_1261) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_571), .A2(n_573), .B1(n_602), .B2(n_603), .C1(n_605), .C2(n_608), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_579), .B1(n_582), .B2(n_587), .Y(n_574) );
INVx1_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
INVx3_ASAP7_75t_L g1516 ( .A(n_578), .Y(n_1516) );
BUFx2_ASAP7_75t_L g638 ( .A(n_580), .Y(n_638) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g627 ( .A(n_584), .Y(n_627) );
AOI33xp33_ASAP7_75t_L g803 ( .A1(n_584), .A2(n_804), .A3(n_806), .B1(n_810), .B2(n_811), .B3(n_813), .Y(n_803) );
AOI33xp33_ASAP7_75t_L g933 ( .A1(n_584), .A2(n_693), .A3(n_934), .B1(n_936), .B2(n_939), .B3(n_940), .Y(n_933) );
INVx2_ASAP7_75t_SL g674 ( .A(n_586), .Y(n_674) );
INVx1_ASAP7_75t_L g732 ( .A(n_586), .Y(n_732) );
OAI31xp33_ASAP7_75t_L g1179 ( .A1(n_586), .A2(n_1180), .A3(n_1181), .B(n_1197), .Y(n_1179) );
OAI31xp33_ASAP7_75t_SL g1503 ( .A1(n_586), .A2(n_1504), .A3(n_1505), .B(n_1509), .Y(n_1503) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_610), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_589), .A2(n_824), .B(n_834), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g1155 ( .A1(n_589), .A2(n_1156), .B(n_1163), .Y(n_1155) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .C(n_601), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_592), .A2(n_593), .B1(n_612), .B2(n_613), .Y(n_611) );
BUFx2_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g604 ( .A(n_599), .Y(n_604) );
INVx2_ASAP7_75t_SL g659 ( .A(n_599), .Y(n_659) );
INVx2_ASAP7_75t_L g754 ( .A(n_599), .Y(n_754) );
INVx1_ASAP7_75t_L g886 ( .A(n_599), .Y(n_886) );
BUFx3_ASAP7_75t_L g712 ( .A(n_600), .Y(n_712) );
INVx1_ASAP7_75t_SL g888 ( .A(n_600), .Y(n_888) );
INVx1_ASAP7_75t_L g672 ( .A(n_602), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_602), .B(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g673 ( .A(n_608), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_609), .A2(n_1002), .B1(n_1003), .B2(n_1004), .Y(n_1001) );
INVx2_ASAP7_75t_SL g1021 ( .A(n_613), .Y(n_1021) );
INVxp67_ASAP7_75t_L g699 ( .A(n_614), .Y(n_699) );
OAI22x1_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_679), .B2(n_733), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
XNOR2x1_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND3x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_646), .C(n_677), .Y(n_620) );
NOR2xp33_ASAP7_75t_SL g621 ( .A(n_622), .B(n_639), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_626), .B(n_633), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AOI33xp33_ASAP7_75t_L g686 ( .A1(n_627), .A2(n_687), .A3(n_688), .B1(n_691), .B2(n_693), .B3(n_694), .Y(n_686) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .C(n_643), .Y(n_639) );
NAND4xp25_ASAP7_75t_SL g794 ( .A(n_640), .B(n_795), .C(n_800), .D(n_803), .Y(n_794) );
INVx1_ASAP7_75t_L g942 ( .A(n_640), .Y(n_942) );
NAND4xp25_ASAP7_75t_SL g947 ( .A(n_640), .B(n_948), .C(n_951), .D(n_953), .Y(n_947) );
AOI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_674), .B(n_675), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_651), .C(n_661), .Y(n_647) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_655), .Y(n_724) );
INVx1_ASAP7_75t_L g751 ( .A(n_655), .Y(n_751) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI31xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .A3(n_668), .B(n_671), .Y(n_661) );
BUFx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g768 ( .A(n_670), .Y(n_768) );
INVx1_ASAP7_75t_L g733 ( .A(n_679), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_701), .C(n_704), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_695), .C(n_700), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_686), .Y(n_682) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_696), .B(n_1039), .Y(n_1038) );
OR2x6_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
OR2x2_ASAP7_75t_L g822 ( .A(n_697), .B(n_699), .Y(n_822) );
INVx2_ASAP7_75t_SL g866 ( .A(n_697), .Y(n_866) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g1137 ( .A(n_700), .B(n_1138), .C(n_1154), .Y(n_1137) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_720), .B(n_729), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_717), .B2(n_718), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_715), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_889) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OR2x6_ASAP7_75t_L g1282 ( .A(n_727), .B(n_1283), .Y(n_1282) );
OAI21xp5_ASAP7_75t_L g877 ( .A1(n_729), .A2(n_878), .B(n_881), .Y(n_877) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g924 ( .A(n_731), .Y(n_924) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_731), .Y(n_1019) );
A2O1A1Ixp33_ASAP7_75t_L g1090 ( .A1(n_731), .A2(n_1091), .B(n_1106), .C(n_1124), .Y(n_1090) );
BUFx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_732), .Y(n_1248) );
XNOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_850), .Y(n_734) );
OAI22x1_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_789), .B1(n_790), .B2(n_849), .Y(n_735) );
INVx2_ASAP7_75t_L g849 ( .A(n_736), .Y(n_849) );
AO21x2_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_788), .Y(n_736) );
NAND3xp33_ASAP7_75t_SL g738 ( .A(n_739), .B(n_743), .C(n_769), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_742), .B(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_762), .B1(n_763), .B2(n_766), .C(n_767), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g1050 ( .A(n_764), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_791), .B(n_816), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_814), .Y(n_792) );
INVxp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_SL g846 ( .A(n_794), .B(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_802), .B(n_952), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_802), .B(n_1043), .Y(n_1042) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_814), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_823), .Y(n_818) );
INVx1_ASAP7_75t_L g844 ( .A(n_828), .Y(n_844) );
OAI211xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B(n_842), .C(n_845), .Y(n_836) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g1000 ( .A(n_839), .Y(n_1000) );
INVx1_ASAP7_75t_L g1165 ( .A(n_839), .Y(n_1165) );
INVx4_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx4f_ASAP7_75t_L g913 ( .A(n_840), .Y(n_913) );
BUFx4f_ASAP7_75t_L g1056 ( .A(n_840), .Y(n_1056) );
OR2x6_ASAP7_75t_L g1066 ( .A(n_840), .B(n_1067), .Y(n_1066) );
BUFx6f_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
BUFx3_ASAP7_75t_L g981 ( .A(n_841), .Y(n_981) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
AND3x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_877), .C(n_893), .Y(n_852) );
NOR4xp25_ASAP7_75t_L g853 ( .A(n_854), .B(n_857), .C(n_858), .D(n_876), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI22xp5_ASAP7_75t_SL g1250 ( .A1(n_859), .A2(n_1251), .B1(n_1256), .B2(n_1257), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_861), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_SL g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g1267 ( .A(n_898), .Y(n_1267) );
XNOR2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_1169), .Y(n_898) );
XNOR2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_986), .Y(n_899) );
XNOR2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_943), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_925), .C(n_928), .Y(n_902) );
OAI31xp33_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_910), .A3(n_922), .B(n_923), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_905), .B(n_907), .Y(n_904) );
OAI211xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B(n_914), .C(n_915), .Y(n_911) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
NOR3xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_941), .C(n_942), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_933), .Y(n_929) );
BUFx2_ASAP7_75t_L g955 ( .A(n_935), .Y(n_955) );
XNOR2x2_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_968), .Y(n_964) );
OAI211xp5_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_979), .B(n_982), .C(n_983), .Y(n_977) );
OAI211xp5_ASAP7_75t_L g1015 ( .A1(n_979), .A2(n_1016), .B(n_1017), .C(n_1018), .Y(n_1015) );
OAI211xp5_ASAP7_75t_L g1243 ( .A1(n_979), .A2(n_1244), .B(n_1245), .C(n_1247), .Y(n_1243) );
INVx5_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx2_ASAP7_75t_SL g980 ( .A(n_981), .Y(n_980) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_981), .B(n_1082), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_981), .B(n_1082), .Y(n_1214) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
XNOR2xp5_ASAP7_75t_L g986 ( .A(n_987), .B(n_1130), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B1(n_1044), .B2(n_1129), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_1019), .B(n_1020), .Y(n_991) );
NAND4xp25_ASAP7_75t_L g992 ( .A(n_993), .B(n_995), .C(n_1011), .D(n_1015), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_997), .B1(n_1006), .B2(n_1007), .Y(n_995) );
INVx4_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_1003), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_1009), .Y(n_1054) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1009), .Y(n_1218) );
OAI221xp5_ASAP7_75t_L g1510 ( .A1(n_1033), .A2(n_1097), .B1(n_1511), .B2(n_1512), .C(n_1513), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1039), .Y(n_1089) );
INVx3_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_1040), .A2(n_1126), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1498 ( .A(n_1040), .Y(n_1498) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1041), .B(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1044), .Y(n_1129) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
XNOR2x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1128), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1090), .Y(n_1046) );
NAND3xp33_ASAP7_75t_SL g1047 ( .A(n_1048), .B(n_1075), .C(n_1087), .Y(n_1047) );
AOI211xp5_ASAP7_75t_SL g1048 ( .A1(n_1049), .A2(n_1052), .B(n_1059), .C(n_1068), .Y(n_1048) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_1054), .A2(n_1056), .B1(n_1071), .B2(n_1072), .C(n_1073), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1055 ( .A(n_1056), .Y(n_1055) );
OAI21xp5_ASAP7_75t_L g1215 ( .A1(n_1057), .A2(n_1066), .B(n_1216), .Y(n_1215) );
INVx2_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1212 ( .A(n_1060), .Y(n_1212) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1060), .Y(n_1539) );
NAND2x2_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1063), .Y(n_1060) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1061), .Y(n_1067) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_SL g1210 ( .A(n_1065), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1543 ( .A(n_1066), .Y(n_1543) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1073), .B(n_1207), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1530 ( .A(n_1073), .Y(n_1530) );
AOI222xp33_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1079), .B1(n_1080), .B2(n_1083), .C1(n_1084), .C2(n_1086), .Y(n_1075) );
AOI21xp33_ASAP7_75t_SL g1541 ( .A1(n_1076), .A2(n_1542), .B(n_1543), .Y(n_1541) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1080), .Y(n_1224) );
AOI222xp33_ASAP7_75t_L g1537 ( .A1(n_1080), .A2(n_1507), .B1(n_1518), .B2(n_1538), .C1(n_1539), .C2(n_1540), .Y(n_1537) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
AOI211xp5_ASAP7_75t_L g1106 ( .A1(n_1083), .A2(n_1107), .B(n_1110), .C(n_1118), .Y(n_1106) );
AOI222xp33_ASAP7_75t_L g1524 ( .A1(n_1084), .A2(n_1508), .B1(n_1525), .B2(n_1530), .C1(n_1531), .C2(n_1534), .Y(n_1524) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1094), .B1(n_1095), .B2(n_1099), .C(n_1100), .Y(n_1091) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_1097), .A2(n_1116), .B1(n_1187), .B2(n_1188), .C(n_1189), .Y(n_1186) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
AOI22xp5_ASAP7_75t_L g1517 ( .A1(n_1102), .A2(n_1105), .B1(n_1499), .B2(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx4_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_1112), .A2(n_1114), .B1(n_1507), .B2(n_1508), .Y(n_1506) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_1115), .A2(n_1182), .B1(n_1186), .B2(n_1190), .C(n_1193), .Y(n_1181) );
OR2x6_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1121), .Y(n_1202) );
INVx3_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1126), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1126), .B(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
AND4x1_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1137), .C(n_1155), .D(n_1168), .Y(n_1133) );
OAI22xp5_ASAP7_75t_SL g1138 ( .A1(n_1139), .A2(n_1140), .B1(n_1147), .B2(n_1148), .Y(n_1138) );
OAI221xp5_ASAP7_75t_L g1251 ( .A1(n_1142), .A2(n_1252), .B1(n_1253), .B2(n_1254), .C(n_1255), .Y(n_1251) );
INVx3_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_1149), .A2(n_1150), .B1(n_1151), .B2(n_1152), .C(n_1153), .Y(n_1148) );
OAI211xp5_ASAP7_75t_L g1164 ( .A1(n_1150), .A2(n_1165), .B(n_1166), .C(n_1167), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g1257 ( .A1(n_1151), .A2(n_1244), .B1(n_1252), .B2(n_1258), .C(n_1259), .Y(n_1257) );
OAI22xp33_ASAP7_75t_SL g1169 ( .A1(n_1170), .A2(n_1171), .B1(n_1229), .B2(n_1265), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
XNOR2xp5_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
NOR2x1_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1203), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1179), .Y(n_1175) );
OAI211xp5_ASAP7_75t_L g1216 ( .A1(n_1187), .A2(n_1217), .B(n_1219), .C(n_1220), .Y(n_1216) );
OAI21xp5_ASAP7_75t_SL g1193 ( .A1(n_1194), .A2(n_1195), .B(n_1196), .Y(n_1193) );
OAI211xp5_ASAP7_75t_L g1519 ( .A1(n_1194), .A2(n_1520), .B(n_1521), .C(n_1522), .Y(n_1519) );
AOI22xp5_ASAP7_75t_L g1209 ( .A1(n_1199), .A2(n_1210), .B1(n_1211), .B2(n_1212), .Y(n_1209) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
NAND3xp33_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1221), .C(n_1225), .Y(n_1203) );
NOR3xp33_ASAP7_75t_SL g1204 ( .A(n_1205), .B(n_1213), .C(n_1215), .Y(n_1204) );
OAI21xp5_ASAP7_75t_SL g1205 ( .A1(n_1206), .A2(n_1208), .B(n_1209), .Y(n_1205) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1229), .Y(n_1265) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
AND4x1_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1249), .C(n_1261), .D(n_1264), .Y(n_1231) );
OAI21xp5_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1242), .B(n_1248), .Y(n_1232) );
INVx2_ASAP7_75t_SL g1236 ( .A(n_1237), .Y(n_1236) );
BUFx4f_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx3_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1277), .Y(n_1270) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1271), .B(n_1280), .Y(n_1549) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1275), .Y(n_1272) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_1273), .B(n_1276), .Y(n_1555) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1273), .Y(n_1563) );
HB1xp67_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1565 ( .A(n_1276), .B(n_1563), .Y(n_1565) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1281), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
AND2x4_ASAP7_75t_SL g1548 ( .A(n_1281), .B(n_1549), .Y(n_1548) );
INVx3_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
OAI221xp5_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1492), .B1(n_1495), .B2(n_1544), .C(n_1550), .Y(n_1284) );
AND4x1_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1447), .C(n_1465), .D(n_1481), .Y(n_1285) );
OAI33xp33_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1379), .A3(n_1397), .B1(n_1403), .B2(n_1415), .B3(n_1426), .Y(n_1286) );
OAI211xp5_ASAP7_75t_SL g1287 ( .A1(n_1288), .A2(n_1307), .B(n_1328), .C(n_1360), .Y(n_1287) );
INVx2_ASAP7_75t_L g1381 ( .A(n_1288), .Y(n_1381) );
AOI331xp33_ASAP7_75t_L g1404 ( .A1(n_1288), .A2(n_1309), .A3(n_1374), .B1(n_1402), .B2(n_1405), .B3(n_1407), .C1(n_1408), .Y(n_1404) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1288), .B(n_1330), .Y(n_1439) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1288), .B(n_1310), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1303), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1289), .B(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1289), .Y(n_1352) );
INVx2_ASAP7_75t_SL g1373 ( .A(n_1289), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1289), .B(n_1310), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1289), .B(n_1485), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1297), .Y(n_1289) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1291), .Y(n_1494) );
AND2x6_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1293), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1292), .B(n_1296), .Y(n_1295) );
AND2x4_ASAP7_75t_L g1298 ( .A(n_1292), .B(n_1299), .Y(n_1298) );
AND2x6_ASAP7_75t_L g1301 ( .A(n_1292), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1292), .B(n_1296), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1292), .B(n_1296), .Y(n_1377) );
OAI21xp5_ASAP7_75t_L g1562 ( .A1(n_1293), .A2(n_1563), .B(n_1564), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1294), .B(n_1300), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g1345 ( .A(n_1303), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1303), .B(n_1352), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1303), .B(n_1311), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1303), .B(n_1410), .Y(n_1409) );
AOI22xp5_ASAP7_75t_L g1416 ( .A1(n_1303), .A2(n_1395), .B1(n_1417), .B2(n_1420), .Y(n_1416) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_1303), .A2(n_1389), .B1(n_1457), .B2(n_1463), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1303), .B(n_1340), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1303), .B(n_1341), .Y(n_1491) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1306), .Y(n_1303) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1314), .Y(n_1308) );
O2A1O1Ixp33_ASAP7_75t_SL g1353 ( .A1(n_1309), .A2(n_1354), .B(n_1355), .C(n_1357), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1309), .B(n_1468), .Y(n_1467) );
CKINVDCx14_ASAP7_75t_R g1309 ( .A(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1310), .B(n_1315), .Y(n_1386) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1310), .B(n_1389), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1310), .B(n_1349), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1310), .B(n_1381), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1310), .B(n_1419), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1310), .B(n_1314), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1310), .B(n_1373), .Y(n_1453) );
INVx3_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_1311), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1311), .B(n_1356), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1311), .B(n_1384), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1311), .B(n_1316), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1311), .B(n_1389), .Y(n_1413) );
AND2x4_ASAP7_75t_SL g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1319), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1315), .B(n_1325), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1315), .B(n_1348), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1315), .B(n_1368), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1315), .B(n_1362), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1315), .B(n_1349), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1315), .B(n_1320), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1315), .B(n_1331), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1315), .B(n_1393), .Y(n_1475) );
INVx2_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1316), .B(n_1331), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1316), .B(n_1325), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1316), .B(n_1362), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1316), .B(n_1332), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1384 ( .A(n_1316), .B(n_1321), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1316), .B(n_1402), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1316), .B(n_1363), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1316), .B(n_1321), .Y(n_1462) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_1316), .B(n_1478), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1318), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1319), .B(n_1356), .Y(n_1478) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1324), .Y(n_1320) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1321), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1321), .B(n_1325), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1325), .B(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1325), .Y(n_1363) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1325), .Y(n_1368) );
NAND2x1_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1327), .Y(n_1325) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_1329), .A2(n_1337), .B1(n_1346), .B2(n_1350), .C(n_1353), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1333), .Y(n_1329) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1330), .Y(n_1468) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1331), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1332), .B(n_1363), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1335), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1334), .B(n_1336), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1334), .B(n_1362), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1334), .B(n_1371), .Y(n_1420) );
OR2x2_ASAP7_75t_L g1432 ( .A(n_1334), .B(n_1351), .Y(n_1432) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1334), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1334), .B(n_1412), .Y(n_1472) );
AOI22xp5_ASAP7_75t_L g1423 ( .A1(n_1335), .A2(n_1345), .B1(n_1390), .B2(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1337), .B(n_1346), .Y(n_1414) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1344), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1340), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1340), .B(n_1358), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1340), .B(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1341), .Y(n_1374) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1341), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1341), .B(n_1345), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1341), .B(n_1438), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1341), .B(n_1453), .Y(n_1452) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1345), .B(n_1373), .Y(n_1372) );
OAI32xp33_ASAP7_75t_L g1385 ( .A1(n_1345), .A2(n_1354), .A3(n_1362), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
HB1xp67_ASAP7_75t_SL g1398 ( .A(n_1345), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1345), .B(n_1392), .Y(n_1458) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1486 ( .A(n_1348), .B(n_1386), .Y(n_1486) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1349), .B(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1351), .Y(n_1480) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1352), .Y(n_1358) );
AOI31xp33_ASAP7_75t_L g1469 ( .A1(n_1352), .A2(n_1429), .A3(n_1470), .B(n_1471), .Y(n_1469) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1354), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1354), .B(n_1406), .Y(n_1405) );
OAI221xp5_ASAP7_75t_L g1415 ( .A1(n_1357), .A2(n_1374), .B1(n_1416), .B2(n_1421), .C(n_1423), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1359), .Y(n_1357) );
OAI221xp5_ASAP7_75t_SL g1379 ( .A1(n_1358), .A2(n_1380), .B1(n_1392), .B2(n_1393), .C(n_1394), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1358), .B(n_1390), .Y(n_1464) );
AOI221xp5_ASAP7_75t_L g1360 ( .A1(n_1361), .A2(n_1364), .B1(n_1365), .B2(n_1374), .C(n_1375), .Y(n_1360) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1361), .Y(n_1488) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1362), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1362), .B(n_1391), .Y(n_1460) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1369), .B1(n_1370), .B2(n_1372), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVxp33_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1372), .Y(n_1419) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1373), .Y(n_1389) );
O2A1O1Ixp33_ASAP7_75t_L g1397 ( .A1(n_1373), .A2(n_1398), .B(n_1399), .C(n_1400), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1373), .B(n_1390), .Y(n_1449) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1374), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1481 ( .A1(n_1374), .A2(n_1468), .B1(n_1482), .B2(n_1483), .C(n_1487), .Y(n_1481) );
INVx3_ASAP7_75t_L g1440 ( .A(n_1375), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1378), .Y(n_1375) );
AOI211xp5_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1382), .B(n_1385), .C(n_1390), .Y(n_1380) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1389), .B(n_1407), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1396), .Y(n_1394) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1396), .Y(n_1451) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1414), .Y(n_1403) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1407), .Y(n_1443) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_1407), .A2(n_1458), .B1(n_1459), .B2(n_1461), .Y(n_1457) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVxp33_ASAP7_75t_SL g1489 ( .A(n_1410), .Y(n_1489) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1413), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1420), .Y(n_1470) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
NAND3xp33_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1433), .C(n_1441), .Y(n_1426) );
INVxp67_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
AOI21xp33_ASAP7_75t_L g1428 ( .A1(n_1429), .A2(n_1431), .B(n_1432), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
NOR2xp33_ASAP7_75t_L g1454 ( .A(n_1430), .B(n_1455), .Y(n_1454) );
AOI211xp5_ASAP7_75t_L g1433 ( .A1(n_1434), .A2(n_1436), .B(n_1439), .C(n_1440), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
NOR2xp33_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1444), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1446), .Y(n_1444) );
INVx2_ASAP7_75t_L g1455 ( .A(n_1446), .Y(n_1455) );
AOI211xp5_ASAP7_75t_L g1447 ( .A1(n_1448), .A2(n_1449), .B(n_1450), .C(n_1456), .Y(n_1447) );
AOI21xp33_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1452), .B(n_1454), .Y(n_1450) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVxp33_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
O2A1O1Ixp33_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1469), .B(n_1473), .C(n_1474), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
AOI21xp5_ASAP7_75t_L g1474 ( .A1(n_1475), .A2(n_1476), .B(n_1479), .Y(n_1474) );
INVxp33_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVxp67_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
AOI21xp33_ASAP7_75t_L g1487 ( .A1(n_1488), .A2(n_1489), .B(n_1490), .Y(n_1487) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
CKINVDCx20_ASAP7_75t_R g1492 ( .A(n_1493), .Y(n_1492) );
CKINVDCx20_ASAP7_75t_R g1493 ( .A(n_1494), .Y(n_1493) );
HB1xp67_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVxp33_ASAP7_75t_L g1559 ( .A(n_1497), .Y(n_1559) );
AOI211x1_ASAP7_75t_L g1497 ( .A1(n_1498), .A2(n_1499), .B(n_1500), .C(n_1523), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1503), .Y(n_1500) );
NAND3xp33_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1517), .C(n_1519), .Y(n_1509) );
INVx3_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
NAND3xp33_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1537), .C(n_1541), .Y(n_1523) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
CKINVDCx20_ASAP7_75t_R g1544 ( .A(n_1545), .Y(n_1544) );
CKINVDCx20_ASAP7_75t_R g1545 ( .A(n_1546), .Y(n_1545) );
INVx3_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
BUFx3_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
HB1xp67_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
BUFx3_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVxp67_ASAP7_75t_SL g1556 ( .A(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
HB1xp67_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
endmodule