module real_jpeg_10360_n_16 (n_301, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_301;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_243;
wire n_173;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_293;
wire n_164;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx24_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_73),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_40),
.B1(n_49),
.B2(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_57),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_57),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_4),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_27),
.B1(n_33),
.B2(n_161),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_4),
.B(n_51),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_42),
.B(n_46),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_4),
.A2(n_40),
.B1(n_49),
.B2(n_159),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_57),
.B(n_60),
.C(n_61),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_7),
.B(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_36),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_10),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_10),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_40),
.B1(n_49),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_13),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_150),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_150),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_13),
.A2(n_40),
.B1(n_49),
.B2(n_150),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_14),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_141),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_141),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_14),
.A2(n_40),
.B1(n_49),
.B2(n_141),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_15),
.A2(n_40),
.B1(n_49),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_15),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_99),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_99),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_99),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_20),
.B(n_107),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_21),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_21),
.B(n_292),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_69),
.CI(n_88),
.CON(n_21),
.SN(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_54),
.B2(n_68),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_25),
.A2(n_38),
.B(n_68),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_25),
.A2(n_26),
.B1(n_55),
.B2(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_27),
.A2(n_33),
.B1(n_140),
.B2(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_27),
.A2(n_93),
.B(n_143),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_27),
.A2(n_34),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_27),
.A2(n_33),
.B1(n_206),
.B2(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_27),
.A2(n_192),
.B(n_228),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_28),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_28),
.A2(n_32),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_29),
.B(n_62),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_29),
.B(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_30),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_32),
.B(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_32),
.B(n_92),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_33),
.B(n_159),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_33),
.A2(n_91),
.B(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_47),
.B(n_50),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_39),
.A2(n_98),
.B(n_100),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_39),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_39),
.A2(n_44),
.B1(n_242),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_39),
.A2(n_44),
.B1(n_98),
.B2(n_251),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_40),
.A2(n_41),
.B(n_159),
.C(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_44),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_75),
.B(n_77),
.C(n_78),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_75),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g184 ( 
.A(n_46),
.B(n_159),
.CON(n_184),
.SN(n_184)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_48),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_51),
.A2(n_115),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_55),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_65),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_61),
.B1(n_63),
.B2(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_56),
.A2(n_61),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_56),
.A2(n_61),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_56),
.A2(n_61),
.B1(n_149),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_56),
.A2(n_61),
.B1(n_174),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_56),
.A2(n_81),
.B(n_182),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_58),
.B1(n_75),
.B2(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_57),
.B(n_75),
.Y(n_190)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_77),
.B1(n_184),
.B2(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_61),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_61),
.A2(n_84),
.B(n_95),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_66),
.A2(n_83),
.B(n_86),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_80),
.B(n_87),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_80),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_74),
.B(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_74),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_74),
.A2(n_78),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_74),
.A2(n_122),
.B(n_254),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_78),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_79),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_109),
.B1(n_110),
.B2(n_127),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.C(n_101),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_89),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_90),
.B(n_94),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_159),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_103),
.A2(n_119),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_103),
.A2(n_119),
.B1(n_202),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_128),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_119),
.A2(n_238),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_279),
.A3(n_291),
.B1(n_293),
.B2(n_299),
.C(n_301),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_244),
.C(n_275),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_218),
.B(n_243),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_195),
.B(n_217),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_177),
.B(n_194),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_168),
.B(n_176),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_156),
.B(n_167),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_144),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_151),
.B2(n_155),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_145),
.B(n_155),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_162),
.B(n_166),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_169),
.B(n_170),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_178),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.CI(n_175),
.CON(n_171),
.SN(n_171)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_188),
.B2(n_193),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_187),
.C(n_193),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_211),
.B2(n_212),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_214),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_203),
.B1(n_204),
.B2(n_210),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_208),
.C(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_232),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_231),
.C(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_236),
.C(n_239),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_262),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_262),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_256),
.C(n_260),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_249),
.C(n_255),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_255),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_252),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_271),
.C(n_272),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_267),
.C(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_280),
.A2(n_294),
.B(n_298),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_288),
.C(n_290),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B(n_297),
.Y(n_294)
);


endmodule