module fake_jpeg_16193_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_21),
.B1(n_20),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_58),
.B1(n_68),
.B2(n_21),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_21),
.B1(n_34),
.B2(n_25),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_25),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_98),
.B1(n_102),
.B2(n_19),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_49),
.B1(n_45),
.B2(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_106),
.B1(n_18),
.B2(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_45),
.B1(n_40),
.B2(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_92),
.B1(n_94),
.B2(n_105),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_31),
.B(n_17),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_82),
.C(n_88),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_97),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_92)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_32),
.A3(n_26),
.B1(n_33),
.B2(n_23),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_28),
.B(n_24),
.C(n_30),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_41),
.B1(n_37),
.B2(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_32),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_100),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_36),
.B1(n_33),
.B2(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_36),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_51),
.A2(n_29),
.B1(n_18),
.B2(n_24),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_23),
.B1(n_16),
.B2(n_14),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_47),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_110),
.B1(n_83),
.B2(n_103),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_66),
.B1(n_35),
.B2(n_19),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_127),
.B(n_88),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_135),
.Y(n_137)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_35),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_100),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_66),
.B1(n_55),
.B2(n_59),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_104),
.B1(n_97),
.B2(n_57),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_19),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_130),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_106),
.B1(n_77),
.B2(n_86),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_30),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_99),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_125),
.B1(n_99),
.B2(n_121),
.Y(n_153)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_30),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_144),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_150),
.B(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_76),
.C(n_81),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_119),
.C(n_109),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_146),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_113),
.B1(n_131),
.B2(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_101),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_149),
.B1(n_154),
.B2(n_155),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_91),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_101),
.B1(n_80),
.B2(n_94),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_107),
.B(n_84),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_52),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_156),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_104),
.B1(n_105),
.B2(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_57),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_57),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_111),
.A2(n_48),
.B(n_22),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_48),
.B(n_30),
.C(n_104),
.D(n_9),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_14),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_48),
.B(n_53),
.C(n_52),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_125),
.B1(n_112),
.B2(n_136),
.Y(n_185)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_0),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_123),
.B1(n_111),
.B2(n_124),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_53),
.B1(n_14),
.B2(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_161),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_173),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_115),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_177),
.C(n_180),
.Y(n_208)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_131),
.B1(n_113),
.B2(n_119),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_176),
.B1(n_185),
.B2(n_186),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_134),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_134),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_181),
.A2(n_160),
.B(n_169),
.Y(n_223)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_183),
.Y(n_233)
);

CKINVDCx12_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_109),
.C(n_125),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_164),
.C(n_159),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_135),
.B1(n_9),
.B2(n_10),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_30),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_196),
.B1(n_160),
.B2(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_203),
.Y(n_224)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_145),
.B1(n_149),
.B2(n_168),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_13),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_53),
.B1(n_11),
.B2(n_10),
.Y(n_203)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_138),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_216),
.C(n_229),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_142),
.CI(n_147),
.CON(n_209),
.SN(n_209)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_225),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_220),
.B(n_223),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_227),
.B(n_201),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_151),
.Y(n_218)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_228),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_178),
.A2(n_137),
.B(n_162),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_175),
.B(n_167),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_155),
.Y(n_229)
);

OAI22x1_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_162),
.B1(n_167),
.B2(n_3),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_192),
.B1(n_186),
.B2(n_162),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_162),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_170),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_239),
.C(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_237),
.B(n_254),
.Y(n_274)
);

AO22x1_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_181),
.B1(n_171),
.B2(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_180),
.C(n_184),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_248),
.B(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_193),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_251),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_198),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_188),
.C(n_190),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_256),
.C(n_222),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_215),
.B(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_173),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_219),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_196),
.C(n_204),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_212),
.B(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_222),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_182),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_266),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_261),
.A2(n_265),
.B(n_226),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_218),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_228),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_223),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_277),
.C(n_234),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_225),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_247),
.A2(n_224),
.B1(n_213),
.B2(n_217),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_278),
.B1(n_263),
.B2(n_280),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_247),
.A2(n_224),
.B1(n_213),
.B2(n_226),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_270),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_280),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_235),
.B1(n_256),
.B2(n_244),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_251),
.B1(n_246),
.B2(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_239),
.C(n_236),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_252),
.C(n_245),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_264),
.B(n_260),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_297),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_262),
.B(n_248),
.CI(n_238),
.CON(n_295),
.SN(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_241),
.C(n_221),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_233),
.C(n_211),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_311),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_295),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_261),
.B1(n_267),
.B2(n_266),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_309),
.B1(n_291),
.B2(n_242),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_297),
.C(n_281),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_2),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_273),
.B1(n_265),
.B2(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_279),
.B1(n_267),
.B2(n_278),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_295),
.B1(n_286),
.B2(n_296),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_285),
.A2(n_276),
.B(n_238),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_211),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_270),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_323),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_321),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_275),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_319),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_324),
.C(n_300),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_292),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_305),
.A3(n_309),
.B1(n_308),
.B2(n_304),
.C1(n_310),
.C2(n_303),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_1),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_332),
.C(n_4),
.Y(n_334)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_327),
.Y(n_339)
);

NAND4xp25_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_315),
.C(n_318),
.D(n_320),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_316),
.B1(n_3),
.B2(n_4),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_7),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_2),
.C(n_3),
.Y(n_332)
);

AOI31xp33_ASAP7_75t_L g333 ( 
.A1(n_314),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_336),
.C(n_332),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_335),
.B(n_337),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_6),
.C(n_7),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_330),
.B(n_329),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_326),
.B1(n_342),
.B2(n_339),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_329),
.C(n_331),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_340),
.B(n_337),
.Y(n_346)
);


endmodule