module fake_jpeg_11473_n_182 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_17),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_62),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_39),
.B1(n_49),
.B2(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_37),
.B(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_15),
.C(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_33),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_29),
.B1(n_28),
.B2(n_18),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_90),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_99),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_96),
.B1(n_68),
.B2(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_41),
.B1(n_36),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_46),
.B1(n_43),
.B2(n_41),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_78),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_36),
.B1(n_45),
.B2(n_32),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_35),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_12),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_87),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_73),
.C(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_109),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_83),
.B1(n_81),
.B2(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_110),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_74),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_75),
.B1(n_65),
.B2(n_60),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_121),
.B(n_95),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_134),
.B(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_94),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_97),
.B(n_59),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_120),
.B(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_117),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_150),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_103),
.C(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_135),
.C(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_114),
.B1(n_108),
.B2(n_84),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_122),
.B1(n_131),
.B2(n_126),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_154),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_144),
.C(n_142),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_129),
.B1(n_120),
.B2(n_128),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_60),
.C(n_82),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_149),
.C(n_147),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_140),
.B(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_151),
.B1(n_145),
.B2(n_141),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_145),
.C(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_153),
.C(n_151),
.Y(n_169)
);

NOR4xp25_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.D(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_164),
.A3(n_165),
.B1(n_141),
.B2(n_159),
.C1(n_13),
.C2(n_14),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_174),
.B(n_9),
.Y(n_177)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_173),
.C(n_11),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_12),
.B(n_5),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_180),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_181),
.Y(n_182)
);


endmodule