module real_aes_9729_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_2043;
wire n_476;
wire n_887;
wire n_599;
wire n_2003;
wire n_2014;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_2006;
wire n_963;
wire n_551;
wire n_884;
wire n_2035;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_2031;
wire n_1160;
wire n_1849;
wire n_2040;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1994;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1959;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_1301;
wire n_728;
wire n_2004;
wire n_1201;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_2038;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_2041;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1648;
wire n_724;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_2012;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2045;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_2036;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_2033;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_402;
wire n_733;
wire n_602;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2039;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_2023;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_2019;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_2042;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1638;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_2032;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_2034;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_719;
wire n_465;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1931;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_2037;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_2030;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_2044;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_2010;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g1214 ( .A(n_0), .B(n_1215), .Y(n_1214) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_1), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_2), .A2(n_339), .B1(n_473), .B2(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g575 ( .A(n_2), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g1685 ( .A1(n_3), .A2(n_364), .B1(n_1686), .B2(n_1694), .Y(n_1685) );
CKINVDCx5p33_ASAP7_75t_R g757 ( .A(n_4), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_5), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g1635 ( .A1(n_6), .A2(n_264), .B1(n_545), .B2(n_1636), .C(n_1638), .Y(n_1635) );
INVx1_ASAP7_75t_L g1653 ( .A(n_6), .Y(n_1653) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_7), .A2(n_111), .B1(n_998), .B2(n_1000), .Y(n_997) );
INVx1_ASAP7_75t_L g1042 ( .A(n_7), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1593 ( .A1(n_8), .A2(n_334), .B1(n_411), .B2(n_422), .Y(n_1593) );
INVx1_ASAP7_75t_L g1612 ( .A(n_8), .Y(n_1612) );
INVx1_ASAP7_75t_L g618 ( .A(n_9), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_9), .A2(n_155), .B1(n_685), .B2(n_688), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_10), .Y(n_445) );
INVx1_ASAP7_75t_L g882 ( .A(n_11), .Y(n_882) );
INVx1_ASAP7_75t_L g1110 ( .A(n_12), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_12), .A2(n_120), .B1(n_479), .B2(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1234 ( .A(n_13), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_13), .A2(n_207), .B1(n_928), .B2(n_929), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1505 ( .A1(n_14), .A2(n_35), .B1(n_795), .B2(n_1506), .C(n_1507), .Y(n_1505) );
INVx1_ASAP7_75t_L g1533 ( .A(n_14), .Y(n_1533) );
OAI22xp33_ASAP7_75t_L g1075 ( .A1(n_15), .A2(n_109), .B1(n_517), .B2(n_558), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_15), .A2(n_109), .B1(n_485), .B2(n_1078), .C(n_1084), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_16), .A2(n_128), .B1(n_1124), .B2(n_1126), .Y(n_1123) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_16), .A2(n_128), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
INVx1_ASAP7_75t_L g912 ( .A(n_17), .Y(n_912) );
OAI211xp5_ASAP7_75t_SL g938 ( .A1(n_17), .A2(n_517), .B(n_939), .C(n_948), .Y(n_938) );
AOI221xp5_ASAP7_75t_L g1415 ( .A1(n_18), .A2(n_314), .B1(n_612), .B2(n_613), .C(n_947), .Y(n_1415) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_18), .A2(n_314), .B1(n_479), .B2(n_1422), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_19), .Y(n_906) );
INVx1_ASAP7_75t_L g1588 ( .A(n_20), .Y(n_1588) );
CKINVDCx20_ASAP7_75t_R g1462 ( .A(n_21), .Y(n_1462) );
AOI22xp5_ASAP7_75t_L g1697 ( .A1(n_22), .A2(n_321), .B1(n_1698), .B2(n_1702), .Y(n_1697) );
CKINVDCx16_ASAP7_75t_R g1628 ( .A(n_23), .Y(n_1628) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_24), .A2(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g645 ( .A(n_24), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g1440 ( .A(n_25), .B(n_1441), .Y(n_1440) );
CKINVDCx16_ASAP7_75t_R g1735 ( .A(n_25), .Y(n_1735) );
INVx1_ASAP7_75t_L g1948 ( .A(n_26), .Y(n_1948) );
AOI22xp33_ASAP7_75t_L g1977 ( .A1(n_26), .A2(n_133), .B1(n_799), .B2(n_1199), .Y(n_1977) );
AOI22xp33_ASAP7_75t_SL g1127 ( .A1(n_27), .A2(n_103), .B1(n_1124), .B2(n_1128), .Y(n_1127) );
INVxp67_ASAP7_75t_SL g1157 ( .A(n_27), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1499 ( .A1(n_28), .A2(n_144), .B1(n_1500), .B2(n_1501), .Y(n_1499) );
INVx1_ASAP7_75t_L g1519 ( .A(n_28), .Y(n_1519) );
XNOR2xp5_ASAP7_75t_L g1930 ( .A(n_29), .B(n_1931), .Y(n_1930) );
OAI222xp33_ASAP7_75t_L g1312 ( .A1(n_30), .A2(n_76), .B1(n_159), .B2(n_1148), .C1(n_1151), .C2(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1327 ( .A(n_30), .Y(n_1327) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_31), .Y(n_1385) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_32), .Y(n_1502) );
CKINVDCx5p33_ASAP7_75t_R g1999 ( .A(n_33), .Y(n_1999) );
INVx1_ASAP7_75t_L g1643 ( .A(n_34), .Y(n_1643) );
AOI22xp33_ASAP7_75t_SL g1674 ( .A1(n_34), .A2(n_322), .B1(n_694), .B2(n_780), .Y(n_1674) );
INVx1_ASAP7_75t_L g1531 ( .A(n_35), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_36), .A2(n_79), .B1(n_627), .B2(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1656 ( .A(n_36), .Y(n_1656) );
AOI221xp5_ASAP7_75t_L g1403 ( .A1(n_37), .A2(n_215), .B1(n_545), .B2(n_1404), .C(n_1405), .Y(n_1403) );
INVx1_ASAP7_75t_L g1429 ( .A(n_37), .Y(n_1429) );
INVx1_ASAP7_75t_L g713 ( .A(n_38), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_38), .A2(n_169), .B1(n_774), .B2(n_775), .C(n_777), .Y(n_773) );
INVx1_ASAP7_75t_L g1639 ( .A(n_39), .Y(n_1639) );
AOI22xp33_ASAP7_75t_L g1673 ( .A1(n_39), .A2(n_178), .B1(n_688), .B2(n_1669), .Y(n_1673) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_40), .B(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1040 ( .A(n_40), .Y(n_1040) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_41), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_42), .A2(n_164), .B1(n_491), .B2(n_1358), .Y(n_1357) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_42), .A2(n_164), .B1(n_630), .B2(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g381 ( .A(n_43), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_44), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g1640 ( .A1(n_45), .A2(n_127), .B1(n_555), .B2(n_1408), .Y(n_1640) );
INVx1_ASAP7_75t_L g1664 ( .A(n_45), .Y(n_1664) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_46), .A2(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g680 ( .A(n_46), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g2020 ( .A(n_47), .Y(n_2020) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_48), .A2(n_168), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
INVx1_ASAP7_75t_L g1430 ( .A(n_48), .Y(n_1430) );
AOI22xp5_ASAP7_75t_L g1721 ( .A1(n_49), .A2(n_167), .B1(n_1686), .B2(n_1694), .Y(n_1721) );
XOR2xp5_ASAP7_75t_L g1584 ( .A(n_50), .B(n_1585), .Y(n_1584) );
AOI22xp33_ASAP7_75t_L g1754 ( .A1(n_50), .A2(n_241), .B1(n_1723), .B2(n_1755), .Y(n_1754) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_51), .Y(n_1113) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_51), .A2(n_190), .B1(n_1148), .B2(n_1151), .Y(n_1147) );
INVx1_ASAP7_75t_L g1164 ( .A(n_52), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_52), .A2(n_232), .B1(n_1121), .B2(n_1191), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_53), .A2(n_161), .B1(n_542), .B2(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_53), .A2(n_161), .B1(n_1078), .B2(n_1138), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_54), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_55), .A2(n_265), .B1(n_479), .B2(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g566 ( .A(n_55), .Y(n_566) );
INVx1_ASAP7_75t_L g739 ( .A(n_56), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_56), .A2(n_142), .B1(n_799), .B2(n_800), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g1957 ( .A(n_57), .Y(n_1957) );
AOI22xp5_ASAP7_75t_L g1705 ( .A1(n_58), .A2(n_145), .B1(n_1686), .B2(n_1694), .Y(n_1705) );
AO221x2_ASAP7_75t_L g1711 ( .A1(n_59), .A2(n_279), .B1(n_1698), .B2(n_1702), .C(n_1712), .Y(n_1711) );
CKINVDCx16_ASAP7_75t_R g1737 ( .A(n_60), .Y(n_1737) );
INVx1_ASAP7_75t_L g851 ( .A(n_61), .Y(n_851) );
INVx1_ASAP7_75t_L g1492 ( .A(n_62), .Y(n_1492) );
XNOR2xp5_ASAP7_75t_L g889 ( .A(n_63), .B(n_890), .Y(n_889) );
AOI22xp5_ASAP7_75t_SL g1741 ( .A1(n_63), .A2(n_258), .B1(n_1702), .B2(n_1723), .Y(n_1741) );
INVx1_ASAP7_75t_L g1552 ( .A(n_64), .Y(n_1552) );
OAI221xp5_ASAP7_75t_L g1565 ( .A1(n_64), .A2(n_517), .B1(n_1566), .B2(n_1570), .C(n_1574), .Y(n_1565) );
INVx1_ASAP7_75t_L g1604 ( .A(n_65), .Y(n_1604) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_65), .A2(n_250), .B1(n_1360), .B2(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1284 ( .A(n_66), .Y(n_1284) );
INVx1_ASAP7_75t_L g1481 ( .A(n_67), .Y(n_1481) );
OAI22xp33_ASAP7_75t_L g1487 ( .A1(n_67), .A2(n_143), .B1(n_422), .B2(n_1262), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1647 ( .A1(n_68), .A2(n_256), .B1(n_1648), .B2(n_1649), .Y(n_1647) );
AOI22xp33_ASAP7_75t_L g1667 ( .A1(n_68), .A2(n_256), .B1(n_1199), .B2(n_1506), .Y(n_1667) );
INVx1_ASAP7_75t_L g1330 ( .A(n_69), .Y(n_1330) );
AOI22xp33_ASAP7_75t_SL g1346 ( .A1(n_69), .A2(n_126), .B1(n_1078), .B2(n_1207), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_70), .A2(n_375), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
INVx1_ASAP7_75t_L g1470 ( .A(n_70), .Y(n_1470) );
CKINVDCx14_ASAP7_75t_R g1793 ( .A(n_71), .Y(n_1793) );
INVx1_ASAP7_75t_L g1599 ( .A(n_72), .Y(n_1599) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_72), .A2(n_210), .B1(n_874), .B2(n_1451), .Y(n_1619) );
INVx1_ASAP7_75t_L g1057 ( .A(n_73), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_73), .A2(n_272), .B1(n_1078), .B2(n_1080), .C(n_1082), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_74), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g1396 ( .A(n_75), .B(n_1397), .Y(n_1396) );
AOI22xp33_ASAP7_75t_SL g1334 ( .A1(n_76), .A2(n_326), .B1(n_542), .B2(n_1335), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_77), .A2(n_209), .B1(n_1124), .B2(n_1189), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_77), .A2(n_209), .B1(n_1135), .B2(n_1199), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g1546 ( .A(n_78), .Y(n_1546) );
INVx1_ASAP7_75t_L g1654 ( .A(n_79), .Y(n_1654) );
INVxp33_ASAP7_75t_SL g827 ( .A(n_80), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_80), .A2(n_365), .B1(n_867), .B2(n_869), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1752 ( .A1(n_81), .A2(n_222), .B1(n_1686), .B2(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1595 ( .A(n_82), .Y(n_1595) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_83), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g1511 ( .A(n_84), .Y(n_1511) );
OAI22xp33_ASAP7_75t_L g920 ( .A1(n_85), .A2(n_366), .B1(n_921), .B2(n_923), .Y(n_920) );
INVx1_ASAP7_75t_L g950 ( .A(n_85), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_86), .Y(n_1274) );
OAI22xp5_ASAP7_75t_L g1503 ( .A1(n_87), .A2(n_268), .B1(n_784), .B2(n_787), .Y(n_1503) );
OAI221xp5_ASAP7_75t_L g1524 ( .A1(n_87), .A2(n_268), .B1(n_724), .B2(n_731), .C(n_734), .Y(n_1524) );
INVx1_ASAP7_75t_L g1567 ( .A(n_88), .Y(n_1567) );
OAI22xp33_ASAP7_75t_L g1578 ( .A1(n_88), .A2(n_182), .B1(n_411), .B2(n_422), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_89), .A2(n_369), .B1(n_480), .B2(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_89), .A2(n_558), .B1(n_560), .B2(n_574), .C(n_580), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g1962 ( .A(n_90), .Y(n_1962) );
INVx1_ASAP7_75t_L g1165 ( .A(n_91), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_91), .A2(n_180), .B1(n_1124), .B2(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g709 ( .A(n_92), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_92), .A2(n_240), .B1(n_780), .B2(n_781), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_93), .Y(n_1226) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_94), .Y(n_1447) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_95), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_95), .A2(n_371), .B1(n_874), .B2(n_876), .C(n_877), .Y(n_873) );
INVx1_ASAP7_75t_L g1277 ( .A(n_96), .Y(n_1277) );
OAI221xp5_ASAP7_75t_L g1287 ( .A1(n_96), .A2(n_558), .B1(n_638), .B2(n_1288), .C(n_1289), .Y(n_1287) );
INVx1_ASAP7_75t_L g918 ( .A(n_97), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_97), .A2(n_315), .B1(n_928), .B2(n_929), .Y(n_927) );
CKINVDCx14_ASAP7_75t_R g1713 ( .A(n_98), .Y(n_1713) );
XNOR2x2_ASAP7_75t_L g1048 ( .A(n_99), .B(n_1049), .Y(n_1048) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_100), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_100), .A2(n_277), .B1(n_800), .B2(n_1135), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_101), .A2(n_132), .B1(n_724), .B2(n_731), .C(n_734), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_101), .A2(n_132), .B1(n_784), .B2(n_787), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_102), .Y(n_1068) );
INVxp33_ASAP7_75t_L g1156 ( .A(n_103), .Y(n_1156) );
INVx1_ASAP7_75t_L g419 ( .A(n_104), .Y(n_419) );
BUFx2_ASAP7_75t_L g471 ( .A(n_104), .Y(n_471) );
BUFx2_ASAP7_75t_L g493 ( .A(n_104), .Y(n_493) );
OR2x2_ASAP7_75t_L g730 ( .A(n_104), .B(n_511), .Y(n_730) );
INVx1_ASAP7_75t_L g602 ( .A(n_105), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_105), .A2(n_146), .B1(n_490), .B2(n_694), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g2016 ( .A1(n_106), .A2(n_330), .B1(n_613), .B2(n_719), .C(n_2017), .Y(n_2016) );
INVx1_ASAP7_75t_L g2028 ( .A(n_106), .Y(n_2028) );
OAI22xp33_ASAP7_75t_L g1282 ( .A1(n_107), .A2(n_115), .B1(n_447), .B2(n_460), .Y(n_1282) );
INVx1_ASAP7_75t_L g1301 ( .A(n_107), .Y(n_1301) );
CKINVDCx5p33_ASAP7_75t_R g1960 ( .A(n_108), .Y(n_1960) );
CKINVDCx5p33_ASAP7_75t_R g1937 ( .A(n_110), .Y(n_1937) );
INVx1_ASAP7_75t_L g986 ( .A(n_111), .Y(n_986) );
INVx1_ASAP7_75t_L g1571 ( .A(n_112), .Y(n_1571) );
OAI22xp33_ASAP7_75t_L g1579 ( .A1(n_112), .A2(n_211), .B1(n_954), .B2(n_957), .Y(n_1579) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_113), .Y(n_1055) );
INVx1_ASAP7_75t_L g429 ( .A(n_114), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_114), .A2(n_310), .B1(n_540), .B2(n_542), .C(n_545), .Y(n_539) );
INVx1_ASAP7_75t_L g1300 ( .A(n_115), .Y(n_1300) );
INVx1_ASAP7_75t_L g1555 ( .A(n_116), .Y(n_1555) );
OAI22xp5_ASAP7_75t_L g1560 ( .A1(n_116), .A2(n_121), .B1(n_928), .B2(n_929), .Y(n_1560) );
OAI221xp5_ASAP7_75t_L g828 ( .A1(n_117), .A2(n_198), .B1(n_724), .B2(n_734), .C(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_117), .A2(n_198), .B1(n_784), .B2(n_871), .Y(n_870) );
AOI221xp5_ASAP7_75t_L g1645 ( .A1(n_118), .A2(n_200), .B1(n_613), .B2(n_1111), .C(n_1646), .Y(n_1645) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_118), .A2(n_200), .B1(n_1669), .B2(n_1672), .Y(n_1668) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_119), .A2(n_219), .B1(n_1121), .B2(n_1130), .Y(n_1129) );
INVxp67_ASAP7_75t_SL g1146 ( .A(n_119), .Y(n_1146) );
INVxp33_ASAP7_75t_L g1105 ( .A(n_120), .Y(n_1105) );
INVx1_ASAP7_75t_L g1554 ( .A(n_121), .Y(n_1554) );
AO221x1_ASAP7_75t_L g1380 ( .A1(n_122), .A2(n_214), .B1(n_635), .B2(n_636), .C(n_1131), .Y(n_1380) );
INVx1_ASAP7_75t_L g1389 ( .A(n_122), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_123), .A2(n_292), .B1(n_799), .B2(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1534 ( .A(n_123), .Y(n_1534) );
INVx1_ASAP7_75t_L g1324 ( .A(n_124), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_124), .A2(n_237), .B1(n_491), .B2(n_1135), .Y(n_1347) );
OAI221xp5_ASAP7_75t_L g1597 ( .A1(n_125), .A2(n_558), .B1(n_638), .B2(n_1598), .C(n_1602), .Y(n_1597) );
AOI22xp33_ASAP7_75t_SL g1620 ( .A1(n_125), .A2(n_284), .B1(n_799), .B2(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1326 ( .A(n_126), .Y(n_1326) );
INVx1_ASAP7_75t_L g1663 ( .A(n_127), .Y(n_1663) );
CKINVDCx5p33_ASAP7_75t_R g2021 ( .A(n_129), .Y(n_2021) );
INVx1_ASAP7_75t_L g1281 ( .A(n_130), .Y(n_1281) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_130), .A2(n_246), .B1(n_928), .B2(n_929), .Y(n_1286) );
AO22x2_ASAP7_75t_L g1307 ( .A1(n_131), .A2(n_1308), .B1(n_1309), .B2(n_1350), .Y(n_1307) );
INVxp67_ASAP7_75t_SL g1308 ( .A(n_131), .Y(n_1308) );
INVx1_ASAP7_75t_L g1952 ( .A(n_133), .Y(n_1952) );
XNOR2xp5_ASAP7_75t_L g1264 ( .A(n_134), .B(n_1265), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_135), .A2(n_299), .B1(n_1138), .B2(n_1360), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g1377 ( .A1(n_135), .A2(n_299), .B1(n_612), .B2(n_613), .C(n_715), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_136), .A2(n_217), .B1(n_540), .B2(n_542), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_136), .A2(n_217), .B1(n_1078), .B2(n_1138), .Y(n_1343) );
INVx1_ASAP7_75t_L g1997 ( .A(n_137), .Y(n_1997) );
AOI221xp5_ASAP7_75t_L g2009 ( .A1(n_137), .A2(n_150), .B1(n_722), .B2(n_944), .C(n_2010), .Y(n_2009) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_138), .A2(n_208), .B1(n_460), .B2(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1485 ( .A(n_138), .Y(n_1485) );
INVx1_ASAP7_75t_L g1549 ( .A(n_139), .Y(n_1549) );
OA22x2_ASAP7_75t_L g966 ( .A1(n_140), .A2(n_967), .B1(n_1046), .B2(n_1047), .Y(n_966) );
INVxp67_ASAP7_75t_SL g1047 ( .A(n_140), .Y(n_1047) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_141), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g751 ( .A(n_142), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g1482 ( .A1(n_143), .A2(n_323), .B1(n_636), .B2(n_1121), .C(n_1122), .Y(n_1482) );
INVx1_ASAP7_75t_L g1523 ( .A(n_144), .Y(n_1523) );
INVx1_ASAP7_75t_L g603 ( .A(n_146), .Y(n_603) );
INVx1_ASAP7_75t_L g1592 ( .A(n_147), .Y(n_1592) );
INVx1_ASAP7_75t_L g1180 ( .A(n_148), .Y(n_1180) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_148), .A2(n_335), .B1(n_1078), .B2(n_1207), .Y(n_1206) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_149), .Y(n_1063) );
INVx1_ASAP7_75t_L g2006 ( .A(n_150), .Y(n_2006) );
OAI22xp5_ASAP7_75t_L g1614 ( .A1(n_151), .A2(n_304), .B1(n_583), .B2(n_588), .Y(n_1614) );
AOI22xp33_ASAP7_75t_L g1622 ( .A1(n_151), .A2(n_304), .B1(n_1623), .B2(n_1624), .Y(n_1622) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_152), .A2(n_212), .B1(n_489), .B2(n_491), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_152), .A2(n_212), .B1(n_583), .B2(n_588), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_153), .Y(n_438) );
INVx1_ASAP7_75t_L g1477 ( .A(n_154), .Y(n_1477) );
OAI22xp33_ASAP7_75t_L g1488 ( .A1(n_154), .A2(n_323), .B1(n_954), .B2(n_957), .Y(n_1488) );
INVx1_ASAP7_75t_L g607 ( .A(n_155), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g987 ( .A(n_156), .Y(n_987) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_157), .Y(n_632) );
AOI22xp5_ASAP7_75t_SL g1740 ( .A1(n_158), .A2(n_174), .B1(n_1686), .B2(n_1694), .Y(n_1740) );
INVx1_ASAP7_75t_L g1328 ( .A(n_159), .Y(n_1328) );
XOR2xp5_ASAP7_75t_L g817 ( .A(n_160), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g1690 ( .A(n_162), .Y(n_1690) );
INVx1_ASAP7_75t_L g1175 ( .A(n_163), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_163), .A2(n_206), .B1(n_440), .B2(n_1199), .Y(n_1208) );
CKINVDCx16_ASAP7_75t_R g1732 ( .A(n_165), .Y(n_1732) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_166), .A2(n_327), .B1(n_1401), .B2(n_1417), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_166), .A2(n_327), .B1(n_771), .B2(n_782), .Y(n_1420) );
INVx1_ASAP7_75t_L g1426 ( .A(n_168), .Y(n_1426) );
INVx1_ASAP7_75t_L g717 ( .A(n_169), .Y(n_717) );
INVx1_ASAP7_75t_L g1106 ( .A(n_170), .Y(n_1106) );
INVx1_ASAP7_75t_L g1949 ( .A(n_171), .Y(n_1949) );
AOI221xp5_ASAP7_75t_L g1974 ( .A1(n_171), .A2(n_224), .B1(n_771), .B2(n_861), .C(n_1975), .Y(n_1974) );
INVx1_ASAP7_75t_L g1691 ( .A(n_172), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_172), .B(n_1689), .Y(n_1696) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_173), .A2(n_324), .B1(n_627), .B2(n_628), .C(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g658 ( .A(n_173), .Y(n_658) );
INVx1_ASAP7_75t_L g1939 ( .A(n_175), .Y(n_1939) );
AOI21xp33_ASAP7_75t_L g1971 ( .A1(n_175), .A2(n_1364), .B(n_1972), .Y(n_1971) );
INVx2_ASAP7_75t_L g393 ( .A(n_176), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g1996 ( .A(n_177), .Y(n_1996) );
INVx1_ASAP7_75t_L g1650 ( .A(n_178), .Y(n_1650) );
INVx1_ASAP7_75t_L g1940 ( .A(n_179), .Y(n_1940) );
AOI22xp33_ASAP7_75t_L g1970 ( .A1(n_179), .A2(n_247), .B1(n_792), .B2(n_1200), .Y(n_1970) );
INVx1_ASAP7_75t_L g1168 ( .A(n_180), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_181), .A2(n_289), .B1(n_627), .B2(n_1339), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_181), .A2(n_289), .B1(n_473), .B2(n_491), .Y(n_1344) );
INVx1_ASAP7_75t_L g1572 ( .A(n_182), .Y(n_1572) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_183), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_184), .A2(n_370), .B1(n_1199), .B2(n_1457), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1464 ( .A1(n_184), .A2(n_370), .B1(n_583), .B2(n_588), .Y(n_1464) );
INVx1_ASAP7_75t_L g415 ( .A(n_185), .Y(n_415) );
BUFx3_ASAP7_75t_L g435 ( .A(n_185), .Y(n_435) );
INVx1_ASAP7_75t_L g1414 ( .A(n_186), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_186), .A2(n_280), .B1(n_431), .B2(n_498), .Y(n_1423) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_187), .Y(n_1006) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_188), .Y(n_1383) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_189), .A2(n_351), .B1(n_447), .B2(n_460), .Y(n_1239) );
INVx1_ASAP7_75t_L g1255 ( .A(n_189), .Y(n_1255) );
INVx1_ASAP7_75t_L g1116 ( .A(n_190), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_191), .Y(n_993) );
INVxp33_ASAP7_75t_SL g824 ( .A(n_192), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g860 ( .A1(n_192), .A2(n_316), .B1(n_799), .B2(n_861), .C(n_863), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_193), .A2(n_361), .B1(n_635), .B2(n_636), .C(n_715), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_193), .A2(n_213), .B1(n_954), .B2(n_957), .Y(n_1263) );
INVx1_ASAP7_75t_L g1295 ( .A(n_194), .Y(n_1295) );
OAI22xp33_ASAP7_75t_L g1304 ( .A1(n_194), .A2(n_196), .B1(n_954), .B2(n_957), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_195), .A2(n_341), .B1(n_928), .B2(n_929), .Y(n_1074) );
INVx1_ASAP7_75t_L g1086 ( .A(n_195), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_196), .A2(n_234), .B1(n_635), .B2(n_636), .C(n_947), .Y(n_1298) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_197), .A2(n_271), .B1(n_1151), .B2(n_1170), .C(n_1171), .Y(n_1169) );
INVx1_ASAP7_75t_L g1178 ( .A(n_197), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g2015 ( .A1(n_199), .A2(n_342), .B1(n_1401), .B2(n_1611), .Y(n_2015) );
AOI22xp33_ASAP7_75t_L g2032 ( .A1(n_199), .A2(n_342), .B1(n_1510), .B2(n_2033), .Y(n_2032) );
CKINVDCx5p33_ASAP7_75t_R g1368 ( .A(n_201), .Y(n_1368) );
AOI22xp33_ASAP7_75t_SL g1365 ( .A1(n_202), .A2(n_373), .B1(n_440), .B2(n_1136), .Y(n_1365) );
INVx1_ASAP7_75t_L g1372 ( .A(n_202), .Y(n_1372) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_203), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g1498 ( .A1(n_204), .A2(n_216), .B1(n_774), .B2(n_777), .C(n_793), .Y(n_1498) );
INVx1_ASAP7_75t_L g1522 ( .A(n_204), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g946 ( .A1(n_205), .A2(n_374), .B1(n_545), .B2(n_612), .C(n_947), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g953 ( .A1(n_205), .A2(n_308), .B1(n_954), .B2(n_957), .Y(n_953) );
INVx1_ASAP7_75t_L g1176 ( .A(n_206), .Y(n_1176) );
INVx1_ASAP7_75t_L g1237 ( .A(n_207), .Y(n_1237) );
INVx1_ASAP7_75t_L g1484 ( .A(n_208), .Y(n_1484) );
INVx1_ASAP7_75t_L g1601 ( .A(n_210), .Y(n_1601) );
INVx1_ASAP7_75t_L g1568 ( .A(n_211), .Y(n_1568) );
INVx1_ASAP7_75t_L g1251 ( .A(n_213), .Y(n_1251) );
INVx1_ASAP7_75t_L g1391 ( .A(n_214), .Y(n_1391) );
INVx1_ASAP7_75t_L g1427 ( .A(n_215), .Y(n_1427) );
INVx1_ASAP7_75t_L g1520 ( .A(n_216), .Y(n_1520) );
INVx1_ASAP7_75t_L g418 ( .A(n_218), .Y(n_418) );
INVx1_ASAP7_75t_L g469 ( .A(n_218), .Y(n_469) );
INVxp33_ASAP7_75t_L g1153 ( .A(n_219), .Y(n_1153) );
INVx1_ASAP7_75t_L g2002 ( .A(n_220), .Y(n_2002) );
OAI221xp5_ASAP7_75t_L g2013 ( .A1(n_220), .A2(n_253), .B1(n_555), .B2(n_1408), .C(n_2014), .Y(n_2013) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_221), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g1791 ( .A(n_223), .Y(n_1791) );
INVx1_ASAP7_75t_L g1951 ( .A(n_224), .Y(n_1951) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_225), .Y(n_755) );
INVx1_ASAP7_75t_L g1411 ( .A(n_226), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_226), .A2(n_274), .B1(n_771), .B2(n_1200), .Y(n_1424) );
INVx1_ASAP7_75t_L g853 ( .A(n_227), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_228), .A2(n_350), .B1(n_1078), .B2(n_1362), .Y(n_1361) );
OAI221xp5_ASAP7_75t_L g1379 ( .A1(n_228), .A2(n_517), .B1(n_1380), .B2(n_1381), .C(n_1384), .Y(n_1379) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_229), .Y(n_761) );
INVx1_ASAP7_75t_L g911 ( .A(n_230), .Y(n_911) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_230), .A2(n_558), .B1(n_638), .B2(n_931), .C(n_937), .Y(n_930) );
XOR2xp5_ASAP7_75t_L g704 ( .A(n_231), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g1172 ( .A(n_232), .Y(n_1172) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_233), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_233), .A2(n_319), .B1(n_682), .B2(n_879), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g1303 ( .A1(n_234), .A2(n_337), .B1(n_422), .B2(n_1262), .Y(n_1303) );
INVx1_ASAP7_75t_L g742 ( .A(n_235), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_235), .A2(n_252), .B1(n_791), .B2(n_793), .C(n_795), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_236), .Y(n_599) );
INVx1_ASAP7_75t_L g1323 ( .A(n_237), .Y(n_1323) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_238), .Y(n_1072) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_238), .A2(n_447), .B1(n_460), .B2(n_497), .C(n_1088), .Y(n_1087) );
CKINVDCx5p33_ASAP7_75t_R g1954 ( .A(n_239), .Y(n_1954) );
INVx1_ASAP7_75t_L g720 ( .A(n_240), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_242), .Y(n_597) );
CKINVDCx14_ASAP7_75t_R g1715 ( .A(n_243), .Y(n_1715) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_244), .A2(n_267), .B1(n_555), .B2(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1433 ( .A(n_244), .Y(n_1433) );
INVx1_ASAP7_75t_L g1558 ( .A(n_245), .Y(n_1558) );
INVx1_ASAP7_75t_L g1280 ( .A(n_246), .Y(n_1280) );
INVx1_ASAP7_75t_L g1935 ( .A(n_247), .Y(n_1935) );
INVx1_ASAP7_75t_L g1591 ( .A(n_248), .Y(n_1591) );
INVx1_ASAP7_75t_L g1434 ( .A(n_249), .Y(n_1434) );
INVx1_ASAP7_75t_L g1603 ( .A(n_250), .Y(n_1603) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_251), .Y(n_1219) );
INVx1_ASAP7_75t_L g745 ( .A(n_252), .Y(n_745) );
INVx1_ASAP7_75t_L g2003 ( .A(n_253), .Y(n_2003) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_254), .Y(n_1167) );
OAI22xp33_ASAP7_75t_L g1556 ( .A1(n_255), .A2(n_347), .B1(n_921), .B2(n_923), .Y(n_1556) );
INVx1_ASAP7_75t_L g1576 ( .A(n_255), .Y(n_1576) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_257), .Y(n_622) );
INVx1_ASAP7_75t_L g1455 ( .A(n_259), .Y(n_1455) );
OAI211xp5_ASAP7_75t_SL g1474 ( .A1(n_259), .A2(n_517), .B(n_1475), .C(n_1483), .Y(n_1474) );
CKINVDCx16_ASAP7_75t_R g1094 ( .A(n_260), .Y(n_1094) );
INVx1_ASAP7_75t_L g1228 ( .A(n_261), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1244 ( .A1(n_261), .A2(n_558), .B1(n_638), .B2(n_1245), .C(n_1246), .Y(n_1244) );
INVx1_ASAP7_75t_L g1454 ( .A(n_262), .Y(n_1454) );
OAI221xp5_ASAP7_75t_L g1465 ( .A1(n_262), .A2(n_558), .B1(n_638), .B2(n_1466), .C(n_1472), .Y(n_1465) );
INVx1_ASAP7_75t_L g1551 ( .A(n_263), .Y(n_1551) );
OAI221xp5_ASAP7_75t_L g1561 ( .A1(n_263), .A2(n_558), .B1(n_638), .B2(n_1562), .C(n_1564), .Y(n_1561) );
INVx1_ASAP7_75t_L g1657 ( .A(n_264), .Y(n_1657) );
INVx1_ASAP7_75t_L g570 ( .A(n_265), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g1223 ( .A(n_266), .Y(n_1223) );
INVx1_ASAP7_75t_L g1432 ( .A(n_267), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_269), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_270), .A2(n_291), .B1(n_973), .B2(n_976), .Y(n_972) );
INVx1_ASAP7_75t_L g1029 ( .A(n_270), .Y(n_1029) );
INVx1_ASAP7_75t_L g1179 ( .A(n_271), .Y(n_1179) );
AOI21xp33_ASAP7_75t_L g1059 ( .A1(n_272), .A2(n_512), .B(n_613), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g1446 ( .A(n_273), .Y(n_1446) );
INVx1_ASAP7_75t_L g1412 ( .A(n_274), .Y(n_1412) );
INVx1_ASAP7_75t_L g1515 ( .A(n_275), .Y(n_1515) );
OAI211xp5_ASAP7_75t_L g979 ( .A1(n_276), .A2(n_561), .B(n_980), .C(n_984), .Y(n_979) );
INVx1_ASAP7_75t_L g1026 ( .A(n_276), .Y(n_1026) );
INVx1_ASAP7_75t_L g1100 ( .A(n_277), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_278), .Y(n_1513) );
INVx1_ASAP7_75t_L g1406 ( .A(n_280), .Y(n_1406) );
INVx1_ASAP7_75t_L g1545 ( .A(n_281), .Y(n_1545) );
CKINVDCx20_ASAP7_75t_R g1729 ( .A(n_282), .Y(n_1729) );
BUFx3_ASAP7_75t_L g414 ( .A(n_283), .Y(n_414) );
INVx1_ASAP7_75t_L g427 ( .A(n_283), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g1605 ( .A1(n_284), .A2(n_517), .B1(n_1606), .B2(n_1608), .C(n_1613), .Y(n_1605) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_285), .Y(n_600) );
INVx1_ASAP7_75t_L g1231 ( .A(n_286), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1248 ( .A1(n_286), .A2(n_517), .B(n_1249), .C(n_1254), .Y(n_1248) );
AO221x2_ASAP7_75t_L g1788 ( .A1(n_287), .A2(n_354), .B1(n_1755), .B2(n_1789), .C(n_1790), .Y(n_1788) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_288), .Y(n_1367) );
AO22x2_ASAP7_75t_L g1160 ( .A1(n_290), .A2(n_1161), .B1(n_1209), .B2(n_1210), .Y(n_1160) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_290), .Y(n_1209) );
AOI22xp5_ASAP7_75t_L g1706 ( .A1(n_290), .A2(n_293), .B1(n_1698), .B2(n_1702), .Y(n_1706) );
INVx1_ASAP7_75t_L g1028 ( .A(n_291), .Y(n_1028) );
INVx1_ASAP7_75t_L g1529 ( .A(n_292), .Y(n_1529) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_294), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_294), .B(n_356), .Y(n_511) );
AND2x2_ASAP7_75t_L g521 ( .A(n_294), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g549 ( .A(n_294), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_295), .Y(n_1382) );
AOI21xp33_ASAP7_75t_L g1066 ( .A1(n_296), .A2(n_635), .B(n_636), .Y(n_1066) );
INVx1_ASAP7_75t_L g1090 ( .A(n_296), .Y(n_1090) );
OR2x2_ASAP7_75t_L g417 ( .A(n_297), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g456 ( .A(n_297), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_298), .Y(n_1514) );
INVx1_ASAP7_75t_L g1252 ( .A(n_300), .Y(n_1252) );
OAI22xp33_ASAP7_75t_L g1261 ( .A1(n_300), .A2(n_361), .B1(n_422), .B2(n_1262), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_301), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g1053 ( .A(n_302), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_303), .Y(n_1013) );
INVx1_ASAP7_75t_L g1241 ( .A(n_305), .Y(n_1241) );
INVx1_ASAP7_75t_L g847 ( .A(n_306), .Y(n_847) );
INVx1_ASAP7_75t_L g1278 ( .A(n_307), .Y(n_1278) );
OAI211xp5_ASAP7_75t_L g1293 ( .A1(n_307), .A2(n_517), .B(n_1294), .C(n_1299), .Y(n_1293) );
INVx1_ASAP7_75t_L g942 ( .A(n_308), .Y(n_942) );
INVx1_ASAP7_75t_L g2024 ( .A(n_309), .Y(n_2024) );
AOI22xp33_ASAP7_75t_L g2037 ( .A1(n_309), .A2(n_338), .B1(n_474), .B2(n_2033), .Y(n_2037) );
INVx1_ASAP7_75t_L g420 ( .A(n_310), .Y(n_420) );
INVx1_ASAP7_75t_L g945 ( .A(n_311), .Y(n_945) );
OAI22xp33_ASAP7_75t_L g952 ( .A1(n_311), .A2(n_374), .B1(n_411), .B2(n_422), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_312), .Y(n_1061) );
AOI22xp5_ASAP7_75t_SL g1722 ( .A1(n_313), .A2(n_318), .B1(n_1702), .B2(n_1723), .Y(n_1722) );
INVx1_ASAP7_75t_L g915 ( .A(n_315), .Y(n_915) );
INVxp33_ASAP7_75t_L g826 ( .A(n_316), .Y(n_826) );
INVx1_ASAP7_75t_L g1320 ( .A(n_317), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_317), .A2(n_331), .B1(n_935), .B2(n_1124), .Y(n_1336) );
AOI22xp5_ASAP7_75t_L g1984 ( .A1(n_318), .A2(n_1985), .B1(n_1989), .B2(n_2038), .Y(n_1984) );
XNOR2xp5_ASAP7_75t_L g1992 ( .A(n_318), .B(n_1993), .Y(n_1992) );
INVxp33_ASAP7_75t_L g832 ( .A(n_319), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g1022 ( .A(n_320), .Y(n_1022) );
INVx1_ASAP7_75t_L g1642 ( .A(n_322), .Y(n_1642) );
INVx1_ASAP7_75t_L g650 ( .A(n_324), .Y(n_650) );
AOI22x1_ASAP7_75t_L g1352 ( .A1(n_325), .A2(n_1353), .B1(n_1354), .B2(n_1392), .Y(n_1352) );
INVxp67_ASAP7_75t_SL g1392 ( .A(n_325), .Y(n_1392) );
INVx1_ASAP7_75t_L g1316 ( .A(n_326), .Y(n_1316) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_328), .A2(n_372), .B1(n_1121), .B2(n_1122), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_328), .A2(n_372), .B1(n_776), .B2(n_1138), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_329), .Y(n_458) );
INVx1_ASAP7_75t_L g2031 ( .A(n_330), .Y(n_2031) );
INVx1_ASAP7_75t_L g1319 ( .A(n_331), .Y(n_1319) );
CKINVDCx5p33_ASAP7_75t_R g1959 ( .A(n_332), .Y(n_1959) );
CKINVDCx5p33_ASAP7_75t_R g1270 ( .A(n_333), .Y(n_1270) );
INVx1_ASAP7_75t_L g1607 ( .A(n_334), .Y(n_1607) );
INVx1_ASAP7_75t_L g1185 ( .A(n_335), .Y(n_1185) );
INVx1_ASAP7_75t_L g1589 ( .A(n_336), .Y(n_1589) );
INVx1_ASAP7_75t_L g1297 ( .A(n_337), .Y(n_1297) );
INVx1_ASAP7_75t_L g2023 ( .A(n_338), .Y(n_2023) );
INVx1_ASAP7_75t_L g577 ( .A(n_339), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_340), .Y(n_1271) );
INVx1_ASAP7_75t_L g1085 ( .A(n_341), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1693 ( .A(n_343), .B(n_381), .Y(n_1693) );
AND3x2_ASAP7_75t_L g1699 ( .A(n_343), .B(n_381), .C(n_1690), .Y(n_1699) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_344), .Y(n_925) );
INVx2_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g1548 ( .A(n_346), .Y(n_1548) );
INVx1_ASAP7_75t_L g1575 ( .A(n_347), .Y(n_1575) );
CKINVDCx5p33_ASAP7_75t_R g1221 ( .A(n_348), .Y(n_1221) );
INVx1_ASAP7_75t_L g1273 ( .A(n_349), .Y(n_1273) );
AOI21xp33_ASAP7_75t_L g1291 ( .A1(n_349), .A2(n_613), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1378 ( .A(n_350), .Y(n_1378) );
INVx1_ASAP7_75t_L g1257 ( .A(n_351), .Y(n_1257) );
XNOR2xp5_ASAP7_75t_L g1540 ( .A(n_352), .B(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g501 ( .A(n_353), .Y(n_501) );
OAI221xp5_ASAP7_75t_L g1942 ( .A1(n_355), .A2(n_357), .B1(n_724), .B2(n_731), .C(n_1943), .Y(n_1942) );
OAI221xp5_ASAP7_75t_L g1965 ( .A1(n_355), .A2(n_357), .B1(n_787), .B2(n_1966), .C(n_1968), .Y(n_1965) );
INVx1_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
INVx2_ASAP7_75t_L g522 ( .A(n_356), .Y(n_522) );
AO22x2_ASAP7_75t_L g593 ( .A1(n_358), .A2(n_594), .B1(n_698), .B2(n_699), .Y(n_593) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_358), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_359), .Y(n_971) );
INVx1_ASAP7_75t_L g856 ( .A(n_360), .Y(n_856) );
INVx1_ASAP7_75t_L g1071 ( .A(n_362), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_362), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1001 ( .A1(n_363), .A2(n_1002), .B(n_1004), .C(n_1008), .Y(n_1001) );
INVx1_ASAP7_75t_L g1043 ( .A(n_363), .Y(n_1043) );
INVxp33_ASAP7_75t_SL g822 ( .A(n_365), .Y(n_822) );
INVx1_ASAP7_75t_L g949 ( .A(n_366), .Y(n_949) );
INVx1_ASAP7_75t_L g2005 ( .A(n_367), .Y(n_2005) );
AOI21xp5_ASAP7_75t_L g2012 ( .A1(n_367), .A2(n_542), .B(n_545), .Y(n_2012) );
NOR2xp33_ASAP7_75t_L g1658 ( .A(n_368), .B(n_1659), .Y(n_1658) );
OAI211xp5_ASAP7_75t_SL g516 ( .A1(n_369), .A2(n_517), .B(n_527), .C(n_550), .Y(n_516) );
INVxp33_ASAP7_75t_SL g836 ( .A(n_371), .Y(n_836) );
INVx1_ASAP7_75t_L g1373 ( .A(n_373), .Y(n_1373) );
INVx1_ASAP7_75t_L g1471 ( .A(n_375), .Y(n_1471) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_397), .B(n_1677), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1988 ( .A(n_379), .B(n_385), .Y(n_1988) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1983 ( .A(n_380), .Y(n_1983) );
NAND2xp5_ASAP7_75t_L g2045 ( .A(n_380), .B(n_382), .Y(n_2045) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1982 ( .A(n_382), .B(n_1983), .Y(n_1982) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g968 ( .A(n_387), .B(n_493), .Y(n_968) );
OR2x6_ASAP7_75t_L g1097 ( .A(n_387), .B(n_493), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g573 ( .A(n_388), .B(n_396), .Y(n_573) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g613 ( .A(n_389), .B(n_614), .Y(n_613) );
INVx8_ASAP7_75t_L g970 ( .A(n_390), .Y(n_970) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_391), .Y(n_569) );
INVx1_ASAP7_75t_L g741 ( .A(n_391), .Y(n_741) );
OR2x2_ASAP7_75t_L g815 ( .A(n_391), .B(n_730), .Y(n_815) );
INVx2_ASAP7_75t_SL g835 ( .A(n_391), .Y(n_835) );
OR2x6_ASAP7_75t_L g1108 ( .A(n_391), .B(n_975), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1947 ( .A(n_391), .Y(n_1947) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g514 ( .A(n_393), .B(n_394), .Y(n_514) );
INVx1_ASAP7_75t_L g525 ( .A(n_393), .Y(n_525) );
INVx2_ASAP7_75t_L g532 ( .A(n_393), .Y(n_532) );
AND2x4_ASAP7_75t_L g538 ( .A(n_393), .B(n_526), .Y(n_538) );
INVx1_ASAP7_75t_L g565 ( .A(n_393), .Y(n_565) );
INVx2_ASAP7_75t_L g526 ( .A(n_394), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_394), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g553 ( .A(n_394), .Y(n_553) );
INVx1_ASAP7_75t_L g564 ( .A(n_394), .Y(n_564) );
INVx1_ASAP7_75t_L g587 ( .A(n_394), .Y(n_587) );
AND2x4_ASAP7_75t_L g988 ( .A(n_395), .B(n_553), .Y(n_988) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
XNOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_959), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_886), .B2(n_887), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22x1_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_702), .B1(n_884), .B2(n_885), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g884 ( .A(n_402), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_593), .B1(n_700), .B2(n_701), .Y(n_402) );
INVx1_ASAP7_75t_L g700 ( .A(n_403), .Y(n_700) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_500), .C(n_515), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_443), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_428), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_420), .B2(n_421), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_409), .A2(n_438), .B1(n_528), .B2(n_533), .C(n_539), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_410), .A2(n_421), .B1(n_1063), .B2(n_1065), .Y(n_1091) );
AOI222xp33_ASAP7_75t_L g1388 ( .A1(n_410), .A2(n_430), .B1(n_503), .B2(n_1382), .C1(n_1385), .C2(n_1389), .Y(n_1388) );
AOI22xp5_ASAP7_75t_L g1425 ( .A1(n_410), .A2(n_421), .B1(n_1426), .B2(n_1427), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1655 ( .A1(n_410), .A2(n_421), .B1(n_1656), .B2(n_1657), .Y(n_1655) );
CKINVDCx6p67_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
INVx2_ASAP7_75t_L g782 ( .A(n_412), .Y(n_782) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_412), .B(n_416), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_412), .A2(n_898), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g477 ( .A(n_413), .Y(n_477) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_413), .Y(n_660) );
INVx1_ASAP7_75t_L g683 ( .A(n_413), .Y(n_683) );
BUFx6f_ASAP7_75t_L g1200 ( .A(n_413), .Y(n_1200) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g436 ( .A(n_414), .Y(n_436) );
AND2x2_ASAP7_75t_L g483 ( .A(n_414), .B(n_435), .Y(n_483) );
INVx1_ASAP7_75t_L g425 ( .A(n_415), .Y(n_425) );
OR2x6_ASAP7_75t_L g422 ( .A(n_416), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
OR2x2_ASAP7_75t_L g954 ( .A(n_416), .B(n_955), .Y(n_954) );
OR2x2_ASAP7_75t_L g957 ( .A(n_416), .B(n_958), .Y(n_957) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx2_ASAP7_75t_L g772 ( .A(n_417), .Y(n_772) );
OR2x2_ASAP7_75t_L g809 ( .A(n_417), .B(n_679), .Y(n_809) );
OR2x2_ASAP7_75t_L g811 ( .A(n_417), .B(n_477), .Y(n_811) );
INVx1_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
AND2x4_ASAP7_75t_L g712 ( .A(n_419), .B(n_521), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g1390 ( .A1(n_421), .A2(n_439), .B1(n_1383), .B2(n_1391), .Y(n_1390) );
CKINVDCx6p67_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_423), .A2(n_677), .B1(n_911), .B2(n_912), .Y(n_910) );
BUFx3_ASAP7_75t_L g1025 ( .A(n_423), .Y(n_1025) );
INVx1_ASAP7_75t_L g2030 ( .A(n_423), .Y(n_2030) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g692 ( .A(n_424), .Y(n_692) );
INVx1_ASAP7_75t_L g908 ( .A(n_424), .Y(n_908) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_424), .Y(n_1225) );
BUFx4f_ASAP7_75t_L g1230 ( .A(n_424), .Y(n_1230) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OR2x2_ASAP7_75t_L g679 ( .A(n_425), .B(n_426), .Y(n_679) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g442 ( .A(n_427), .B(n_435), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_438), .B2(n_439), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g1089 ( .A1(n_430), .A2(n_439), .B1(n_503), .B2(n_1061), .C1(n_1068), .C2(n_1090), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g1428 ( .A1(n_430), .A2(n_439), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
AOI221xp5_ASAP7_75t_L g1590 ( .A1(n_430), .A2(n_439), .B1(n_1591), .B2(n_1592), .C(n_1593), .Y(n_1590) );
AOI22xp33_ASAP7_75t_L g1652 ( .A1(n_430), .A2(n_439), .B1(n_1653), .B2(n_1654), .Y(n_1652) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_437), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g799 ( .A(n_432), .Y(n_799) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g479 ( .A(n_433), .Y(n_479) );
INVx6_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
AND2x2_ASAP7_75t_L g504 ( .A(n_433), .B(n_453), .Y(n_504) );
AND2x4_ASAP7_75t_L g655 ( .A(n_433), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g463 ( .A(n_434), .Y(n_463) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g450 ( .A(n_436), .Y(n_450) );
AND2x2_ASAP7_75t_L g439 ( .A(n_437), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_441), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g1358 ( .A(n_441), .Y(n_1358) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g473 ( .A(n_442), .Y(n_473) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_442), .Y(n_490) );
AND2x6_ASAP7_75t_L g651 ( .A(n_442), .B(n_652), .Y(n_651) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_442), .Y(n_687) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_442), .Y(n_771) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_442), .Y(n_792) );
BUFx3_ASAP7_75t_L g899 ( .A(n_442), .Y(n_899) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_442), .Y(n_1135) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_464), .C(n_495), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_458), .B2(n_459), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_445), .A2(n_458), .B1(n_551), .B2(n_554), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g1587 ( .A1(n_446), .A2(n_459), .B1(n_893), .B2(n_1588), .C(n_1589), .Y(n_1587) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g922 ( .A(n_447), .Y(n_922) );
HB1xp67_ASAP7_75t_L g1460 ( .A(n_447), .Y(n_1460) );
INVx2_ASAP7_75t_L g1662 ( .A(n_447), .Y(n_1662) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g786 ( .A(n_449), .Y(n_786) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g667 ( .A(n_450), .Y(n_667) );
INVx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_L g460 ( .A(n_452), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g499 ( .A(n_452), .Y(n_499) );
OR2x2_ASAP7_75t_L g923 ( .A(n_452), .B(n_461), .Y(n_923) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
AND2x4_ASAP7_75t_L g785 ( .A(n_453), .B(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g788 ( .A(n_453), .B(n_462), .Y(n_788) );
INVx1_ASAP7_75t_L g805 ( .A(n_453), .Y(n_805) );
AND2x4_ASAP7_75t_L g1967 ( .A(n_453), .B(n_786), .Y(n_1967) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x4_ASAP7_75t_L g494 ( .A(n_455), .B(n_469), .Y(n_494) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g468 ( .A(n_456), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g648 ( .A(n_456), .Y(n_648) );
INVx1_ASAP7_75t_L g653 ( .A(n_456), .Y(n_653) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_456), .Y(n_657) );
OR2x6_ASAP7_75t_L g764 ( .A(n_457), .B(n_547), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g1366 ( .A1(n_459), .A2(n_893), .B1(n_922), .B2(n_1367), .C(n_1368), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1431 ( .A1(n_459), .A2(n_893), .B1(n_922), .B2(n_1432), .C(n_1433), .Y(n_1431) );
AOI22xp5_ASAP7_75t_L g1661 ( .A1(n_459), .A2(n_1662), .B1(n_1663), .B2(n_1664), .Y(n_1661) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g871 ( .A(n_461), .B(n_805), .Y(n_871) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x6_ASAP7_75t_L g668 ( .A(n_463), .B(n_653), .Y(n_668) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_472), .A3(n_478), .B1(n_484), .B2(n_488), .B3(n_492), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_465), .A2(n_697), .B1(n_1077), .B2(n_1083), .C(n_1087), .Y(n_1076) );
INVx1_ASAP7_75t_L g2026 ( .A(n_465), .Y(n_2026) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_466), .A2(n_675), .B1(n_689), .B2(n_695), .Y(n_674) );
OAI22xp5_ASAP7_75t_SL g1444 ( .A1(n_466), .A2(n_919), .B1(n_1445), .B2(n_1453), .Y(n_1444) );
CKINVDCx5p33_ASAP7_75t_R g1616 ( .A(n_466), .Y(n_1616) );
CKINVDCx5p33_ASAP7_75t_R g1666 ( .A(n_466), .Y(n_1666) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
OR2x2_ASAP7_75t_L g896 ( .A(n_467), .B(n_470), .Y(n_896) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g797 ( .A(n_468), .Y(n_797) );
INVx1_ASAP7_75t_L g877 ( .A(n_468), .Y(n_877) );
INVx1_ASAP7_75t_L g1204 ( .A(n_468), .Y(n_1204) );
BUFx3_ASAP7_75t_L g1976 ( .A(n_468), .Y(n_1976) );
INVx1_ASAP7_75t_L g641 ( .A(n_469), .Y(n_641) );
INVx2_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
BUFx2_ASAP7_75t_L g592 ( .A(n_470), .Y(n_592) );
AND2x4_ASAP7_75t_L g1119 ( .A(n_470), .B(n_573), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_470), .B(n_1204), .Y(n_1203) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g642 ( .A(n_471), .Y(n_642) );
OR2x6_ASAP7_75t_L g737 ( .A(n_471), .B(n_613), .Y(n_737) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g491 ( .A(n_475), .Y(n_491) );
INVx2_ASAP7_75t_SL g902 ( .A(n_475), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_475), .A2(n_686), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g869 ( .A(n_476), .Y(n_869) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g1018 ( .A(n_477), .Y(n_1018) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g1672 ( .A(n_481), .Y(n_1672) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_482), .Y(n_498) );
INVx1_ASAP7_75t_L g663 ( .A(n_482), .Y(n_663) );
AND2x4_ASAP7_75t_L g802 ( .A(n_482), .B(n_772), .Y(n_802) );
INVx1_ASAP7_75t_L g1142 ( .A(n_482), .Y(n_1142) );
BUFx4f_ASAP7_75t_L g1360 ( .A(n_482), .Y(n_1360) );
BUFx3_ASAP7_75t_L g1621 ( .A(n_482), .Y(n_1621) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_483), .Y(n_673) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g774 ( .A(n_486), .Y(n_774) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g649 ( .A(n_487), .Y(n_649) );
INVx2_ASAP7_75t_L g880 ( .A(n_487), .Y(n_880) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_487), .Y(n_1081) );
INVx2_ASAP7_75t_L g1139 ( .A(n_487), .Y(n_1139) );
INVx1_ASAP7_75t_L g1207 ( .A(n_487), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1364 ( .A(n_487), .Y(n_1364) );
INVx1_ASAP7_75t_L g1671 ( .A(n_487), .Y(n_1671) );
BUFx4f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g958 ( .A(n_490), .Y(n_958) );
BUFx2_ASAP7_75t_L g1450 ( .A(n_490), .Y(n_1450) );
AOI33xp33_ASAP7_75t_L g1132 ( .A1(n_492), .A2(n_1133), .A3(n_1134), .B1(n_1137), .B2(n_1140), .B3(n_1143), .Y(n_1132) );
NAND3xp33_ASAP7_75t_L g1205 ( .A(n_492), .B(n_1206), .C(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g1238 ( .A(n_492), .Y(n_1238) );
INVx1_ASAP7_75t_L g1349 ( .A(n_492), .Y(n_1349) );
AOI33xp33_ASAP7_75t_L g1356 ( .A1(n_492), .A2(n_1133), .A3(n_1357), .B1(n_1359), .B2(n_1361), .B3(n_1365), .Y(n_1356) );
AOI33xp33_ASAP7_75t_L g1419 ( .A1(n_492), .A2(n_1202), .A3(n_1420), .B1(n_1421), .B2(n_1423), .B3(n_1424), .Y(n_1419) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x4_ASAP7_75t_L g503 ( .A(n_493), .B(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g697 ( .A(n_493), .B(n_494), .Y(n_697) );
INVx2_ASAP7_75t_L g778 ( .A(n_494), .Y(n_778) );
INVx2_ASAP7_75t_SL g865 ( .A(n_494), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g1972 ( .A(n_494), .Y(n_1972) );
NAND3xp33_ASAP7_75t_SL g1660 ( .A(n_495), .B(n_1661), .C(n_1665), .Y(n_1660) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_498), .Y(n_688) );
BUFx2_ASAP7_75t_SL g876 ( .A(n_498), .Y(n_876) );
AND2x2_ASAP7_75t_L g893 ( .A(n_499), .B(n_894), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_502), .B(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_502), .B(n_1241), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_502), .B(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1397 ( .A(n_502), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_502), .B(n_1462), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_502), .B(n_1558), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_502), .B(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1659 ( .A(n_502), .Y(n_1659) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
INVx2_ASAP7_75t_L g816 ( .A(n_503), .Y(n_816) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g767 ( .A(n_506), .Y(n_767) );
INVx1_ASAP7_75t_L g598 ( .A(n_507), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AND2x2_ASAP7_75t_L g551 ( .A(n_508), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_508), .B(n_552), .Y(n_1256) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x6_ASAP7_75t_L g555 ( .A(n_509), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g580 ( .A(n_509), .B(n_581), .Y(n_580) );
OR2x6_ASAP7_75t_L g638 ( .A(n_509), .B(n_581), .Y(n_638) );
INVx1_ASAP7_75t_L g1073 ( .A(n_509), .Y(n_1073) );
INVx1_ASAP7_75t_L g1409 ( .A(n_509), .Y(n_1409) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_512), .Y(n_1121) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g635 ( .A(n_513), .Y(n_635) );
INVx2_ASAP7_75t_SL g719 ( .A(n_513), .Y(n_719) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_514), .Y(n_544) );
OAI31xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_557), .A3(n_582), .B(n_590), .Y(n_515) );
INVx8_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI222xp33_ASAP7_75t_L g596 ( .A1(n_518), .A2(n_559), .B1(n_597), .B2(n_598), .C1(n_599), .C2(n_600), .Y(n_596) );
AOI221xp5_ASAP7_75t_SL g1399 ( .A1(n_518), .A2(n_1400), .B1(n_1403), .B2(n_1406), .C(n_1407), .Y(n_1399) );
AOI221xp5_ASAP7_75t_L g1631 ( .A1(n_518), .A2(n_1632), .B1(n_1635), .B2(n_1639), .C(n_1640), .Y(n_1631) );
AOI222xp33_ASAP7_75t_L g2019 ( .A1(n_518), .A2(n_559), .B1(n_598), .B2(n_1996), .C1(n_2020), .C2(n_2021), .Y(n_2019) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
AND2x4_ASAP7_75t_L g589 ( .A(n_519), .B(n_536), .Y(n_589) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g559 ( .A(n_521), .B(n_544), .Y(n_559) );
AND2x2_ASAP7_75t_L g584 ( .A(n_521), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g548 ( .A(n_522), .Y(n_548) );
INVx1_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
INVx1_ASAP7_75t_L g541 ( .A(n_523), .Y(n_541) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g715 ( .A(n_524), .Y(n_715) );
BUFx6f_ASAP7_75t_L g947 ( .A(n_524), .Y(n_947) );
AND2x4_ASAP7_75t_L g981 ( .A(n_524), .B(n_982), .Y(n_981) );
BUFx6f_ASAP7_75t_L g1131 ( .A(n_524), .Y(n_1131) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_524), .Y(n_1183) );
INVx1_ASAP7_75t_L g2018 ( .A(n_524), .Y(n_2018) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g1609 ( .A(n_529), .Y(n_1609) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_530), .Y(n_933) );
INVx1_ASAP7_75t_L g1250 ( .A(n_530), .Y(n_1250) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g617 ( .A(n_531), .Y(n_617) );
INVx1_ASAP7_75t_L g750 ( .A(n_531), .Y(n_750) );
INVx1_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
AND2x4_ASAP7_75t_L g585 ( .A(n_532), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_535), .A2(n_940), .B1(n_1013), .B2(n_1016), .Y(n_1035) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g1417 ( .A(n_537), .Y(n_1417) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g579 ( .A(n_538), .Y(n_579) );
INVx3_ASAP7_75t_L g621 ( .A(n_538), .Y(n_621) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_538), .Y(n_630) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g1405 ( .A(n_541), .Y(n_1405) );
A2O1A1Ixp33_ASAP7_75t_L g1384 ( .A1(n_542), .A2(n_1073), .B(n_1385), .C(n_1386), .Y(n_1384) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g985 ( .A(n_543), .Y(n_985) );
INVx2_ASAP7_75t_SL g1292 ( .A(n_543), .Y(n_1292) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_544), .Y(n_612) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_544), .Y(n_1404) );
INVx1_ASAP7_75t_L g1569 ( .A(n_545), .Y(n_1569) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g636 ( .A(n_547), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g983 ( .A(n_548), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_551), .A2(n_554), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_551), .A2(n_554), .B1(n_949), .B2(n_950), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_551), .A2(n_554), .B1(n_1484), .B2(n_1485), .Y(n_1483) );
AOI22xp5_ASAP7_75t_L g1613 ( .A1(n_551), .A2(n_554), .B1(n_1588), .B2(n_1589), .Y(n_1613) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g728 ( .A(n_553), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_553), .A2(n_733), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_554), .A2(n_1255), .B1(n_1256), .B2(n_1257), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_554), .A2(n_1256), .B1(n_1300), .B2(n_1301), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_554), .A2(n_1256), .B1(n_1575), .B2(n_1576), .Y(n_1574) );
CKINVDCx11_ASAP7_75t_R g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g733 ( .A(n_556), .Y(n_733) );
CKINVDCx6p67_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g1374 ( .A1(n_559), .A2(n_1375), .B1(n_1377), .B2(n_1378), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1413 ( .A1(n_559), .A2(n_637), .B1(n_1414), .B2(n_1415), .C(n_1416), .Y(n_1413) );
AOI221xp5_ASAP7_75t_L g1644 ( .A1(n_559), .A2(n_637), .B1(n_1645), .B2(n_1647), .C(n_1650), .Y(n_1644) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_566), .B1(n_567), .B2(n_570), .C(n_571), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g1945 ( .A1(n_561), .A2(n_1946), .B1(n_1948), .B2(n_1949), .Y(n_1945) );
OAI22xp33_ASAP7_75t_L g1958 ( .A1(n_561), .A2(n_1473), .B1(n_1959), .B2(n_1960), .Y(n_1958) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g581 ( .A(n_563), .Y(n_581) );
INVx2_ASAP7_75t_L g633 ( .A(n_563), .Y(n_633) );
INVx3_ASAP7_75t_L g1058 ( .A(n_563), .Y(n_1058) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_564), .B(n_565), .Y(n_610) );
INVx1_ASAP7_75t_L g991 ( .A(n_565), .Y(n_991) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_569), .A2(n_571), .B1(n_609), .B2(n_906), .C(n_909), .Y(n_937) );
OAI22xp33_ASAP7_75t_L g1032 ( .A1(n_569), .A2(n_1020), .B1(n_1022), .B2(n_1033), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_569), .A2(n_854), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
BUFx2_ASAP7_75t_L g1473 ( .A(n_569), .Y(n_1473) );
OAI221xp5_ASAP7_75t_L g1602 ( .A1(n_569), .A2(n_609), .B1(n_1247), .B2(n_1603), .C(n_1604), .Y(n_1602) );
OAI221xp5_ASAP7_75t_L g1606 ( .A1(n_569), .A2(n_1058), .B1(n_1569), .B2(n_1592), .C(n_1607), .Y(n_1606) );
OAI221xp5_ASAP7_75t_L g1472 ( .A1(n_571), .A2(n_633), .B1(n_1446), .B2(n_1447), .C(n_1473), .Y(n_1472) );
OAI221xp5_ASAP7_75t_L g1564 ( .A1(n_571), .A2(n_834), .B1(n_1058), .B2(n_1548), .C(n_1549), .Y(n_1564) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_SL g1247 ( .A(n_573), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_576), .A2(n_1053), .B1(n_1054), .B2(n_1055), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_576), .A2(n_1061), .B1(n_1062), .B2(n_1063), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1381 ( .A1(n_576), .A2(n_1062), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
INVx1_ASAP7_75t_L g753 ( .A(n_578), .Y(n_753) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g978 ( .A(n_579), .Y(n_978) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_581), .Y(n_837) );
INVx1_ASAP7_75t_L g1034 ( .A(n_581), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_581), .B(n_1070), .Y(n_1069) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_584), .A2(n_589), .B1(n_602), .B2(n_603), .Y(n_601) );
INVx3_ASAP7_75t_L g928 ( .A(n_584), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_584), .A2(n_589), .B1(n_1372), .B2(n_1373), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_584), .A2(n_589), .B1(n_1411), .B2(n_1412), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1641 ( .A1(n_584), .A2(n_589), .B1(n_1642), .B2(n_1643), .Y(n_1641) );
AOI22xp33_ASAP7_75t_L g2022 ( .A1(n_584), .A2(n_589), .B1(n_2023), .B2(n_2024), .Y(n_2022) );
BUFx2_ASAP7_75t_L g627 ( .A(n_585), .Y(n_627) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_585), .Y(n_722) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_585), .B(n_975), .Y(n_1101) );
INVx1_ASAP7_75t_L g1125 ( .A(n_585), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g1376 ( .A(n_585), .Y(n_1376) );
BUFx6f_ASAP7_75t_L g1401 ( .A(n_585), .Y(n_1401) );
BUFx2_ASAP7_75t_L g1648 ( .A(n_585), .Y(n_1648) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx3_ASAP7_75t_L g929 ( .A(n_589), .Y(n_929) );
OAI31xp33_ASAP7_75t_L g1559 ( .A1(n_590), .A2(n_1560), .A3(n_1561), .B(n_1565), .Y(n_1559) );
AOI31xp33_ASAP7_75t_L g1963 ( .A1(n_590), .A2(n_1964), .A3(n_1973), .B(n_1978), .Y(n_1963) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI31xp33_ASAP7_75t_SL g1630 ( .A1(n_591), .A2(n_1631), .A3(n_1641), .B(n_1644), .Y(n_1630) );
CKINVDCx8_ASAP7_75t_R g591 ( .A(n_592), .Y(n_591) );
AOI221x1_ASAP7_75t_SL g594 ( .A1(n_592), .A2(n_595), .B1(n_639), .B2(n_643), .C(n_674), .Y(n_594) );
OAI31xp33_ASAP7_75t_SL g1463 ( .A1(n_592), .A2(n_1464), .A3(n_1465), .B(n_1474), .Y(n_1463) );
INVx2_ASAP7_75t_SL g701 ( .A(n_593), .Y(n_701) );
INVx1_ASAP7_75t_L g699 ( .A(n_594), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_601), .C(n_604), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_597), .A2(n_655), .B1(n_658), .B2(n_659), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_599), .A2(n_600), .B1(n_677), .B2(n_690), .C(n_693), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_626), .C(n_637), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_615), .B(n_623), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_611), .Y(n_606) );
BUFx3_ASAP7_75t_L g743 ( .A(n_608), .Y(n_743) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g855 ( .A(n_609), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g1246 ( .A1(n_609), .A2(n_759), .B1(n_1223), .B2(n_1226), .C(n_1247), .Y(n_1246) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_609), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_609), .B(n_1387), .Y(n_1386) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g1067 ( .A1(n_612), .A2(n_1068), .B(n_1069), .C(n_1073), .Y(n_1067) );
INVx1_ASAP7_75t_L g975 ( .A(n_614), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B1(n_619), .B2(n_622), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_616), .A2(n_847), .B1(n_848), .B2(n_851), .Y(n_846) );
BUFx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g941 ( .A(n_617), .Y(n_941) );
OR2x2_ASAP7_75t_L g973 ( .A(n_617), .B(n_974), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_619), .A2(n_940), .B1(n_1270), .B2(n_1271), .Y(n_1288) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g711 ( .A(n_620), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g1340 ( .A(n_620), .Y(n_1340) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g845 ( .A(n_621), .Y(n_845) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_621), .Y(n_850) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_622), .A2(n_676), .B1(n_680), .B2(n_681), .C(n_684), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_624), .A2(n_625), .B1(n_632), .B2(n_662), .C1(n_664), .C2(n_668), .Y(n_661) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_629), .A2(n_1037), .B1(n_1219), .B2(n_1221), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1535 ( .A1(n_629), .A2(n_746), .B1(n_1502), .B2(n_1514), .Y(n_1535) );
INVx2_ASAP7_75t_SL g1649 ( .A(n_629), .Y(n_1649) );
INVx4_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g756 ( .A(n_630), .Y(n_756) );
INVx2_ASAP7_75t_SL g1296 ( .A(n_630), .Y(n_1296) );
INVx2_ASAP7_75t_SL g1600 ( .A(n_630), .Y(n_1600) );
INVx2_ASAP7_75t_SL g1634 ( .A(n_630), .Y(n_1634) );
BUFx3_ASAP7_75t_L g1956 ( .A(n_630), .Y(n_1956) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_633), .B(n_634), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g758 ( .A1(n_633), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
OAI21xp33_ASAP7_75t_L g1064 ( .A1(n_633), .A2(n_1065), .B(n_1066), .Y(n_1064) );
NOR3xp33_ASAP7_75t_SL g2008 ( .A(n_637), .B(n_2009), .C(n_2013), .Y(n_2008) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI221x1_ASAP7_75t_L g1161 ( .A1(n_639), .A2(n_1096), .B1(n_1162), .B2(n_1173), .C(n_1186), .Y(n_1161) );
AOI221x1_ASAP7_75t_L g1309 ( .A1(n_639), .A2(n_1096), .B1(n_1310), .B2(n_1321), .C(n_1332), .Y(n_1309) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI221x1_ASAP7_75t_SL g1993 ( .A1(n_640), .A2(n_1258), .B1(n_1994), .B2(n_2007), .C(n_2025), .Y(n_1993) );
AND2x4_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_641), .B(n_642), .Y(n_1009) );
INVx2_ASAP7_75t_L g1259 ( .A(n_642), .Y(n_1259) );
NAND4xp25_ASAP7_75t_SL g643 ( .A(n_644), .B(n_654), .C(n_661), .D(n_669), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_650), .B2(n_651), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_646), .A2(n_659), .B1(n_1164), .B2(n_1165), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_646), .A2(n_655), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
AND2x4_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
AND2x6_ASAP7_75t_L g659 ( .A(n_647), .B(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_647), .B(n_649), .Y(n_1154) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_648), .B(n_1150), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_651), .A2(n_659), .B1(n_1156), .B2(n_1157), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g1166 ( .A1(n_651), .A2(n_655), .B1(n_1167), .B2(n_1168), .C(n_1169), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_651), .A2(n_659), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g2004 ( .A1(n_651), .A2(n_1154), .B1(n_2005), .B2(n_2006), .Y(n_2004) );
INVx1_ASAP7_75t_L g672 ( .A(n_652), .Y(n_672) );
INVx1_ASAP7_75t_L g999 ( .A(n_652), .Y(n_999) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_652), .B(n_776), .Y(n_1003) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx4_ASAP7_75t_L g1000 ( .A(n_655), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_655), .A2(n_1106), .B1(n_1153), .B2(n_1154), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1995 ( .A1(n_655), .A2(n_659), .B1(n_1996), .B2(n_1997), .Y(n_1995) );
AND2x4_ASAP7_75t_L g665 ( .A(n_656), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_SL g1007 ( .A(n_656), .B(n_666), .Y(n_1007) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx4_ASAP7_75t_L g996 ( .A(n_659), .Y(n_996) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_660), .Y(n_800) );
INVx1_ASAP7_75t_L g1030 ( .A(n_660), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_660), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g1236 ( .A(n_660), .Y(n_1236) );
INVx2_ASAP7_75t_L g1625 ( .A(n_660), .Y(n_1625) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g1998 ( .A1(n_664), .A2(n_668), .B1(n_1999), .B2(n_2000), .C1(n_2002), .C2(n_2003), .Y(n_1998) );
BUFx4f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g1150 ( .A(n_667), .Y(n_1150) );
AOI322xp5_ASAP7_75t_L g1004 ( .A1(n_668), .A2(n_687), .A3(n_987), .B1(n_993), .B2(n_1005), .C1(n_1006), .C2(n_1007), .Y(n_1004) );
INVx3_ASAP7_75t_L g1151 ( .A(n_668), .Y(n_1151) );
NAND4xp25_ASAP7_75t_L g1994 ( .A(n_669), .B(n_1995), .C(n_1998), .D(n_2004), .Y(n_1994) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx5_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
CKINVDCx8_ASAP7_75t_R g1008 ( .A(n_671), .Y(n_1008) );
AOI211xp5_ASAP7_75t_L g1145 ( .A1(n_671), .A2(n_1003), .B(n_1146), .C(n_1147), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_671), .B(n_1312), .Y(n_1311) );
AND2x4_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g1171 ( .A1(n_672), .A2(n_806), .B(n_1172), .Y(n_1171) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_673), .Y(n_776) );
INVx1_ASAP7_75t_L g794 ( .A(n_673), .Y(n_794) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_673), .Y(n_806) );
INVx2_ASAP7_75t_L g1079 ( .A(n_673), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1445 ( .A1(n_676), .A2(n_1446), .B1(n_1447), .B2(n_1448), .C(n_1449), .Y(n_1445) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g905 ( .A(n_679), .Y(n_905) );
INVx2_ASAP7_75t_L g956 ( .A(n_679), .Y(n_956) );
OR2x2_ASAP7_75t_L g998 ( .A(n_679), .B(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g694 ( .A(n_683), .Y(n_694) );
INVx1_ASAP7_75t_L g917 ( .A(n_683), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_683), .A2(n_875), .B1(n_1053), .B2(n_1055), .Y(n_1082) );
OAI22xp33_ASAP7_75t_L g1268 ( .A1(n_683), .A2(n_1269), .B1(n_1270), .B2(n_1271), .Y(n_1268) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g1015 ( .A(n_686), .Y(n_1015) );
INVx2_ASAP7_75t_SL g1623 ( .A(n_686), .Y(n_1623) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g1233 ( .A(n_687), .Y(n_1233) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_687), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1275 ( .A1(n_690), .A2(n_1276), .B1(n_1277), .B2(n_1278), .Y(n_1275) );
OAI221xp5_ASAP7_75t_L g1453 ( .A1(n_690), .A2(n_1276), .B1(n_1454), .B2(n_1455), .C(n_1456), .Y(n_1453) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_692), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
AOI33xp33_ASAP7_75t_L g1615 ( .A1(n_696), .A2(n_1616), .A3(n_1617), .B1(n_1619), .B2(n_1620), .B3(n_1622), .Y(n_1615) );
BUFx4f_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx4_ASAP7_75t_L g919 ( .A(n_697), .Y(n_919) );
BUFx4f_ASAP7_75t_L g1675 ( .A(n_697), .Y(n_1675) );
INVx1_ASAP7_75t_L g885 ( .A(n_702), .Y(n_885) );
AO22x2_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_817), .B2(n_883), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_765), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_723), .C(n_736), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_716), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_713), .B2(n_714), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_710), .A2(n_714), .B1(n_1519), .B2(n_1520), .Y(n_1518) );
BUFx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g823 ( .A(n_711), .Y(n_823) );
BUFx2_ASAP7_75t_L g1936 ( .A(n_711), .Y(n_1936) );
AND2x6_ASAP7_75t_L g714 ( .A(n_712), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g718 ( .A(n_712), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g721 ( .A(n_712), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g1941 ( .A(n_712), .B(n_722), .Y(n_1941) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_714), .A2(n_822), .B1(n_823), .B2(n_824), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g1934 ( .A1(n_714), .A2(n_1935), .B1(n_1936), .B2(n_1937), .Y(n_1934) );
NAND2x1p5_ASAP7_75t_L g735 ( .A(n_715), .B(n_729), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_721), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_718), .A2(n_721), .B1(n_826), .B2(n_827), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_718), .A2(n_721), .B1(n_1522), .B2(n_1523), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g1938 ( .A1(n_718), .A2(n_1939), .B1(n_1940), .B2(n_1941), .Y(n_1938) );
INVx1_ASAP7_75t_L g1637 ( .A(n_719), .Y(n_1637) );
BUFx2_ASAP7_75t_L g1646 ( .A(n_719), .Y(n_1646) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2x1_ASAP7_75t_SL g726 ( .A(n_727), .B(n_729), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g1387 ( .A1(n_727), .A2(n_990), .B1(n_1367), .B2(n_1368), .Y(n_1387) );
NAND2x1p5_ASAP7_75t_L g1408 ( .A(n_727), .B(n_1409), .Y(n_1408) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2x1p5_ASAP7_75t_L g732 ( .A(n_729), .B(n_733), .Y(n_732) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx4f_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx4f_ASAP7_75t_L g829 ( .A(n_732), .Y(n_829) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g1943 ( .A(n_735), .Y(n_1943) );
OAI33xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .A3(n_744), .B1(n_754), .B2(n_758), .B3(n_762), .Y(n_736) );
OAI33xp33_ASAP7_75t_L g830 ( .A1(n_737), .A2(n_762), .A3(n_831), .B1(n_838), .B2(n_846), .B3(n_852), .Y(n_830) );
OAI33xp33_ASAP7_75t_L g1031 ( .A1(n_737), .A2(n_1032), .A3(n_1035), .B1(n_1036), .B2(n_1041), .B3(n_1044), .Y(n_1031) );
INVx1_ASAP7_75t_L g1527 ( .A(n_737), .Y(n_1527) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g759 ( .A(n_741), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_751), .B2(n_752), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_746), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_746), .A2(n_756), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g840 ( .A(n_749), .Y(n_840) );
INVx2_ASAP7_75t_SL g1037 ( .A(n_749), .Y(n_1037) );
INVx2_ASAP7_75t_L g1563 ( .A(n_749), .Y(n_1563) );
BUFx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g1469 ( .A(n_750), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1562 ( .A1(n_752), .A2(n_1545), .B1(n_1546), .B2(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_755), .A2(n_770), .B1(n_773), .B2(n_779), .C(n_783), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_756), .A2(n_1250), .B1(n_1251), .B2(n_1252), .C(n_1253), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_757), .A2(n_760), .B1(n_808), .B2(n_810), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g1528 ( .A1(n_759), .A2(n_1529), .B1(n_1530), .B2(n_1531), .Y(n_1528) );
OAI221xp5_ASAP7_75t_L g1566 ( .A1(n_759), .A2(n_854), .B1(n_1567), .B2(n_1568), .C(n_1569), .Y(n_1566) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_761), .A2(n_790), .B1(n_798), .B2(n_801), .C(n_803), .Y(n_789) );
OAI33xp33_ASAP7_75t_L g1525 ( .A1(n_762), .A2(n_1526), .A3(n_1528), .B1(n_1532), .B2(n_1535), .B3(n_1536), .Y(n_1525) );
OAI33xp33_ASAP7_75t_L g1944 ( .A1(n_762), .A2(n_1526), .A3(n_1945), .B1(n_1950), .B2(n_1953), .B3(n_1958), .Y(n_1944) );
CKINVDCx8_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g1193 ( .A(n_763), .B(n_1194), .C(n_1196), .Y(n_1193) );
NAND3xp33_ASAP7_75t_L g1333 ( .A(n_763), .B(n_1334), .C(n_1336), .Y(n_1333) );
INVx5_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx6_ASAP7_75t_L g1045 ( .A(n_764), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B1(n_812), .B2(n_813), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_766), .A2(n_813), .B1(n_858), .B2(n_882), .Y(n_857) );
AOI31xp33_ASAP7_75t_L g1398 ( .A1(n_766), .A2(n_1399), .A3(n_1410), .B(n_1413), .Y(n_1398) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI31xp33_ASAP7_75t_L g926 ( .A1(n_767), .A2(n_927), .A3(n_930), .B(n_938), .Y(n_926) );
OAI31xp33_ASAP7_75t_L g1050 ( .A1(n_767), .A2(n_1051), .A3(n_1074), .B(n_1075), .Y(n_1050) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_789), .C(n_807), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_770), .A2(n_847), .B1(n_860), .B2(n_866), .C(n_870), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g1497 ( .A1(n_770), .A2(n_1498), .B1(n_1499), .B2(n_1502), .C(n_1503), .Y(n_1497) );
AOI21xp5_ASAP7_75t_L g1964 ( .A1(n_770), .A2(n_1954), .B(n_1965), .Y(n_1964) );
AND2x4_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
BUFx3_ASAP7_75t_L g780 ( .A(n_771), .Y(n_780) );
INVx1_ASAP7_75t_L g868 ( .A(n_771), .Y(n_868) );
INVx2_ASAP7_75t_SL g875 ( .A(n_771), .Y(n_875) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
BUFx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g914 ( .A(n_792), .Y(n_914) );
INVx1_ASAP7_75t_L g1458 ( .A(n_792), .Y(n_1458) );
BUFx2_ASAP7_75t_L g1506 ( .A(n_792), .Y(n_1506) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g894 ( .A(n_794), .Y(n_894) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g872 ( .A1(n_801), .A2(n_803), .B1(n_856), .B2(n_873), .C(n_878), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g1504 ( .A1(n_801), .A2(n_803), .B1(n_1505), .B2(n_1509), .C(n_1511), .Y(n_1504) );
AOI221xp5_ASAP7_75t_L g1973 ( .A1(n_801), .A2(n_803), .B1(n_1960), .B2(n_1974), .C(n_1977), .Y(n_1973) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AND2x4_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g862 ( .A(n_806), .Y(n_862) );
INVx1_ASAP7_75t_L g1508 ( .A(n_806), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_808), .A2(n_810), .B1(n_851), .B2(n_853), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_808), .A2(n_810), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1978 ( .A1(n_808), .A2(n_810), .B1(n_1957), .B2(n_1959), .Y(n_1978) );
INVx6_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx4_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_813), .A2(n_1495), .B1(n_1496), .B2(n_1515), .Y(n_1494) );
AOI21xp33_ASAP7_75t_L g1961 ( .A1(n_813), .A2(n_1962), .B(n_1963), .Y(n_1961) );
INVx5_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g883 ( .A(n_817), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_857), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_828), .C(n_830), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_825), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_836), .B2(n_837), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_833), .A2(n_853), .B1(n_854), .B2(n_856), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g1536 ( .A1(n_833), .A2(n_1290), .B1(n_1511), .B2(n_1513), .Y(n_1536) );
BUFx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g1466 ( .A1(n_842), .A2(n_1467), .B1(n_1470), .B2(n_1471), .Y(n_1466) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g936 ( .A(n_845), .Y(n_936) );
INVx2_ASAP7_75t_L g1054 ( .A(n_845), .Y(n_1054) );
INVx2_ASAP7_75t_L g1062 ( .A(n_845), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g1402 ( .A(n_845), .Y(n_1402) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g944 ( .A(n_850), .Y(n_944) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_850), .Y(n_1039) );
INVx2_ASAP7_75t_L g1195 ( .A(n_850), .Y(n_1195) );
INVx3_ASAP7_75t_L g1611 ( .A(n_850), .Y(n_1611) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g1530 ( .A(n_855), .Y(n_1530) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_872), .C(n_881), .Y(n_858) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g1501 ( .A(n_869), .Y(n_1501) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g1500 ( .A(n_875), .Y(n_1500) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
BUFx3_ASAP7_75t_L g1618 ( .A(n_880), .Y(n_1618) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AND4x1_ASAP7_75t_L g890 ( .A(n_891), .B(n_924), .C(n_926), .D(n_951), .Y(n_890) );
NOR3xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_895), .C(n_920), .Y(n_891) );
NOR3xp33_ASAP7_75t_SL g1542 ( .A(n_892), .B(n_1543), .C(n_1556), .Y(n_1542) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NOR3xp33_ASAP7_75t_L g1216 ( .A(n_893), .B(n_1217), .C(n_1239), .Y(n_1216) );
NOR3xp33_ASAP7_75t_L g1266 ( .A(n_893), .B(n_1267), .C(n_1282), .Y(n_1266) );
BUFx2_ASAP7_75t_L g1443 ( .A(n_893), .Y(n_1443) );
OAI33xp33_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .A3(n_904), .B1(n_910), .B2(n_913), .B3(n_919), .Y(n_895) );
OAI33xp33_ASAP7_75t_L g1011 ( .A1(n_896), .A2(n_919), .A3(n_1012), .B1(n_1019), .B2(n_1024), .B3(n_1027), .Y(n_1011) );
INVx1_ASAP7_75t_SL g1133 ( .A(n_896), .Y(n_1133) );
OAI33xp33_ASAP7_75t_L g1217 ( .A1(n_896), .A2(n_1218), .A3(n_1222), .B1(n_1227), .B2(n_1232), .B3(n_1238), .Y(n_1217) );
OAI33xp33_ASAP7_75t_L g1267 ( .A1(n_896), .A2(n_1238), .A3(n_1268), .B1(n_1272), .B2(n_1275), .B3(n_1279), .Y(n_1267) );
OAI33xp33_ASAP7_75t_L g1543 ( .A1(n_896), .A2(n_919), .A3(n_1544), .B1(n_1547), .B2(n_1550), .B3(n_1553), .Y(n_1543) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_900), .B1(n_901), .B2(n_903), .Y(n_897) );
OAI22xp33_ASAP7_75t_L g1218 ( .A1(n_898), .A2(n_1219), .B1(n_1220), .B2(n_1221), .Y(n_1218) );
INVx2_ASAP7_75t_SL g898 ( .A(n_899), .Y(n_898) );
BUFx3_ASAP7_75t_L g2033 ( .A(n_899), .Y(n_2033) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_900), .A2(n_903), .B1(n_932), .B2(n_934), .Y(n_931) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_907), .B2(n_909), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g1547 ( .A1(n_905), .A2(n_1025), .B1(n_1548), .B2(n_1549), .Y(n_1547) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g1314 ( .A(n_908), .Y(n_1314) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_916), .B2(n_918), .Y(n_913) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g2025 ( .A1(n_919), .A2(n_2026), .B1(n_2027), .B2(n_2034), .Y(n_2025) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_942), .B1(n_943), .B2(n_945), .C(n_946), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_947), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g1122 ( .A(n_947), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .Y(n_951) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx2_ASAP7_75t_L g1021 ( .A(n_956), .Y(n_1021) );
INVx2_ASAP7_75t_L g1276 ( .A(n_956), .Y(n_1276) );
HB1xp67_ASAP7_75t_L g2036 ( .A(n_956), .Y(n_2036) );
AOI22xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_1437), .B2(n_1676), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
OAI21x1_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_1393), .B(n_1435), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_963), .B(n_1436), .Y(n_1435) );
XNOR2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_1212), .Y(n_963) );
XNOR2x1_ASAP7_75t_L g964 ( .A(n_965), .B(n_1092), .Y(n_964) );
XNOR2x1_ASAP7_75t_L g965 ( .A(n_966), .B(n_1048), .Y(n_965) );
INVx1_ASAP7_75t_L g1046 ( .A(n_967), .Y(n_1046) );
OAI211xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B(n_994), .C(n_1010), .Y(n_967) );
AOI211xp5_ASAP7_75t_L g969 ( .A1(n_970), .A2(n_971), .B(n_972), .C(n_979), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_970), .A2(n_1105), .B1(n_1106), .B2(n_1107), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_970), .A2(n_1107), .B1(n_1167), .B2(n_1185), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_970), .A2(n_1317), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_971), .A2(n_1021), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
AOI322xp5_ASAP7_75t_L g984 ( .A1(n_974), .A2(n_985), .A3(n_986), .B1(n_987), .B2(n_988), .C1(n_989), .C2(n_993), .Y(n_984) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
AND2x4_ASAP7_75t_L g977 ( .A(n_975), .B(n_978), .Y(n_977) );
AND2x4_ASAP7_75t_L g1103 ( .A(n_975), .B(n_978), .Y(n_1103) );
INVx5_ASAP7_75t_SL g976 ( .A(n_977), .Y(n_976) );
NAND4xp25_ASAP7_75t_SL g1098 ( .A(n_980), .B(n_1099), .C(n_1104), .D(n_1109), .Y(n_1098) );
NAND4xp25_ASAP7_75t_SL g1173 ( .A(n_980), .B(n_1174), .C(n_1177), .D(n_1184), .Y(n_1173) );
NAND4xp25_ASAP7_75t_SL g1321 ( .A(n_980), .B(n_1322), .C(n_1325), .D(n_1329), .Y(n_1321) );
CKINVDCx11_ASAP7_75t_R g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVxp67_ASAP7_75t_L g992 ( .A(n_983), .Y(n_992) );
INVx2_ASAP7_75t_L g1115 ( .A(n_988), .Y(n_1115) );
AOI222xp33_ASAP7_75t_L g1177 ( .A1(n_988), .A2(n_989), .B1(n_1178), .B2(n_1179), .C1(n_1180), .C2(n_1181), .Y(n_1177) );
AOI222xp33_ASAP7_75t_L g1109 ( .A1(n_989), .A2(n_1110), .B1(n_1111), .B2(n_1113), .C1(n_1114), .C2(n_1116), .Y(n_1109) );
AOI222xp33_ASAP7_75t_L g1325 ( .A1(n_989), .A2(n_1111), .B1(n_1114), .B2(n_1326), .C1(n_1327), .C2(n_1328), .Y(n_1325) );
AND2x4_ASAP7_75t_L g989 ( .A(n_990), .B(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI31xp33_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_997), .A3(n_1001), .B(n_1009), .Y(n_994) );
INVx1_ASAP7_75t_L g1005 ( .A(n_999), .Y(n_1005) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_1006), .A2(n_1037), .B1(n_1038), .B2(n_1040), .Y(n_1036) );
INVx1_ASAP7_75t_SL g1158 ( .A(n_1009), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1031), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1014), .B1(n_1016), .B2(n_1017), .Y(n_1012) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
OAI22xp33_ASAP7_75t_SL g1019 ( .A1(n_1020), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1222 ( .A1(n_1021), .A2(n_1223), .B1(n_1224), .B2(n_1226), .Y(n_1222) );
OAI22xp33_ASAP7_75t_L g1227 ( .A1(n_1021), .A2(n_1228), .B1(n_1229), .B2(n_1231), .Y(n_1227) );
OAI22xp33_ASAP7_75t_L g1272 ( .A1(n_1021), .A2(n_1224), .B1(n_1273), .B2(n_1274), .Y(n_1272) );
OAI22xp33_ASAP7_75t_L g1550 ( .A1(n_1021), .A2(n_1025), .B1(n_1551), .B2(n_1552), .Y(n_1550) );
OAI221xp5_ASAP7_75t_L g2027 ( .A1(n_1021), .A2(n_2028), .B1(n_2029), .B2(n_2031), .C(n_2032), .Y(n_2027) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g2011 ( .A(n_1034), .Y(n_2011) );
OAI22xp5_ASAP7_75t_L g1598 ( .A1(n_1037), .A2(n_1599), .B1(n_1600), .B2(n_1601), .Y(n_1598) );
OAI22xp5_ASAP7_75t_L g1950 ( .A1(n_1038), .A2(n_1467), .B1(n_1951), .B2(n_1952), .Y(n_1950) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AOI33xp33_ASAP7_75t_L g1118 ( .A1(n_1045), .A2(n_1119), .A3(n_1120), .B1(n_1123), .B2(n_1127), .B3(n_1129), .Y(n_1118) );
NAND4xp25_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1076), .C(n_1089), .D(n_1091), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1056), .B1(n_1060), .B2(n_1064), .C(n_1067), .Y(n_1051) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1054), .Y(n_1128) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_1054), .Y(n_1189) );
OAI21xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B(n_1059), .Y(n_1056) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1062), .Y(n_1126) );
INVx1_ASAP7_75t_L g2001 ( .A(n_1078), .Y(n_2001) );
INVx3_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1079), .Y(n_1422) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
OA22x2_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1159), .B1(n_1160), .B2(n_1211), .Y(n_1092) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1093), .Y(n_1211) );
XNOR2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
AOI211xp5_ASAP7_75t_L g1095 ( .A1(n_1096), .A2(n_1098), .B(n_1117), .C(n_1144), .Y(n_1095) );
CKINVDCx16_ASAP7_75t_R g1096 ( .A(n_1097), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1101), .B1(n_1102), .B2(n_1103), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_1101), .A2(n_1103), .B1(n_1175), .B2(n_1176), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_1101), .A2(n_1103), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
INVx4_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx5_ASAP7_75t_L g1331 ( .A(n_1108), .Y(n_1331) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1638 ( .A(n_1112), .Y(n_1638) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
NAND2xp5_ASAP7_75t_SL g1117 ( .A(n_1118), .B(n_1132), .Y(n_1117) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_1119), .B(n_1188), .C(n_1190), .Y(n_1187) );
NAND3xp33_ASAP7_75t_L g1337 ( .A(n_1119), .B(n_1338), .C(n_1341), .Y(n_1337) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx2_ASAP7_75t_SL g1192 ( .A(n_1131), .Y(n_1192) );
HB1xp67_ASAP7_75t_L g1335 ( .A(n_1131), .Y(n_1335) );
BUFx6f_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
AOI31xp33_ASAP7_75t_SL g1144 ( .A1(n_1145), .A2(n_1152), .A3(n_1155), .B(n_1158), .Y(n_1144) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1149), .Y(n_1170) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1161), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1166), .Y(n_1162) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND4xp25_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1193), .C(n_1197), .D(n_1205), .Y(n_1186) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1189), .Y(n_1573) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NAND3xp33_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1201), .C(n_1202), .Y(n_1197) );
BUFx6f_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1200), .Y(n_1220) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1200), .Y(n_1452) );
BUFx3_ASAP7_75t_L g1510 ( .A(n_1200), .Y(n_1510) );
NAND3xp33_ASAP7_75t_L g1342 ( .A(n_1202), .B(n_1343), .C(n_1344), .Y(n_1342) );
INVx3_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
XNOR2xp5_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1305), .Y(n_1212) );
XOR2xp5_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1264), .Y(n_1213) );
AND4x1_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1240), .C(n_1242), .D(n_1260), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_1220), .A2(n_1233), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
INVx2_ASAP7_75t_SL g1224 ( .A(n_1225), .Y(n_1224) );
BUFx2_ASAP7_75t_L g1448 ( .A(n_1229), .Y(n_1448) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_SL g1969 ( .A(n_1230), .Y(n_1969) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1234), .B1(n_1235), .B2(n_1237), .Y(n_1232) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_1236), .Y(n_1235) );
OAI31xp33_ASAP7_75t_L g1242 ( .A1(n_1243), .A2(n_1244), .A3(n_1248), .B(n_1258), .Y(n_1242) );
OAI221xp5_ASAP7_75t_L g1294 ( .A1(n_1250), .A2(n_1295), .B1(n_1296), .B2(n_1297), .C(n_1298), .Y(n_1294) );
OAI31xp33_ASAP7_75t_L g1285 ( .A1(n_1258), .A2(n_1286), .A3(n_1287), .B(n_1293), .Y(n_1285) );
OAI21xp5_ASAP7_75t_L g1369 ( .A1(n_1258), .A2(n_1370), .B(n_1379), .Y(n_1369) );
OAI31xp33_ASAP7_75t_L g1596 ( .A1(n_1258), .A2(n_1597), .A3(n_1605), .B(n_1614), .Y(n_1596) );
BUFx8_ASAP7_75t_SL g1258 ( .A(n_1259), .Y(n_1258) );
INVx2_ASAP7_75t_L g1495 ( .A(n_1259), .Y(n_1495) );
NOR2xp33_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1263), .Y(n_1260) );
AND4x1_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1283), .C(n_1285), .D(n_1302), .Y(n_1265) );
OAI21xp33_ASAP7_75t_SL g1289 ( .A1(n_1274), .A2(n_1290), .B(n_1291), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1304), .Y(n_1302) );
OAI22x1_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B1(n_1351), .B2(n_1352), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1309), .Y(n_1350) );
NAND3xp33_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1315), .C(n_1318), .Y(n_1310) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
NAND4xp25_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1337), .C(n_1342), .D(n_1345), .Y(n_1332) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1347), .C(n_1348), .Y(n_1345) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx2_ASAP7_75t_SL g1351 ( .A(n_1352), .Y(n_1351) );
INVx2_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
NAND4xp75_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1369), .C(n_1388), .D(n_1390), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1366), .Y(n_1355) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1374), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx2_ASAP7_75t_L g1436 ( .A(n_1394), .Y(n_1436) );
XOR2x2_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1434), .Y(n_1394) );
NOR3xp33_ASAP7_75t_L g1395 ( .A(n_1396), .B(n_1398), .C(n_1418), .Y(n_1395) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1417), .Y(n_1480) );
NAND4xp25_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1425), .C(n_1428), .D(n_1431), .Y(n_1418) );
INVx1_ASAP7_75t_SL g1676 ( .A(n_1437), .Y(n_1676) );
XNOR2xp5_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1581), .Y(n_1437) );
XOR2xp5_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1489), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
AND4x1_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1461), .C(n_1463), .D(n_1486), .Y(n_1441) );
NOR3xp33_ASAP7_75t_SL g1442 ( .A(n_1443), .B(n_1444), .C(n_1459), .Y(n_1442) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1544 ( .A1(n_1452), .A2(n_1458), .B1(n_1545), .B2(n_1546), .Y(n_1544) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1953 ( .A1(n_1467), .A2(n_1954), .B1(n_1955), .B2(n_1957), .Y(n_1953) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx2_ASAP7_75t_L g1476 ( .A(n_1468), .Y(n_1476) );
INVx2_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
OAI221xp5_ASAP7_75t_L g1475 ( .A1(n_1476), .A2(n_1477), .B1(n_1478), .B2(n_1481), .C(n_1482), .Y(n_1475) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
NOR2xp33_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1488), .Y(n_1486) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_1490), .A2(n_1537), .B1(n_1538), .B2(n_1580), .Y(n_1489) );
INVx2_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
HB1xp67_ASAP7_75t_L g1580 ( .A(n_1491), .Y(n_1580) );
XNOR2x1_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1516), .Y(n_1493) );
NAND3xp33_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1504), .C(n_1512), .Y(n_1496) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
NOR3xp33_ASAP7_75t_SL g1516 ( .A(n_1517), .B(n_1524), .C(n_1525), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1521), .Y(n_1517) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
AND4x1_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1557), .C(n_1559), .D(n_1577), .Y(n_1541) );
OAI22xp5_ASAP7_75t_SL g1570 ( .A1(n_1563), .A2(n_1571), .B1(n_1572), .B2(n_1573), .Y(n_1570) );
NOR2xp33_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1579), .Y(n_1577) );
HB1xp67_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
AOI22xp5_ASAP7_75t_L g1582 ( .A1(n_1583), .A2(n_1584), .B1(n_1626), .B2(n_1627), .Y(n_1582) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
NAND4xp75_ASAP7_75t_SL g1585 ( .A(n_1586), .B(n_1594), .C(n_1596), .D(n_1615), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1590), .Y(n_1586) );
OAI22xp5_ASAP7_75t_L g1608 ( .A1(n_1591), .A2(n_1609), .B1(n_1610), .B2(n_1612), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
XNOR2xp5_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
NOR4xp75_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1651), .C(n_1658), .D(n_1660), .Y(n_1629) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1655), .Y(n_1651) );
AOI33xp33_ASAP7_75t_L g1665 ( .A1(n_1666), .A2(n_1667), .A3(n_1668), .B1(n_1673), .B2(n_1674), .B3(n_1675), .Y(n_1665) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
OAI221xp5_ASAP7_75t_L g1677 ( .A1(n_1678), .A2(n_1928), .B1(n_1930), .B2(n_1979), .C(n_1984), .Y(n_1677) );
O2A1O1Ixp33_ASAP7_75t_L g1678 ( .A1(n_1679), .A2(n_1810), .B(n_1846), .C(n_1896), .Y(n_1678) );
NAND5xp2_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1767), .C(n_1795), .D(n_1804), .E(n_1808), .Y(n_1679) );
AOI221xp5_ASAP7_75t_L g1680 ( .A1(n_1681), .A2(n_1717), .B1(n_1742), .B2(n_1749), .C(n_1756), .Y(n_1680) );
INVxp67_ASAP7_75t_SL g1681 ( .A(n_1682), .Y(n_1681) );
NOR2xp33_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1707), .Y(n_1682) );
AOI221xp5_ASAP7_75t_L g1897 ( .A1(n_1683), .A2(n_1724), .B1(n_1831), .B2(n_1898), .C(n_1899), .Y(n_1897) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1703), .Y(n_1683) );
INVx2_ASAP7_75t_L g1710 ( .A(n_1684), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1684), .B(n_1748), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1762 ( .A(n_1684), .B(n_1711), .Y(n_1762) );
OR2x2_ASAP7_75t_L g1798 ( .A(n_1684), .B(n_1711), .Y(n_1798) );
NOR2xp33_ASAP7_75t_L g1852 ( .A(n_1684), .B(n_1703), .Y(n_1852) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1697), .Y(n_1684) );
AND2x4_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1692), .Y(n_1686) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
OR2x2_ASAP7_75t_L g1714 ( .A(n_1688), .B(n_1693), .Y(n_1714) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1691), .Y(n_1688) );
HB1xp67_ASAP7_75t_L g2044 ( .A(n_1689), .Y(n_2044) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1691), .Y(n_1701) );
AND2x4_ASAP7_75t_L g1694 ( .A(n_1692), .B(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1693), .B(n_1696), .Y(n_1716) );
BUFx2_ASAP7_75t_L g1753 ( .A(n_1694), .Y(n_1753) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
AND2x4_ASAP7_75t_L g1702 ( .A(n_1699), .B(n_1701), .Y(n_1702) );
AND2x4_ASAP7_75t_L g1723 ( .A(n_1699), .B(n_1700), .Y(n_1723) );
HB1xp67_ASAP7_75t_L g2042 ( .A(n_1700), .Y(n_2042) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
INVx2_ASAP7_75t_L g1736 ( .A(n_1702), .Y(n_1736) );
OR2x2_ASAP7_75t_L g1761 ( .A(n_1703), .B(n_1720), .Y(n_1761) );
OR2x2_ASAP7_75t_L g1771 ( .A(n_1703), .B(n_1772), .Y(n_1771) );
NAND2xp5_ASAP7_75t_L g1773 ( .A(n_1703), .B(n_1710), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1703), .B(n_1747), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1858 ( .A(n_1703), .B(n_1859), .Y(n_1858) );
OAI322xp33_ASAP7_75t_L g1868 ( .A1(n_1703), .A2(n_1854), .A3(n_1869), .B1(n_1870), .B2(n_1871), .C1(n_1872), .C2(n_1874), .Y(n_1868) );
AND2x2_ASAP7_75t_L g1873 ( .A(n_1703), .B(n_1748), .Y(n_1873) );
BUFx3_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVxp67_ASAP7_75t_L g1708 ( .A(n_1704), .Y(n_1708) );
BUFx2_ASAP7_75t_L g1778 ( .A(n_1704), .Y(n_1778) );
OR2x2_ASAP7_75t_L g1815 ( .A(n_1704), .B(n_1711), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1824 ( .A(n_1704), .B(n_1825), .Y(n_1824) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1706), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_1707), .B(n_1783), .Y(n_1807) );
NAND2xp5_ASAP7_75t_L g1832 ( .A(n_1707), .B(n_1720), .Y(n_1832) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1709), .Y(n_1707) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1708), .B(n_1747), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1708), .B(n_1797), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1910 ( .A(n_1708), .B(n_1830), .Y(n_1910) );
AND2x2_ASAP7_75t_L g1924 ( .A(n_1708), .B(n_1825), .Y(n_1924) );
AND2x2_ASAP7_75t_L g1764 ( .A(n_1709), .B(n_1719), .Y(n_1764) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1709), .Y(n_1839) );
AND2x2_ASAP7_75t_L g1863 ( .A(n_1709), .B(n_1778), .Y(n_1863) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1711), .Y(n_1709) );
INVx2_ASAP7_75t_SL g1748 ( .A(n_1711), .Y(n_1748) );
OAI22xp5_ASAP7_75t_L g1712 ( .A1(n_1713), .A2(n_1714), .B1(n_1715), .B2(n_1716), .Y(n_1712) );
BUFx6f_ASAP7_75t_L g1728 ( .A(n_1714), .Y(n_1728) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1716), .Y(n_1731) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1724), .Y(n_1718) );
NOR2xp33_ASAP7_75t_L g1797 ( .A(n_1719), .B(n_1798), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1838 ( .A(n_1719), .B(n_1825), .Y(n_1838) );
AND2x2_ASAP7_75t_L g1859 ( .A(n_1719), .B(n_1762), .Y(n_1859) );
NOR2xp33_ASAP7_75t_L g1912 ( .A(n_1719), .B(n_1785), .Y(n_1912) );
INVx2_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
BUFx2_ASAP7_75t_L g1745 ( .A(n_1720), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1720), .B(n_1778), .Y(n_1777) );
INVx2_ASAP7_75t_L g1784 ( .A(n_1720), .Y(n_1784) );
AND2x2_ASAP7_75t_L g1830 ( .A(n_1720), .B(n_1762), .Y(n_1830) );
NAND2xp5_ASAP7_75t_L g1869 ( .A(n_1720), .B(n_1803), .Y(n_1869) );
NAND2xp5_ASAP7_75t_L g1882 ( .A(n_1720), .B(n_1725), .Y(n_1882) );
AND2x2_ASAP7_75t_L g1891 ( .A(n_1720), .B(n_1806), .Y(n_1891) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1722), .Y(n_1720) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1723), .Y(n_1734) );
BUFx3_ASAP7_75t_L g1789 ( .A(n_1723), .Y(n_1789) );
AND2x2_ASAP7_75t_L g1799 ( .A(n_1724), .B(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1886 ( .A(n_1724), .Y(n_1886) );
AND2x4_ASAP7_75t_L g1724 ( .A(n_1725), .B(n_1738), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1725), .B(n_1739), .Y(n_1758) );
HB1xp67_ASAP7_75t_L g1775 ( .A(n_1725), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1725), .B(n_1784), .Y(n_1783) );
INVx2_ASAP7_75t_SL g1821 ( .A(n_1725), .Y(n_1821) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1725), .Y(n_1841) );
NAND2xp5_ASAP7_75t_L g1867 ( .A(n_1725), .B(n_1800), .Y(n_1867) );
NOR2xp33_ASAP7_75t_L g1878 ( .A(n_1725), .B(n_1784), .Y(n_1878) );
CKINVDCx5p33_ASAP7_75t_R g1725 ( .A(n_1726), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_1726), .B(n_1738), .Y(n_1803) );
AND2x2_ASAP7_75t_L g1888 ( .A(n_1726), .B(n_1739), .Y(n_1888) );
OR2x2_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1733), .Y(n_1726) );
OAI22xp5_ASAP7_75t_L g1727 ( .A1(n_1728), .A2(n_1729), .B1(n_1730), .B2(n_1732), .Y(n_1727) );
BUFx3_ASAP7_75t_L g1792 ( .A(n_1728), .Y(n_1792) );
HB1xp67_ASAP7_75t_L g1794 ( .A(n_1730), .Y(n_1794) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
OAI22xp5_ASAP7_75t_L g1733 ( .A1(n_1734), .A2(n_1735), .B1(n_1736), .B2(n_1737), .Y(n_1733) );
INVx2_ASAP7_75t_L g1755 ( .A(n_1736), .Y(n_1755) );
INVx1_ASAP7_75t_L g1929 ( .A(n_1736), .Y(n_1929) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1738), .B(n_1751), .Y(n_1766) );
OR2x2_ASAP7_75t_L g1780 ( .A(n_1738), .B(n_1781), .Y(n_1780) );
AOI22xp5_ASAP7_75t_L g1812 ( .A1(n_1738), .A2(n_1813), .B1(n_1814), .B2(n_1816), .Y(n_1812) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1738), .Y(n_1827) );
NAND3xp33_ASAP7_75t_L g1877 ( .A(n_1738), .B(n_1825), .C(n_1878), .Y(n_1877) );
NOR2xp33_ASAP7_75t_L g1881 ( .A(n_1738), .B(n_1882), .Y(n_1881) );
INVx3_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1739), .B(n_1750), .Y(n_1749) );
OR2x2_ASAP7_75t_L g1822 ( .A(n_1739), .B(n_1751), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1740), .B(n_1741), .Y(n_1739) );
AOI211xp5_ASAP7_75t_L g1901 ( .A1(n_1742), .A2(n_1758), .B(n_1902), .C(n_1913), .Y(n_1901) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
OR2x2_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1746), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1744), .B(n_1749), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1851 ( .A(n_1744), .B(n_1852), .Y(n_1851) );
NAND2xp5_ASAP7_75t_L g1862 ( .A(n_1744), .B(n_1863), .Y(n_1862) );
OAI21xp33_ASAP7_75t_L g1925 ( .A1(n_1744), .A2(n_1839), .B(n_1926), .Y(n_1925) );
INVx2_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1894 ( .A(n_1745), .B(n_1747), .Y(n_1894) );
NAND2xp5_ASAP7_75t_L g1906 ( .A(n_1745), .B(n_1827), .Y(n_1906) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1747), .Y(n_1885) );
NOR2x1_ASAP7_75t_L g1921 ( .A(n_1748), .B(n_1778), .Y(n_1921) );
NAND2xp5_ASAP7_75t_L g1840 ( .A(n_1749), .B(n_1841), .Y(n_1840) );
AOI22xp5_ASAP7_75t_L g1857 ( .A1(n_1749), .A2(n_1807), .B1(n_1827), .B2(n_1858), .Y(n_1857) );
AOI322xp5_ASAP7_75t_L g1922 ( .A1(n_1749), .A2(n_1814), .A3(n_1849), .B1(n_1923), .B2(n_1924), .C1(n_1925), .C2(n_1927), .Y(n_1922) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1750), .Y(n_1800) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1750), .Y(n_1811) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1751), .Y(n_1781) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1751), .Y(n_1806) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1752), .B(n_1754), .Y(n_1751) );
OAI22xp5_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1759), .B1(n_1763), .B2(n_1765), .Y(n_1756) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1762), .Y(n_1759) );
OAI211xp5_ASAP7_75t_SL g1916 ( .A1(n_1760), .A2(n_1859), .B(n_1917), .C(n_1920), .Y(n_1916) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
OR2x2_ASAP7_75t_L g1865 ( .A(n_1761), .B(n_1798), .Y(n_1865) );
OR2x2_ASAP7_75t_L g1884 ( .A(n_1761), .B(n_1885), .Y(n_1884) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1762), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1776 ( .A(n_1762), .B(n_1777), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1762), .B(n_1778), .Y(n_1816) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
OAI21xp33_ASAP7_75t_L g1911 ( .A1(n_1764), .A2(n_1799), .B(n_1912), .Y(n_1911) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_1765), .B(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
AOI221xp5_ASAP7_75t_L g1847 ( .A1(n_1766), .A2(n_1848), .B1(n_1849), .B2(n_1850), .C(n_1853), .Y(n_1847) );
NAND2xp5_ASAP7_75t_L g1871 ( .A(n_1766), .B(n_1841), .Y(n_1871) );
AOI211xp5_ASAP7_75t_SL g1767 ( .A1(n_1768), .A2(n_1770), .B(n_1774), .C(n_1779), .Y(n_1767) );
INVxp67_ASAP7_75t_SL g1768 ( .A(n_1769), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1770 ( .A(n_1771), .B(n_1773), .Y(n_1770) );
INVx1_ASAP7_75t_L g1848 ( .A(n_1771), .Y(n_1848) );
NOR2xp33_ASAP7_75t_L g1801 ( .A(n_1773), .B(n_1802), .Y(n_1801) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1773), .Y(n_1904) );
NOR2xp33_ASAP7_75t_L g1774 ( .A(n_1775), .B(n_1776), .Y(n_1774) );
A2O1A1Ixp33_ASAP7_75t_L g1914 ( .A1(n_1775), .A2(n_1830), .B(n_1864), .C(n_1915), .Y(n_1914) );
NAND2xp5_ASAP7_75t_L g1828 ( .A(n_1776), .B(n_1829), .Y(n_1828) );
AND2x2_ASAP7_75t_L g1908 ( .A(n_1777), .B(n_1825), .Y(n_1908) );
AOI321xp33_ASAP7_75t_L g1889 ( .A1(n_1778), .A2(n_1890), .A3(n_1891), .B1(n_1892), .B2(n_1893), .C(n_1895), .Y(n_1889) );
A2O1A1Ixp33_ASAP7_75t_L g1779 ( .A1(n_1780), .A2(n_1782), .B(n_1785), .C(n_1787), .Y(n_1779) );
INVx1_ASAP7_75t_L g1915 ( .A(n_1780), .Y(n_1915) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1784), .B(n_1803), .Y(n_1802) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
INVx3_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVx3_ASAP7_75t_L g1895 ( .A(n_1788), .Y(n_1895) );
OAI22xp33_ASAP7_75t_L g1790 ( .A1(n_1791), .A2(n_1792), .B1(n_1793), .B2(n_1794), .Y(n_1790) );
AOI21xp5_ASAP7_75t_L g1795 ( .A1(n_1796), .A2(n_1799), .B(n_1801), .Y(n_1795) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1797), .Y(n_1874) );
NOR2xp33_ASAP7_75t_L g1809 ( .A(n_1798), .B(n_1802), .Y(n_1809) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1798), .Y(n_1825) );
AND2x2_ASAP7_75t_L g1855 ( .A(n_1800), .B(n_1841), .Y(n_1855) );
INVx2_ASAP7_75t_L g1870 ( .A(n_1800), .Y(n_1870) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1802), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1803), .B(n_1806), .Y(n_1849) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1805), .B(n_1807), .Y(n_1804) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
NAND2xp5_ASAP7_75t_L g1835 ( .A(n_1806), .B(n_1836), .Y(n_1835) );
INVxp67_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
OAI211xp5_ASAP7_75t_L g1810 ( .A1(n_1811), .A2(n_1812), .B(n_1817), .C(n_1842), .Y(n_1810) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1811), .Y(n_1833) );
OAI211xp5_ASAP7_75t_SL g1896 ( .A1(n_1811), .A2(n_1897), .B(n_1901), .C(n_1922), .Y(n_1896) );
INVx1_ASAP7_75t_L g1919 ( .A(n_1811), .Y(n_1919) );
NAND2xp5_ASAP7_75t_L g1880 ( .A(n_1814), .B(n_1881), .Y(n_1880) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1816), .Y(n_1900) );
AOI221xp5_ASAP7_75t_L g1817 ( .A1(n_1818), .A2(n_1830), .B1(n_1831), .B2(n_1833), .C(n_1834), .Y(n_1817) );
NAND3xp33_ASAP7_75t_L g1818 ( .A(n_1819), .B(n_1823), .C(n_1826), .Y(n_1818) );
INVx1_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
NOR2xp33_ASAP7_75t_L g1820 ( .A(n_1821), .B(n_1822), .Y(n_1820) );
INVx2_ASAP7_75t_L g1829 ( .A(n_1821), .Y(n_1829) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1821), .Y(n_1836) );
AND2x2_ASAP7_75t_L g1907 ( .A(n_1821), .B(n_1908), .Y(n_1907) );
INVxp67_ASAP7_75t_L g1844 ( .A(n_1823), .Y(n_1844) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1824), .Y(n_1856) );
INVxp67_ASAP7_75t_L g1843 ( .A(n_1826), .Y(n_1843) );
NAND2xp5_ASAP7_75t_L g1826 ( .A(n_1827), .B(n_1828), .Y(n_1826) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
OAI22xp5_ASAP7_75t_L g1834 ( .A1(n_1835), .A2(n_1837), .B1(n_1839), .B2(n_1840), .Y(n_1834) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1835), .Y(n_1892) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
NAND2xp5_ASAP7_75t_L g1890 ( .A(n_1839), .B(n_1885), .Y(n_1890) );
INVx1_ASAP7_75t_L g1927 ( .A(n_1840), .Y(n_1927) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1841), .Y(n_1845) );
OAI21xp5_ASAP7_75t_L g1842 ( .A1(n_1843), .A2(n_1844), .B(n_1845), .Y(n_1842) );
NAND5xp2_ASAP7_75t_L g1846 ( .A(n_1847), .B(n_1857), .C(n_1860), .D(n_1875), .E(n_1889), .Y(n_1846) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
NOR2xp33_ASAP7_75t_L g1853 ( .A(n_1854), .B(n_1856), .Y(n_1853) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
O2A1O1Ixp33_ASAP7_75t_L g1860 ( .A1(n_1861), .A2(n_1864), .B(n_1866), .C(n_1868), .Y(n_1860) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
INVx1_ASAP7_75t_L g1926 ( .A(n_1863), .Y(n_1926) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
OAI22xp33_ASAP7_75t_L g1883 ( .A1(n_1865), .A2(n_1884), .B1(n_1886), .B2(n_1887), .Y(n_1883) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1898 ( .A(n_1869), .Y(n_1898) );
OAI221xp5_ASAP7_75t_L g1902 ( .A1(n_1870), .A2(n_1871), .B1(n_1903), .B2(n_1909), .C(n_1911), .Y(n_1902) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
NOR3xp33_ASAP7_75t_SL g1875 ( .A(n_1876), .B(n_1879), .C(n_1883), .Y(n_1875) );
INVxp67_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
INVxp67_ASAP7_75t_SL g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1923 ( .A(n_1882), .Y(n_1923) );
NOR2xp33_ASAP7_75t_L g1899 ( .A(n_1886), .B(n_1900), .Y(n_1899) );
OR2x2_ASAP7_75t_L g1918 ( .A(n_1887), .B(n_1919), .Y(n_1918) );
CKINVDCx5p33_ASAP7_75t_R g1887 ( .A(n_1888), .Y(n_1887) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1894), .Y(n_1893) );
AOI21xp33_ASAP7_75t_L g1903 ( .A1(n_1904), .A2(n_1905), .B(n_1907), .Y(n_1903) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1906), .Y(n_1905) );
INVx1_ASAP7_75t_L g1909 ( .A(n_1910), .Y(n_1909) );
NAND2xp5_ASAP7_75t_SL g1913 ( .A(n_1914), .B(n_1916), .Y(n_1913) );
INVx1_ASAP7_75t_L g1917 ( .A(n_1918), .Y(n_1917) );
INVx1_ASAP7_75t_L g1920 ( .A(n_1921), .Y(n_1920) );
INVx1_ASAP7_75t_L g1928 ( .A(n_1929), .Y(n_1928) );
AND2x2_ASAP7_75t_L g1931 ( .A(n_1932), .B(n_1961), .Y(n_1931) );
NOR3xp33_ASAP7_75t_SL g1932 ( .A(n_1933), .B(n_1942), .C(n_1944), .Y(n_1932) );
NAND2xp5_ASAP7_75t_L g1933 ( .A(n_1934), .B(n_1938), .Y(n_1933) );
OAI211xp5_ASAP7_75t_L g1968 ( .A1(n_1937), .A2(n_1969), .B(n_1970), .C(n_1971), .Y(n_1968) );
INVx3_ASAP7_75t_L g1946 ( .A(n_1947), .Y(n_1946) );
INVx1_ASAP7_75t_L g1955 ( .A(n_1956), .Y(n_1955) );
INVx1_ASAP7_75t_SL g1966 ( .A(n_1967), .Y(n_1966) );
INVx1_ASAP7_75t_L g1975 ( .A(n_1976), .Y(n_1975) );
CKINVDCx14_ASAP7_75t_R g1979 ( .A(n_1980), .Y(n_1979) );
INVx2_ASAP7_75t_L g1980 ( .A(n_1981), .Y(n_1980) );
CKINVDCx5p33_ASAP7_75t_R g1981 ( .A(n_1982), .Y(n_1981) );
A2O1A1Ixp33_ASAP7_75t_L g2040 ( .A1(n_1983), .A2(n_2041), .B(n_2043), .C(n_2045), .Y(n_2040) );
BUFx2_ASAP7_75t_L g1985 ( .A(n_1986), .Y(n_1985) );
INVx1_ASAP7_75t_L g1986 ( .A(n_1987), .Y(n_1986) );
INVx1_ASAP7_75t_L g1987 ( .A(n_1988), .Y(n_1987) );
INVx1_ASAP7_75t_L g1989 ( .A(n_1990), .Y(n_1989) );
INVx1_ASAP7_75t_L g1990 ( .A(n_1991), .Y(n_1990) );
INVx1_ASAP7_75t_L g1991 ( .A(n_1992), .Y(n_1991) );
OAI21xp5_ASAP7_75t_SL g2010 ( .A1(n_1999), .A2(n_2011), .B(n_2012), .Y(n_2010) );
INVx1_ASAP7_75t_L g2000 ( .A(n_2001), .Y(n_2000) );
NAND3xp33_ASAP7_75t_L g2007 ( .A(n_2008), .B(n_2019), .C(n_2022), .Y(n_2007) );
NAND2xp5_ASAP7_75t_L g2014 ( .A(n_2015), .B(n_2016), .Y(n_2014) );
INVx2_ASAP7_75t_L g2017 ( .A(n_2018), .Y(n_2017) );
OAI221xp5_ASAP7_75t_L g2034 ( .A1(n_2020), .A2(n_2021), .B1(n_2029), .B2(n_2035), .C(n_2037), .Y(n_2034) );
INVx2_ASAP7_75t_L g2029 ( .A(n_2030), .Y(n_2029) );
INVx1_ASAP7_75t_L g2035 ( .A(n_2036), .Y(n_2035) );
BUFx2_ASAP7_75t_L g2038 ( .A(n_2039), .Y(n_2038) );
HB1xp67_ASAP7_75t_L g2039 ( .A(n_2040), .Y(n_2039) );
INVx1_ASAP7_75t_L g2041 ( .A(n_2042), .Y(n_2041) );
INVx1_ASAP7_75t_L g2043 ( .A(n_2044), .Y(n_2043) );
endmodule