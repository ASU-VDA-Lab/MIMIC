module fake_aes_7526_n_730 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_730);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_730;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g80 ( .A(n_20), .B(n_46), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_41), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_71), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_66), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_77), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_7), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_44), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_9), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_6), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_12), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_16), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_74), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_15), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_7), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_55), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
BUFx10_ASAP7_75t_L g100 ( .A(n_26), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_31), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_54), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_53), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_3), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_9), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_68), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_64), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_57), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_52), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_39), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_72), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_78), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_30), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_17), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_67), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_75), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_21), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_32), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_8), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_48), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_10), .B(n_15), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_65), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_122), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_109), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_125), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_122), .B(n_0), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_81), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_97), .B(n_1), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_102), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_96), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_86), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
NOR2x1_ASAP7_75t_L g144 ( .A(n_118), .B(n_42), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_117), .B(n_4), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVxp33_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_81), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_104), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_95), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_118), .B(n_5), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_113), .B(n_5), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_113), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_98), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_89), .B(n_10), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_82), .B(n_11), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_89), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_98), .Y(n_166) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_110), .B(n_79), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_101), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_112), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_112), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_90), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_130), .B(n_119), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_130), .B(n_103), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_157), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_131), .B(n_99), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_138), .Y(n_183) );
OR2x6_ASAP7_75t_L g184 ( .A(n_136), .B(n_115), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_161), .B(n_90), .Y(n_185) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_167), .B(n_128), .Y(n_186) );
NOR2xp33_ASAP7_75t_SL g187 ( .A(n_138), .B(n_103), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_148), .B(n_123), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_152), .B(n_120), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
BUFx10_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_135), .B(n_123), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_135), .B(n_101), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_151), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_161), .A2(n_120), .B1(n_91), .B2(n_93), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
BUFx10_ASAP7_75t_L g203 ( .A(n_169), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_140), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_169), .B(n_100), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_129), .Y(n_207) );
BUFx10_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_143), .B(n_126), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_140), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_154), .B(n_100), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_167), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_165), .B(n_100), .Y(n_214) );
INVx6_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_129), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_143), .B(n_87), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_145), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_145), .B(n_126), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_153), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_150), .B(n_107), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_150), .B(n_106), .Y(n_225) );
INVxp67_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_162), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_171), .B(n_91), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_134), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_134), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_155), .Y(n_231) );
NAND2xp33_ASAP7_75t_R g232 ( .A(n_146), .B(n_93), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_142), .B(n_115), .Y(n_234) );
BUFx10_ASAP7_75t_L g235 ( .A(n_155), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_156), .A2(n_127), .B1(n_128), .B2(n_124), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_156), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_147), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_237), .A2(n_170), .B(n_168), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_188), .B(n_171), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_184), .B(n_132), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_218), .B(n_170), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_184), .B(n_168), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_182), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_195), .B(n_206), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_235), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_194), .B(n_166), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_235), .Y(n_248) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_184), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_235), .B(n_166), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_231), .B(n_160), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_199), .B(n_160), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_230), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_210), .B(n_164), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_179), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_226), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_230), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_222), .B(n_158), .C(n_124), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_228), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_195), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_175), .A2(n_163), .B(n_159), .C(n_149), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_221), .B(n_141), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_198), .Y(n_267) );
AND3x1_ASAP7_75t_L g268 ( .A(n_187), .B(n_144), .C(n_141), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_179), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_213), .B(n_141), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_212), .B(n_163), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_229), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_186), .A2(n_159), .B1(n_149), .B2(n_116), .Y(n_273) );
NAND2x1p5_ASAP7_75t_L g274 ( .A(n_206), .B(n_114), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_184), .B(n_108), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_176), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_191), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_231), .B(n_84), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_212), .B(n_83), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_182), .B(n_80), .Y(n_280) );
AOI22xp33_ASAP7_75t_SL g281 ( .A1(n_213), .A2(n_105), .B1(n_12), .B2(n_13), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_183), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_200), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_186), .A2(n_11), .B1(n_14), .B2(n_16), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_177), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_214), .B(n_17), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_185), .B(n_18), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_191), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_178), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_185), .B(n_23), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_209), .B(n_25), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_182), .B(n_27), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_213), .A2(n_28), .B1(n_35), .B2(n_36), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_181), .B(n_38), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_220), .B(n_40), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_196), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_185), .B(n_43), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_190), .B(n_45), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_178), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_201), .B(n_47), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_193), .B(n_49), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_197), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_192), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_174), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_208), .A2(n_50), .B1(n_51), .B2(n_56), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_207), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_243), .B(n_173), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_243), .B(n_178), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_243), .B(n_298), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_283), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_246), .B(n_208), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_253), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_307), .B(n_208), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_282), .B(n_203), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_291), .B(n_205), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_279), .B(n_222), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_302), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_246), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
OAI22xp5_ASAP7_75t_SL g325 ( .A1(n_259), .A2(n_234), .B1(n_236), .B2(n_203), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_259), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_263), .B(n_203), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_245), .B(n_193), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_240), .B(n_193), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_270), .B(n_234), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_241), .A2(n_232), .B1(n_234), .B2(n_225), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_270), .B(n_234), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_262), .A2(n_207), .B1(n_217), .B2(n_238), .Y(n_334) );
AO22x1_ASAP7_75t_L g335 ( .A1(n_241), .A2(n_207), .B1(n_217), .B2(n_233), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_271), .B(n_223), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_263), .B(n_217), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
AOI21xp33_ASAP7_75t_L g339 ( .A1(n_286), .A2(n_238), .B(n_233), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_239), .A2(n_189), .B(n_180), .C(n_216), .Y(n_340) );
INVx6_ASAP7_75t_SL g341 ( .A(n_270), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_264), .A2(n_189), .B(n_180), .C(n_216), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_274), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_245), .B(n_219), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_275), .B(n_219), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_289), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_276), .Y(n_347) );
NOR2x1_ASAP7_75t_R g348 ( .A(n_241), .B(n_219), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_285), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_250), .A2(n_204), .B(n_202), .Y(n_350) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_249), .B(n_227), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_289), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_242), .A2(n_227), .B1(n_204), .B2(n_211), .C(n_202), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_249), .A2(n_215), .B1(n_211), .B2(n_197), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_287), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_266), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_274), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_272), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_306), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_249), .Y(n_360) );
BUFx12f_ASAP7_75t_L g361 ( .A(n_270), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_275), .B(n_215), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_265), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_255), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_312), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_314), .B(n_248), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_355), .A2(n_287), .B1(n_290), .B2(n_273), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_361), .B(n_290), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_327), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_355), .A2(n_290), .B1(n_301), .B2(n_275), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_294), .B(n_297), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_356), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_SL g373 ( .A1(n_342), .A2(n_294), .B(n_264), .C(n_296), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_356), .A2(n_300), .B(n_295), .Y(n_374) );
NOR2xp33_ASAP7_75t_R g375 ( .A(n_327), .B(n_304), .Y(n_375) );
INVx3_ASAP7_75t_SL g376 ( .A(n_323), .Y(n_376) );
BUFx12f_ASAP7_75t_L g377 ( .A(n_361), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_358), .A2(n_308), .B(n_268), .Y(n_378) );
O2A1O1Ixp5_ASAP7_75t_L g379 ( .A1(n_335), .A2(n_280), .B(n_304), .C(n_293), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_358), .A2(n_280), .B(n_278), .Y(n_380) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_342), .A2(n_278), .B(n_301), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_354), .A2(n_303), .B(n_251), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_357), .B(n_244), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_337), .A2(n_251), .B(n_247), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_355), .A2(n_284), .B1(n_254), .B2(n_260), .Y(n_385) );
BUFx4f_ASAP7_75t_SL g386 ( .A(n_341), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_321), .B(n_257), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
OAI21x1_ASAP7_75t_SL g389 ( .A1(n_357), .A2(n_309), .B(n_305), .Y(n_389) );
INVx4_ASAP7_75t_SL g390 ( .A(n_324), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_340), .A2(n_224), .B(n_250), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_332), .A2(n_261), .B1(n_281), .B2(n_244), .C(n_260), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_315), .A2(n_224), .B(n_305), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_336), .B(n_255), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_331), .B(n_244), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_320), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_330), .A2(n_299), .B(n_292), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_387), .B(n_313), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_370), .A2(n_348), .B(n_328), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_373), .A2(n_367), .B(n_340), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_339), .B(n_353), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_372), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_343), .B1(n_324), .B2(n_360), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_395), .B(n_363), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_377), .Y(n_408) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_359), .B(n_349), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_375), .A2(n_319), .B(n_318), .C(n_310), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_368), .A2(n_324), .B1(n_360), .B2(n_317), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_397), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_394), .A2(n_347), .B(n_334), .Y(n_413) );
AO31x2_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_326), .A3(n_316), .B(n_322), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_396), .B(n_331), .Y(n_415) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_368), .B(n_324), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_368), .A2(n_333), .B1(n_331), .B2(n_325), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_392), .A2(n_333), .B1(n_319), .B2(n_328), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_369), .A2(n_334), .B1(n_311), .B2(n_329), .C(n_345), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_376), .A2(n_333), .B1(n_323), .B2(n_364), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_397), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_376), .B(n_344), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_396), .A2(n_320), .B1(n_338), .B2(n_322), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_338), .B1(n_352), .B2(n_346), .Y(n_425) );
OAI22xp33_ASAP7_75t_SL g426 ( .A1(n_388), .A2(n_351), .B1(n_315), .B2(n_346), .Y(n_426) );
AO21x1_ASAP7_75t_SL g427 ( .A1(n_390), .A2(n_362), .B(n_323), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_409), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_403), .B(n_390), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_403), .B(n_381), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_404), .B(n_381), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_404), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_421), .B(n_390), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_421), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_409), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_412), .B(n_390), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_412), .B(n_323), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_427), .Y(n_440) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_401), .A2(n_389), .B(n_378), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_408), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_422), .B(n_381), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_422), .B(n_376), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_407), .B(n_380), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_424), .B(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_414), .B(n_383), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_414), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_414), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_406), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_378), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_416), .B(n_383), .Y(n_458) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_405), .B(n_388), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_414), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_418), .B(n_384), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_416), .B(n_383), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_384), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_417), .B(n_391), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_444), .B(n_402), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_444), .B(n_402), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_445), .B(n_410), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_430), .B(n_402), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_443), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_430), .B(n_402), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_428), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_433), .B(n_419), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_455), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_440), .B(n_391), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_440), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_440), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_456), .A2(n_411), .B1(n_400), .B2(n_415), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_428), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g481 ( .A(n_429), .B(n_393), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_443), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_427), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_431), .B(n_391), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_433), .B(n_423), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_432), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_435), .B(n_425), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_440), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_455), .A2(n_393), .B1(n_366), .B2(n_379), .C(n_420), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_440), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_435), .B(n_382), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_439), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_439), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_456), .A2(n_426), .B1(n_389), .B2(n_398), .C(n_198), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_432), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
AOI211xp5_ASAP7_75t_L g497 ( .A1(n_458), .A2(n_386), .B(n_377), .C(n_352), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_463), .B(n_382), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_463), .B(n_58), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_436), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_436), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_464), .B(n_352), .Y(n_503) );
XNOR2x2_ASAP7_75t_L g504 ( .A(n_459), .B(n_371), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_451), .Y(n_505) );
OAI31xp33_ASAP7_75t_L g506 ( .A1(n_449), .A2(n_346), .A3(n_269), .B(n_288), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_451), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_446), .B(n_59), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_446), .B(n_60), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_459), .B(n_198), .C(n_252), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_464), .B(n_371), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_449), .B(n_198), .Y(n_513) );
INVx4_ASAP7_75t_L g514 ( .A(n_440), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_453), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_461), .B(n_252), .C(n_267), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_490), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_474), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_465), .B(n_449), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_514), .B(n_434), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_465), .B(n_449), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_468), .B(n_462), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_506), .A2(n_460), .B(n_452), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_466), .B(n_453), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_470), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_474), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_472), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_466), .B(n_452), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_467), .B(n_461), .C(n_462), .D(n_458), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_483), .B(n_460), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_498), .B(n_453), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_483), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_514), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_490), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_487), .B(n_429), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_476), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_498), .B(n_457), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_492), .B(n_457), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_484), .B(n_454), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_484), .B(n_454), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_482), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_482), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_472), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_469), .B(n_450), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_469), .B(n_450), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_487), .A2(n_429), .B1(n_434), .B2(n_441), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_493), .B(n_448), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_481), .B(n_442), .Y(n_551) );
AOI211x1_ASAP7_75t_L g552 ( .A1(n_489), .A2(n_448), .B(n_434), .C(n_429), .Y(n_552) );
NAND3x1_ASAP7_75t_L g553 ( .A(n_506), .B(n_434), .C(n_437), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_479), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_485), .B(n_437), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_485), .B(n_437), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_493), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_471), .B(n_447), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_514), .B(n_447), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_473), .B(n_437), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_471), .B(n_447), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_514), .B(n_447), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_495), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_476), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_491), .B(n_441), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_478), .A2(n_441), .B1(n_438), .B2(n_215), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_505), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_491), .B(n_441), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_476), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_477), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_438), .Y(n_571) );
OR3x1_ASAP7_75t_L g572 ( .A(n_504), .B(n_438), .C(n_62), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_507), .B(n_438), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_479), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_479), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_503), .B(n_61), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_507), .B(n_63), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_525), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_558), .B(n_475), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_528), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_558), .B(n_475), .Y(n_581) );
NAND4xp25_ASAP7_75t_L g582 ( .A(n_552), .B(n_497), .C(n_478), .D(n_473), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_531), .A2(n_510), .B1(n_481), .B2(n_477), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_561), .B(n_475), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_535), .B(n_488), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_534), .B(n_495), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_530), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_532), .B(n_502), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_535), .B(n_488), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_526), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_561), .B(n_475), .Y(n_594) );
NAND2x1_ASAP7_75t_L g595 ( .A(n_535), .B(n_510), .Y(n_595) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_572), .B(n_488), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_531), .B(n_481), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_535), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_532), .B(n_496), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_543), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_543), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_519), .B(n_477), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_519), .B(n_499), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_529), .B(n_518), .Y(n_605) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_563), .Y(n_606) );
INVxp33_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
AND2x4_ASAP7_75t_SL g608 ( .A(n_538), .B(n_499), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_527), .B(n_496), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_529), .B(n_502), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_546), .B(n_515), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_521), .B(n_503), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_521), .B(n_508), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_544), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_524), .B(n_512), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_527), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_524), .B(n_533), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_545), .Y(n_618) );
AND2x2_ASAP7_75t_SL g619 ( .A(n_559), .B(n_508), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_555), .B(n_480), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_546), .B(n_515), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_533), .B(n_512), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_556), .B(n_480), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_549), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_547), .B(n_512), .Y(n_626) );
XOR2xp5_ASAP7_75t_L g627 ( .A(n_522), .B(n_504), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_549), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_551), .Y(n_629) );
NAND2xp33_ASAP7_75t_SL g630 ( .A(n_576), .B(n_509), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_557), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_606), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_597), .A2(n_553), .B1(n_560), .B2(n_537), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_583), .A2(n_553), .B(n_576), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_588), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_597), .A2(n_568), .B1(n_565), .B2(n_557), .C1(n_539), .C2(n_541), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_590), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_608), .A2(n_497), .B(n_523), .C(n_520), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_617), .B(n_547), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_582), .B(n_494), .C(n_513), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_578), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_617), .B(n_541), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_627), .A2(n_548), .B1(n_565), .B2(n_568), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_619), .A2(n_572), .B1(n_552), .B2(n_562), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_608), .A2(n_517), .B(n_564), .C(n_569), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_626), .B(n_542), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_585), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_592), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_598), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_583), .A2(n_513), .B(n_536), .C(n_509), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_593), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_609), .A2(n_566), .B(n_577), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_629), .A2(n_542), .B1(n_539), .B2(n_567), .C(n_566), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_600), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_601), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_605), .B(n_540), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_599), .B(n_540), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_602), .B(n_559), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_615), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_619), .B(n_577), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_598), .B(n_559), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_616), .B(n_564), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_614), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_595), .A2(n_559), .B(n_536), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_630), .A2(n_517), .B1(n_562), .B2(n_564), .C(n_570), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_624), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_609), .B(n_567), .C(n_550), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_596), .A2(n_516), .B(n_571), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_630), .A2(n_569), .B1(n_570), .B2(n_573), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g670 ( .A1(n_638), .A2(n_607), .B(n_591), .Y(n_670) );
INVxp33_ASAP7_75t_SL g671 ( .A(n_644), .Y(n_671) );
AOI31xp33_ASAP7_75t_L g672 ( .A1(n_634), .A2(n_591), .A3(n_607), .B(n_587), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_656), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_643), .A2(n_626), .A3(n_603), .B1(n_579), .B2(n_581), .C1(n_594), .C2(n_586), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g675 ( .A1(n_650), .A2(n_587), .B(n_613), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_636), .B(n_611), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_632), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_639), .B(n_610), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_658), .B(n_594), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_633), .A2(n_621), .B1(n_612), .B2(n_625), .C(n_631), .Y(n_680) );
AOI31xp33_ASAP7_75t_L g681 ( .A1(n_660), .A2(n_587), .A3(n_581), .B(n_586), .Y(n_681) );
OAI31xp33_ASAP7_75t_SL g682 ( .A1(n_665), .A2(n_579), .A3(n_615), .B(n_622), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_640), .A2(n_628), .B(n_570), .C(n_569), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_661), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_641), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_636), .B(n_622), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_647), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_662), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_648), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_635), .B(n_623), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_649), .Y(n_691) );
OA21x2_ASAP7_75t_SL g692 ( .A1(n_649), .A2(n_517), .B(n_620), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_637), .B(n_618), .Y(n_693) );
OAI31xp33_ASAP7_75t_L g694 ( .A1(n_671), .A2(n_660), .A3(n_645), .B(n_667), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_676), .B(n_653), .Y(n_695) );
OAI31xp33_ASAP7_75t_L g696 ( .A1(n_671), .A2(n_667), .A3(n_664), .B(n_661), .Y(n_696) );
OAI22xp5_ASAP7_75t_SL g697 ( .A1(n_688), .A2(n_669), .B1(n_652), .B2(n_668), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g698 ( .A1(n_672), .A2(n_642), .B(n_657), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_670), .A2(n_666), .B1(n_663), .B2(n_651), .Y(n_699) );
AO22x2_ASAP7_75t_L g700 ( .A1(n_692), .A2(n_655), .B1(n_654), .B2(n_659), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_683), .A2(n_550), .B(n_511), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_691), .B(n_571), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_681), .A2(n_646), .B1(n_618), .B2(n_604), .Y(n_703) );
AOI322xp5_ASAP7_75t_L g704 ( .A1(n_686), .A2(n_604), .A3(n_589), .B1(n_584), .B2(n_580), .C1(n_573), .C2(n_574), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_685), .Y(n_705) );
AOI221xp5_ASAP7_75t_SL g706 ( .A1(n_680), .A2(n_589), .B1(n_584), .B2(n_580), .C(n_575), .Y(n_706) );
AO22x2_ASAP7_75t_L g707 ( .A1(n_675), .A2(n_684), .B1(n_677), .B2(n_673), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_689), .B1(n_687), .B2(n_684), .C(n_693), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_694), .A2(n_682), .B(n_688), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g710 ( .A(n_696), .B(n_674), .C(n_684), .D(n_690), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_697), .A2(n_678), .B(n_679), .C(n_511), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_699), .A2(n_575), .B1(n_574), .B2(n_554), .C(n_545), .Y(n_712) );
NOR4xp25_ASAP7_75t_L g713 ( .A(n_695), .B(n_516), .C(n_554), .D(n_501), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_698), .A2(n_500), .B1(n_486), .B2(n_480), .C(n_501), .Y(n_714) );
AOI211xp5_ASAP7_75t_L g715 ( .A1(n_703), .A2(n_501), .B(n_500), .C(n_486), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_708), .B(n_706), .C(n_701), .Y(n_716) );
AND3x4_ASAP7_75t_L g717 ( .A(n_713), .B(n_700), .C(n_704), .Y(n_717) );
NOR3xp33_ASAP7_75t_SL g718 ( .A(n_709), .B(n_710), .C(n_714), .Y(n_718) );
OAI321xp33_ASAP7_75t_L g719 ( .A1(n_711), .A2(n_702), .A3(n_700), .B1(n_705), .B2(n_500), .C(n_486), .Y(n_719) );
AOI211xp5_ASAP7_75t_L g720 ( .A1(n_715), .A2(n_69), .B(n_70), .C(n_73), .Y(n_720) );
OA22x2_ASAP7_75t_L g721 ( .A1(n_717), .A2(n_712), .B1(n_76), .B2(n_277), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g722 ( .A(n_718), .B(n_215), .C(n_269), .D(n_258), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_716), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_723), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_722), .B(n_720), .Y(n_725) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_724), .A2(n_721), .B(n_719), .C(n_288), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_726), .Y(n_727) );
AOI222xp33_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_725), .B1(n_258), .B2(n_277), .C1(n_292), .C2(n_299), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_252), .B1(n_267), .B2(n_723), .Y(n_729) );
OAI221xp5_ASAP7_75t_SL g730 ( .A1(n_729), .A2(n_252), .B1(n_267), .B2(n_723), .C(n_724), .Y(n_730) );
endmodule