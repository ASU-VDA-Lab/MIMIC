module real_jpeg_14753_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_29),
.B1(n_33),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_88),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_68),
.B1(n_70),
.B2(n_88),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_58),
.B1(n_63),
.B2(n_88),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_2),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_2),
.A2(n_29),
.B1(n_33),
.B2(n_136),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_2),
.A2(n_68),
.B1(n_70),
.B2(n_136),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_2),
.A2(n_58),
.B1(n_63),
.B2(n_136),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_29),
.B1(n_33),
.B2(n_172),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_4),
.A2(n_68),
.B1(n_70),
.B2(n_172),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_4),
.A2(n_58),
.B1(n_63),
.B2(n_172),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_5),
.A2(n_29),
.B1(n_33),
.B2(n_80),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_68),
.B1(n_70),
.B2(n_80),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_5),
.A2(n_58),
.B1(n_63),
.B2(n_80),
.Y(n_240)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_58),
.B1(n_63),
.B2(n_67),
.Y(n_163)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_9),
.A2(n_40),
.B1(n_58),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_40),
.B1(n_68),
.B2(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_29),
.B1(n_33),
.B2(n_40),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_82),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_68),
.B1(n_70),
.B2(n_82),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_10),
.A2(n_58),
.B1(n_63),
.B2(n_82),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_12),
.Y(n_341)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_16),
.A2(n_29),
.B1(n_33),
.B2(n_187),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_16),
.A2(n_68),
.B1(n_70),
.B2(n_187),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_16),
.A2(n_58),
.B1(n_63),
.B2(n_187),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B(n_340),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_17),
.B(n_341),
.Y(n_340)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_18),
.A2(n_35),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_18),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_18),
.B(n_38),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_18),
.A2(n_68),
.B1(n_70),
.B2(n_185),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_18),
.A2(n_70),
.B(n_73),
.C(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_18),
.B(n_95),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_18),
.B(n_61),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_18),
.B(n_77),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_18),
.A2(n_33),
.B(n_89),
.C(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_19),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_19),
.A2(n_43),
.B1(n_68),
.B2(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_19),
.A2(n_29),
.B1(n_33),
.B2(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_19),
.A2(n_43),
.B1(n_58),
.B2(n_63),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_38),
.B(n_39),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_26),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_26),
.A2(n_38),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_26),
.A2(n_38),
.B1(n_42),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_27),
.A2(n_28),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_28),
.B1(n_81),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_27),
.A2(n_28),
.B1(n_79),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_27),
.A2(n_28),
.B1(n_101),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_27),
.A2(n_28),
.B1(n_135),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_27),
.A2(n_28),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_29),
.A2(n_33),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_29),
.A2(n_32),
.A3(n_35),
.B1(n_184),
.B2(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_29),
.B(n_185),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_31),
.B(n_33),
.Y(n_202)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g236 ( 
.A1(n_33),
.A2(n_68),
.A3(n_91),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_36),
.B(n_185),
.Y(n_184)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_41),
.B(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_45),
.B(n_339),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_335),
.B(n_337),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_323),
.B(n_334),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_150),
.B(n_320),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_137),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_112),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_51),
.B(n_112),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_83),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_52),
.B(n_98),
.C(n_110),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_78),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_54),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_64),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_56),
.B1(n_78),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_62),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_57),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_57),
.A2(n_61),
.B1(n_163),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_57),
.A2(n_61),
.B1(n_199),
.B2(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_57),
.A2(n_61),
.B1(n_210),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_57),
.A2(n_61),
.B1(n_240),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_57),
.A2(n_61),
.B1(n_185),
.B2(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_57),
.A2(n_61),
.B1(n_266),
.B2(n_273),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_58),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_63),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_58),
.B(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_60),
.A2(n_126),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_60),
.A2(n_161),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_63),
.A2(n_74),
.B(n_185),
.Y(n_254)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_66),
.A2(n_71),
.B1(n_77),
.B2(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_70),
.B1(n_91),
.B2(n_92),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_70),
.B(n_92),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_76),
.B1(n_77),
.B2(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_77),
.B(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_71),
.A2(n_77),
.B1(n_166),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_71),
.A2(n_77),
.B1(n_193),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_71),
.A2(n_77),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_71),
.A2(n_77),
.B1(n_252),
.B2(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_75),
.A2(n_130),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_75),
.A2(n_167),
.B1(n_232),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_98),
.B1(n_110),
.B2(n_111),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_85),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_96),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_87),
.A2(n_93),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_89),
.A2(n_95),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_89),
.A2(n_95),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_89),
.A2(n_95),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_108),
.B1(n_132),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_93),
.A2(n_132),
.B1(n_133),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_93),
.A2(n_132),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_93),
.A2(n_206),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_100),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_104),
.C(n_106),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_100),
.B(n_140),
.C(n_143),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_109),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_104),
.B(n_146),
.C(n_148),
.Y(n_333)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_131),
.C(n_134),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_122),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_306)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_137),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_138),
.B(n_139),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_147),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_149),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_175),
.B(n_319),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_173),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_152),
.B(n_173),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_153),
.B(n_156),
.Y(n_317)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_157),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_168),
.C(n_170),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_158),
.A2(n_159),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_164),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_168),
.B(n_170),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_314),
.B(n_318),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_224),
.B(n_302),
.C(n_313),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_211),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_178),
.B(n_211),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_196),
.C(n_203),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_179),
.A2(n_180),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_189),
.C(n_195),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_196),
.B(n_203),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_213),
.B(n_214),
.C(n_215),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_223),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_217),
.B(n_220),
.C(n_223),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_301),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_244),
.B(n_300),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_241),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_227),
.B(n_241),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_230),
.A2(n_233),
.B1(n_234),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_294),
.B(n_299),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_282),
.B(n_293),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_262),
.B(n_281),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_248),
.B(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_258),
.C(n_260),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_261),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_270),
.B(n_280),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_268),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_279),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_304),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_312),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_325),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_331),
.C(n_333),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);


endmodule