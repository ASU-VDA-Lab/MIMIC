module fake_ariane_2994_n_1995 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1995);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1995;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_363;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_197),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_141),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_85),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_97),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_78),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_45),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_90),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_161),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_149),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_89),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_162),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_104),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_185),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_44),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_188),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_105),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_155),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_76),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_127),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_138),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_9),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_5),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_125),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_25),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_17),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_121),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_189),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_92),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_78),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_165),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_58),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_117),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_103),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_79),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_99),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_114),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_107),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_16),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_10),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_166),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_163),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_170),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_172),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_31),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_25),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_72),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_73),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_45),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_110),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_193),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_94),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_59),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_106),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_19),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_62),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_21),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_57),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_57),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_3),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_144),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_122),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_70),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_175),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_27),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_192),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_87),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_50),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_73),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_47),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_8),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_158),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_43),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_132),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_51),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_0),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_19),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_56),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_46),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_126),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_130),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_18),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_115),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_56),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_66),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_198),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_91),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_142),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_29),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_182),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_164),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_65),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_67),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_2),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_76),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_202),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_191),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_157),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_156),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_31),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_168),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_120),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_143),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_180),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_62),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_46),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_1),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_83),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_54),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_118),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_102),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_81),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_123),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_55),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_167),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_96),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_39),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_109),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_139),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_21),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_47),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_44),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_133),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_64),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_16),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_34),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_28),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_79),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_160),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_199),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_0),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_29),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_43),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_20),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_100),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_35),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_68),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_33),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_173),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_77),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_151),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_64),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_195),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_60),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_177),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_24),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_26),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_67),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_11),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_22),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_15),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_35),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_200),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_50),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_136),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_48),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_39),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_71),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_51),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_116),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_169),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_13),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_206),
.B(n_4),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_279),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_346),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_357),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_279),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_234),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_228),
.B(n_4),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_234),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_272),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_343),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_206),
.B(n_5),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_274),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_323),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_343),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_268),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_229),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_325),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_229),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_228),
.B(n_7),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_226),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_211),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_226),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_217),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_212),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_217),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_212),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_212),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_229),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_212),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_360),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_204),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_219),
.B(n_7),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_367),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_365),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_395),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_395),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_305),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_367),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_219),
.B(n_12),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_378),
.B(n_12),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_398),
.B(n_13),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_380),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_213),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_321),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_204),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_216),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_321),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_230),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_321),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_230),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_359),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_218),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_220),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_222),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_247),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_223),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_247),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_232),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_232),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_242),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_242),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_359),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_359),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_250),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_250),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_244),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_320),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_224),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_384),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_244),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_245),
.B(n_14),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_236),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_384),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_291),
.B(n_14),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_267),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_241),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_243),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_246),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_251),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_267),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_271),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_260),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_263),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_271),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_269),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_273),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_273),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_424),
.B(n_284),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_448),
.A2(n_291),
.B(n_214),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_248),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_409),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_430),
.B(n_245),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_435),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_487),
.Y(n_524)
);

BUFx8_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_433),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_410),
.A2(n_306),
.B1(n_333),
.B2(n_257),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_487),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_487),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_259),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_434),
.B(n_436),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_478),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_446),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_259),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_479),
.B(n_248),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_480),
.B(n_284),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_480),
.B(n_285),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_481),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_454),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_486),
.B(n_248),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_486),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_491),
.B(n_285),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_461),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_491),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_443),
.B(n_289),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_440),
.B(n_265),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g559 ( 
.A1(n_462),
.A2(n_275),
.B(n_265),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_489),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_477),
.B(n_289),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_465),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_468),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_406),
.B(n_275),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_459),
.B(n_299),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_464),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_408),
.B(n_277),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_414),
.B(n_299),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_475),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_423),
.B(n_299),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_501),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_505),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_416),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_508),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_434),
.B(n_214),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_439),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_450),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_442),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_412),
.B(n_415),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_492),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_412),
.B(n_327),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_470),
.B(n_277),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_585),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_513),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_589),
.A2(n_415),
.B1(n_421),
.B2(n_417),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_516),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_516),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_513),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_585),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_569),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_581),
.B(n_405),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_581),
.B(n_405),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_539),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_586),
.B(n_411),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_586),
.B(n_411),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_546),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_560),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_539),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_586),
.B(n_438),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_SL g610 ( 
.A(n_586),
.B(n_417),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_526),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_539),
.B(n_214),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_587),
.B(n_438),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_518),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_530),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_568),
.A2(n_407),
.B1(n_428),
.B2(n_413),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_523),
.B(n_484),
.Y(n_622)
);

AO22x2_ASAP7_75t_L g623 ( 
.A1(n_527),
.A2(n_306),
.B1(n_333),
.B2(n_257),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_586),
.B(n_441),
.Y(n_624)
);

AO22x2_ASAP7_75t_L g625 ( 
.A1(n_527),
.A2(n_369),
.B1(n_342),
.B2(n_327),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_589),
.A2(n_421),
.B1(n_441),
.B2(n_463),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_583),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_530),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_569),
.B(n_404),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_586),
.B(n_288),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_560),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_523),
.B(n_288),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_523),
.B(n_304),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_555),
.B(n_444),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_568),
.A2(n_432),
.B1(n_469),
.B2(n_467),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_579),
.B(n_419),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_527),
.A2(n_369),
.B1(n_472),
.B2(n_466),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

NOR2x1p5_ASAP7_75t_L g639 ( 
.A(n_569),
.B(n_453),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_587),
.B(n_588),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_543),
.Y(n_641)
);

OA22x2_ASAP7_75t_L g642 ( 
.A1(n_590),
.A2(n_502),
.B1(n_485),
.B2(n_474),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_471),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_561),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_523),
.B(n_539),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_534),
.B(n_476),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_523),
.B(n_304),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_536),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_539),
.B(n_310),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_539),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_569),
.B(n_418),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_549),
.B(n_310),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_510),
.B(n_482),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_549),
.B(n_371),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_561),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_568),
.A2(n_429),
.B1(n_451),
.B2(n_431),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_561),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_546),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_515),
.A2(n_488),
.B1(n_493),
.B2(n_476),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_510),
.B(n_483),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_536),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_546),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_536),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_561),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_580),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_511),
.B(n_490),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_SL g669 ( 
.A(n_590),
.B(n_504),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_488),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_543),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_543),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_543),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_549),
.B(n_312),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_549),
.B(n_312),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_543),
.Y(n_676)
);

BUFx10_ASAP7_75t_L g677 ( 
.A(n_549),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_549),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_543),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_582),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_544),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_544),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_590),
.B(n_493),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_512),
.B(n_498),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_543),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_582),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_515),
.A2(n_498),
.B1(n_500),
.B2(n_499),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_544),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_511),
.B(n_545),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_583),
.B(n_473),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_580),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_543),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_545),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_565),
.B(n_293),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_511),
.B(n_499),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_550),
.B(n_500),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_550),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_550),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_512),
.B(n_506),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_543),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_554),
.B(n_331),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_568),
.B(n_371),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_568),
.A2(n_494),
.B1(n_295),
.B2(n_297),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_582),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_568),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_554),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_572),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_558),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_554),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_558),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_562),
.A2(n_295),
.B1(n_297),
.B2(n_293),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_562),
.B(n_506),
.C(n_280),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_572),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_558),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_582),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_576),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_558),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_562),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_558),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_555),
.B(n_270),
.Y(n_721)
);

AND2x6_ASAP7_75t_L g722 ( 
.A(n_512),
.B(n_371),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_SL g723 ( 
.A(n_553),
.B(n_452),
.C(n_281),
.Y(n_723)
);

BUFx4f_ASAP7_75t_L g724 ( 
.A(n_559),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_582),
.B(n_420),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_558),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_535),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_573),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_562),
.A2(n_366),
.B1(n_332),
.B2(n_334),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_555),
.A2(n_283),
.B1(n_329),
.B2(n_403),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_540),
.B(n_308),
.Y(n_732)
);

OR2x6_ASAP7_75t_L g733 ( 
.A(n_565),
.B(n_308),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_644),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_683),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_646),
.B(n_614),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_634),
.B(n_540),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_599),
.B(n_570),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_640),
.B(n_576),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_613),
.B(n_580),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_598),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_592),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_596),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_644),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_601),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_625),
.A2(n_565),
.B1(n_575),
.B2(n_572),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_697),
.B(n_576),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_598),
.B(n_553),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_600),
.B(n_570),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_696),
.B(n_575),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_613),
.B(n_580),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_706),
.B(n_575),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_622),
.B(n_540),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_613),
.B(n_580),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_594),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_622),
.B(n_540),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_706),
.B(n_541),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_611),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_719),
.B(n_541),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_657),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_591),
.B(n_570),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_591),
.B(n_517),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_615),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_651),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_719),
.B(n_541),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_724),
.B(n_678),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_636),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_610),
.A2(n_573),
.B1(n_577),
.B2(n_574),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_591),
.B(n_517),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_619),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_602),
.B(n_608),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_625),
.A2(n_722),
.B1(n_703),
.B2(n_623),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_628),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_597),
.B(n_517),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_634),
.B(n_551),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_597),
.B(n_566),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_634),
.B(n_551),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_648),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_625),
.A2(n_722),
.B1(n_703),
.B2(n_623),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_724),
.B(n_580),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_657),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_722),
.B(n_580),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_577),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_649),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_722),
.A2(n_578),
.B1(n_577),
.B2(n_531),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_595),
.B(n_566),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_670),
.B(n_578),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_593),
.A2(n_531),
.B1(n_538),
.B2(n_521),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_670),
.B(n_578),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_659),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_659),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_684),
.B(n_521),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_684),
.B(n_521),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_606),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_724),
.B(n_580),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_663),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_666),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_700),
.B(n_531),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_700),
.B(n_609),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_689),
.A2(n_538),
.B(n_514),
.C(n_563),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_665),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_624),
.B(n_584),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_727),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_681),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_682),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_727),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_688),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_693),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_624),
.B(n_584),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_678),
.B(n_651),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_627),
.B(n_566),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_694),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_639),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_698),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_680),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_606),
.Y(n_817)
);

BUFx5_ASAP7_75t_L g818 ( 
.A(n_722),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_626),
.B(n_571),
.C(n_567),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_651),
.B(n_677),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_699),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_707),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_643),
.A2(n_571),
.B1(n_567),
.B2(n_564),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_677),
.B(n_563),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_690),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_677),
.B(n_717),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_722),
.A2(n_564),
.B1(n_563),
.B2(n_567),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_710),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_717),
.B(n_708),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_728),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_732),
.B(n_645),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_709),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_709),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_732),
.B(n_525),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_597),
.B(n_655),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_717),
.B(n_563),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_645),
.B(n_525),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_629),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_711),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_690),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_689),
.B(n_525),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_703),
.B(n_525),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_680),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_711),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_662),
.B(n_579),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_715),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_625),
.A2(n_559),
.B1(n_525),
.B2(n_564),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_632),
.A2(n_633),
.B(n_647),
.C(n_630),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_612),
.B(n_564),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_723),
.B(n_661),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_668),
.B(n_603),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_612),
.B(n_276),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_703),
.B(n_525),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_703),
.B(n_556),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_715),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_612),
.B(n_282),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_718),
.Y(n_857)
);

OR2x6_ASAP7_75t_L g858 ( 
.A(n_629),
.B(n_571),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_718),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_708),
.B(n_514),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_703),
.B(n_556),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_708),
.B(n_514),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_L g863 ( 
.A(n_612),
.B(n_292),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_686),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_714),
.B(n_686),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_704),
.B(n_422),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_635),
.B(n_725),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_714),
.B(n_514),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_603),
.B(n_557),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_621),
.A2(n_294),
.B1(n_298),
.B2(n_296),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_605),
.B(n_557),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_612),
.B(n_656),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_631),
.Y(n_873)
);

OR2x2_ASAP7_75t_SL g874 ( 
.A(n_637),
.B(n_426),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_714),
.B(n_331),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_720),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_720),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_705),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_623),
.A2(n_559),
.B1(n_557),
.B2(n_552),
.Y(n_879)
);

NAND2xp33_ASAP7_75t_L g880 ( 
.A(n_612),
.B(n_301),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_726),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_705),
.B(n_338),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_716),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_716),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_726),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_652),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_605),
.B(n_535),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_631),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_656),
.B(n_535),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_656),
.B(n_535),
.Y(n_890)
);

NAND2x1_ASAP7_75t_L g891 ( 
.A(n_656),
.B(n_519),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_656),
.B(n_695),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_652),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_734),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_800),
.A2(n_630),
.B(n_632),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_736),
.B(n_713),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_825),
.B(n_658),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_780),
.A2(n_616),
.B(n_650),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_734),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_738),
.A2(n_623),
.B(n_731),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_809),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_795),
.A2(n_616),
.B(n_650),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_766),
.A2(n_616),
.B(n_654),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_786),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_800),
.A2(n_647),
.B(n_633),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_744),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_840),
.B(n_687),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_835),
.B(n_669),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_766),
.A2(n_674),
.B(n_654),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_798),
.B(n_792),
.Y(n_910)
);

O2A1O1Ixp5_ASAP7_75t_L g911 ( 
.A1(n_823),
.A2(n_674),
.B(n_675),
.C(n_702),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_744),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_794),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_760),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_793),
.B(n_695),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_867),
.B(n_695),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_739),
.A2(n_675),
.B(n_667),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_L g918 ( 
.A(n_762),
.B(n_669),
.C(n_324),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_818),
.B(n_641),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_851),
.A2(n_702),
.B(n_729),
.C(n_712),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_749),
.B(n_799),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_794),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_812),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_767),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_836),
.A2(n_691),
.B(n_667),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_760),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_788),
.B(n_733),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_860),
.A2(n_339),
.B(n_338),
.Y(n_928)
);

NOR2x2_ASAP7_75t_L g929 ( 
.A(n_858),
.B(n_629),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_753),
.B(n_733),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_818),
.B(n_641),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_809),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_735),
.A2(n_660),
.B1(n_664),
.B2(n_652),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_750),
.A2(n_309),
.B(n_303),
.Y(n_934)
);

AOI21x1_ASAP7_75t_L g935 ( 
.A1(n_862),
.A2(n_868),
.B(n_810),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_747),
.A2(n_730),
.B(n_664),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_753),
.B(n_733),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_794),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_818),
.B(n_641),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_868),
.A2(n_660),
.B(n_671),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_815),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_755),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_815),
.Y(n_943)
);

BUFx8_ASAP7_75t_L g944 ( 
.A(n_814),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_845),
.A2(n_656),
.B1(n_733),
.B2(n_653),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_769),
.Y(n_946)
);

AOI21x1_ASAP7_75t_L g947 ( 
.A1(n_803),
.A2(n_617),
.B(n_607),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_831),
.B(n_629),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_774),
.B(n_324),
.C(n_322),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_870),
.A2(n_322),
.B(n_334),
.C(n_332),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_794),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_756),
.B(n_642),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_817),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_756),
.B(n_653),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_756),
.B(n_653),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_787),
.B(n_653),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_829),
.A2(n_826),
.B(n_824),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_789),
.B(n_672),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_771),
.A2(n_672),
.B1(n_679),
.B2(n_673),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_819),
.A2(n_617),
.B(n_607),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_775),
.B(n_620),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_781),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_764),
.A2(n_701),
.B1(n_692),
.B2(n_685),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_737),
.B(n_679),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_759),
.B(n_685),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_740),
.A2(n_701),
.B(n_692),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_830),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_765),
.B(n_783),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_817),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_737),
.B(n_777),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_740),
.A2(n_620),
.B(n_604),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_776),
.B(n_866),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_L g973 ( 
.A1(n_761),
.A2(n_313),
.B(n_311),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_757),
.A2(n_388),
.B(n_399),
.C(n_335),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_818),
.B(n_641),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_742),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_892),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_848),
.A2(n_399),
.B(n_397),
.C(n_335),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_743),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_781),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_751),
.A2(n_604),
.B(n_631),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_841),
.A2(n_559),
.B(n_532),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_L g983 ( 
.A(n_850),
.B(n_375),
.C(n_366),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_817),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_864),
.B(n_676),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_817),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_745),
.B(n_676),
.Y(n_987)
);

AO21x1_ASAP7_75t_L g988 ( 
.A1(n_887),
.A2(n_351),
.B(n_350),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_854),
.A2(n_559),
.B(n_316),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_838),
.B(n_559),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_758),
.B(n_676),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_751),
.A2(n_604),
.B(n_631),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_763),
.B(n_537),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_858),
.B(n_559),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_754),
.A2(n_604),
.B(n_638),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_767),
.B(n_537),
.Y(n_996)
);

CKINVDCx10_ASAP7_75t_R g997 ( 
.A(n_741),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_893),
.A2(n_618),
.B(n_542),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_754),
.A2(n_893),
.B(n_875),
.Y(n_999)
);

AOI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_861),
.A2(n_317),
.B(n_315),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_764),
.A2(n_373),
.B1(n_318),
.B2(n_385),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_785),
.A2(n_397),
.B(n_381),
.C(n_375),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_790),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_875),
.A2(n_604),
.B(n_638),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_874),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_770),
.B(n_537),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_790),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_773),
.B(n_542),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_778),
.B(n_542),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_791),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_784),
.B(n_547),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_843),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_741),
.B(n_547),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_843),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_796),
.B(n_547),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_791),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_878),
.B(n_638),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_827),
.A2(n_886),
.B(n_833),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_814),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_802),
.B(n_547),
.Y(n_1020)
);

AND2x4_ASAP7_75t_SL g1021 ( 
.A(n_858),
.B(n_548),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_818),
.B(n_638),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_805),
.B(n_548),
.Y(n_1023)
);

AO21x1_ASAP7_75t_L g1024 ( 
.A1(n_834),
.A2(n_394),
.B(n_351),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_797),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_806),
.B(n_548),
.Y(n_1026)
);

OAI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_768),
.A2(n_345),
.B(n_319),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_808),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_813),
.B(n_548),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_818),
.B(n_618),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_752),
.A2(n_349),
.B(n_347),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_811),
.A2(n_618),
.B(n_532),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_869),
.A2(n_388),
.B(n_381),
.C(n_552),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_811),
.A2(n_618),
.B(n_532),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_871),
.A2(n_532),
.B(n_509),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_820),
.B(n_362),
.C(n_361),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_821),
.B(n_552),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_822),
.B(n_552),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_828),
.B(n_394),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_746),
.B(n_364),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_858),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_820),
.A2(n_509),
.B(n_519),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_772),
.B(n_368),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_882),
.A2(n_396),
.B(n_327),
.C(n_342),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_832),
.A2(n_520),
.B(n_519),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_816),
.A2(n_883),
.B1(n_884),
.B2(n_865),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_816),
.B(n_837),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_818),
.B(n_396),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_865),
.A2(n_509),
.B(n_519),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_832),
.A2(n_509),
.B(n_519),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_L g1051 ( 
.A(n_873),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_849),
.A2(n_342),
.B(n_291),
.C(n_390),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_816),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_873),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_779),
.B(n_372),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_839),
.A2(n_524),
.B(n_520),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_891),
.B(n_374),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_797),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_839),
.B(n_377),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_844),
.A2(n_524),
.B(n_520),
.Y(n_1060)
);

OAI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_882),
.A2(n_383),
.B(n_379),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_873),
.B(n_520),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_846),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_889),
.A2(n_528),
.B(n_524),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_846),
.A2(n_528),
.B(n_524),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_855),
.B(n_387),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_L g1067 ( 
.A1(n_890),
.A2(n_528),
.B(n_524),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_857),
.A2(n_529),
.B(n_528),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_SL g1069 ( 
.A1(n_972),
.A2(n_748),
.B1(n_856),
.B2(n_852),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_SL g1070 ( 
.A(n_1001),
.B(n_391),
.C(n_389),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_896),
.A2(n_908),
.B(n_946),
.C(n_921),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_SL g1072 ( 
.A1(n_910),
.A2(n_876),
.B(n_885),
.C(n_881),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_942),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_968),
.A2(n_782),
.B(n_849),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_896),
.A2(n_852),
.B(n_856),
.C(n_863),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_921),
.B(n_857),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_944),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_970),
.B(n_859),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_927),
.A2(n_863),
.B(n_880),
.C(n_872),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_904),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_915),
.A2(n_847),
.B1(n_879),
.B2(n_881),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1051),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_1051),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_996),
.B(n_923),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_967),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_R g1086 ( 
.A(n_997),
.B(n_880),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_956),
.A2(n_885),
.B(n_877),
.C(n_859),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_976),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_1012),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_956),
.A2(n_853),
.B1(n_842),
.B2(n_392),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_907),
.B(n_877),
.Y(n_1091)
);

NAND2x1_ASAP7_75t_L g1092 ( 
.A(n_1054),
.B(n_888),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_SL g1093 ( 
.A(n_973),
.B(n_400),
.C(n_393),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_979),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_916),
.B(n_804),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_1019),
.Y(n_1096)
);

CKINVDCx8_ASAP7_75t_R g1097 ( 
.A(n_1041),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_922),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_897),
.B(n_804),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_1019),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_944),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1028),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_920),
.B(n_807),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_954),
.B(n_801),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_920),
.B(n_801),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_900),
.A2(n_291),
.B(n_528),
.C(n_529),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_901),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_948),
.B(n_888),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_1012),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_924),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_948),
.B(n_888),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_932),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_SL g1113 ( 
.A(n_955),
.B(n_203),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_911),
.A2(n_533),
.B(n_529),
.C(n_528),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_936),
.A2(n_533),
.B(n_529),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_941),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_894),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_949),
.B(n_15),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_940),
.A2(n_533),
.B(n_529),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_943),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_SL g1121 ( 
.A(n_1027),
.B(n_209),
.C(n_402),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_945),
.B(n_205),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_950),
.A2(n_533),
.B(n_529),
.C(n_20),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_990),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_918),
.A2(n_533),
.B(n_18),
.C(n_22),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_930),
.B(n_207),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1063),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_983),
.B(n_215),
.C(n_401),
.Y(n_1128)
);

NAND2x1_ASAP7_75t_L g1129 ( 
.A(n_1054),
.B(n_533),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_SL g1130 ( 
.A(n_1013),
.B(n_210),
.C(n_386),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_958),
.A2(n_208),
.B(n_382),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_964),
.B(n_221),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_1005),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_937),
.B(n_225),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_978),
.A2(n_17),
.B(n_23),
.C(n_24),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_964),
.B(n_227),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_913),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_952),
.A2(n_1014),
.B1(n_1040),
.B2(n_977),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1014),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_977),
.B(n_26),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_978),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1043),
.A2(n_231),
.B1(n_376),
.B2(n_370),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1047),
.A2(n_290),
.B(n_235),
.C(n_363),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1000),
.B(n_233),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1057),
.B(n_30),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1061),
.B(n_237),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_957),
.A2(n_302),
.B(n_239),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_971),
.A2(n_307),
.B(n_240),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_961),
.B(n_1047),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_938),
.B(n_238),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_913),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_913),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_951),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_966),
.A2(n_965),
.B(n_925),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1066),
.B(n_32),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_913),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_993),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1002),
.A2(n_353),
.B1(n_262),
.B2(n_261),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_895),
.A2(n_249),
.B(n_252),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_953),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_960),
.A2(n_326),
.B(n_254),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1002),
.A2(n_358),
.B1(n_255),
.B2(n_253),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1066),
.B(n_1039),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1006),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1057),
.B(n_32),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_922),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_974),
.A2(n_934),
.B(n_1052),
.C(n_1031),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1053),
.B(n_256),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1055),
.A2(n_905),
.B1(n_969),
.B2(n_929),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_953),
.B(n_258),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_961),
.A2(n_933),
.B1(n_1038),
.B2(n_1037),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_909),
.A2(n_330),
.B(n_266),
.C(n_356),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1008),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_969),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1053),
.B(n_899),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_899),
.B(n_33),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_953),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1022),
.A2(n_336),
.B(n_278),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1009),
.A2(n_264),
.B1(n_286),
.B2(n_287),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_951),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1036),
.B(n_1059),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1011),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_953),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_919),
.A2(n_939),
.B(n_931),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1015),
.A2(n_1029),
.B1(n_1020),
.B2(n_1023),
.Y(n_1185)
);

AND2x2_ASAP7_75t_SL g1186 ( 
.A(n_1021),
.B(n_320),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_938),
.B(n_300),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1052),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_947),
.A2(n_522),
.B(n_518),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1046),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_906),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_912),
.B(n_40),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1021),
.B(n_40),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_R g1194 ( 
.A(n_984),
.B(n_314),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_994),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_984),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_41),
.B(n_42),
.C(n_48),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1033),
.A2(n_41),
.B(n_42),
.C(n_49),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1003),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_986),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_898),
.A2(n_348),
.B(n_337),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_986),
.B(n_49),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_986),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_986),
.B(n_344),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_912),
.B(n_52),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_987),
.B(n_991),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1048),
.A2(n_355),
.B1(n_352),
.B2(n_341),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_999),
.A2(n_328),
.B(n_320),
.C(n_522),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_914),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_919),
.A2(n_931),
.B(n_939),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_SL g1211 ( 
.A(n_1048),
.B(n_320),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_985),
.B(n_1017),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1018),
.A2(n_320),
.B1(n_53),
.B2(n_55),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_975),
.A2(n_518),
.B(n_522),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1062),
.B(n_52),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_975),
.A2(n_522),
.B(n_518),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_985),
.A2(n_522),
.B1(n_518),
.B2(n_60),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_917),
.A2(n_992),
.B(n_995),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1071),
.B(n_1017),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1082),
.B(n_926),
.Y(n_1220)
);

AOI221x1_ASAP7_75t_L g1221 ( 
.A1(n_1213),
.A2(n_1155),
.B1(n_1138),
.B2(n_1075),
.C(n_1169),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1213),
.A2(n_1044),
.B(n_963),
.C(n_1062),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1209),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1073),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1149),
.A2(n_903),
.B1(n_902),
.B2(n_998),
.Y(n_1225)
);

AOI221x1_ASAP7_75t_L g1226 ( 
.A1(n_1218),
.A2(n_989),
.B1(n_1049),
.B2(n_959),
.C(n_1042),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1149),
.A2(n_1030),
.B(n_1004),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1074),
.A2(n_1030),
.B(n_981),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1073),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1185),
.A2(n_1032),
.B(n_1034),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1181),
.B(n_1145),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1084),
.B(n_926),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1099),
.A2(n_1025),
.B1(n_962),
.B2(n_980),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1076),
.A2(n_935),
.B1(n_1045),
.B2(n_1016),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1167),
.A2(n_1068),
.B(n_1056),
.C(n_1065),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1185),
.A2(n_1035),
.B(n_1060),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1091),
.B(n_1058),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1159),
.A2(n_1050),
.B(n_1067),
.Y(n_1238)
);

BUFx4f_ASAP7_75t_L g1239 ( 
.A(n_1101),
.Y(n_1239)
);

INVx3_ASAP7_75t_SL g1240 ( 
.A(n_1101),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1163),
.A2(n_980),
.B(n_1016),
.C(n_1010),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1082),
.B(n_1010),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1083),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1171),
.A2(n_1007),
.B(n_962),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1077),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1089),
.B(n_1109),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1200),
.B(n_1007),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_SL g1248 ( 
.A(n_1118),
.B(n_53),
.C(n_58),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1086),
.Y(n_1249)
);

AO21x1_ASAP7_75t_L g1250 ( 
.A1(n_1212),
.A2(n_982),
.B(n_1064),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1180),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1079),
.A2(n_1210),
.B(n_1184),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1078),
.A2(n_522),
.B(n_518),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1139),
.B(n_61),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1123),
.A2(n_522),
.B(n_518),
.C(n_68),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1103),
.A2(n_518),
.A3(n_113),
.B(n_119),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1080),
.B(n_63),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1100),
.B(n_66),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1126),
.B(n_69),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1134),
.B(n_69),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1119),
.A2(n_128),
.B(n_196),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1096),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1105),
.A2(n_108),
.A3(n_194),
.B(n_190),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1125),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_1264)
);

OAI22x1_ASAP7_75t_L g1265 ( 
.A1(n_1145),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1208),
.A2(n_80),
.A3(n_82),
.B(n_84),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1110),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1146),
.A2(n_93),
.B(n_95),
.C(n_98),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1115),
.A2(n_101),
.B(n_135),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1214),
.A2(n_140),
.B(n_150),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1083),
.B(n_201),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1087),
.A2(n_153),
.A3(n_174),
.B(n_178),
.Y(n_1272)
);

AOI221xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1190),
.A2(n_186),
.B1(n_1135),
.B2(n_1141),
.C(n_1198),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1165),
.B(n_1130),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1143),
.A2(n_1172),
.B(n_1092),
.C(n_1108),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1216),
.A2(n_1106),
.B(n_1192),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1165),
.B(n_1097),
.Y(n_1277)
);

AO22x1_ASAP7_75t_L g1278 ( 
.A1(n_1193),
.A2(n_1202),
.B1(n_1203),
.B2(n_1158),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1179),
.A2(n_1162),
.B(n_1158),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1069),
.A2(n_1168),
.B1(n_1140),
.B2(n_1142),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1192),
.A2(n_1175),
.B(n_1111),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1217),
.A2(n_1070),
.B1(n_1182),
.B2(n_1173),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1193),
.A2(n_1162),
.B1(n_1122),
.B2(n_1093),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1137),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1094),
.B(n_1102),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1179),
.A2(n_1161),
.B(n_1114),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1191),
.A2(n_1211),
.A3(n_1164),
.B(n_1157),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1072),
.A2(n_1201),
.B(n_1206),
.Y(n_1289)
);

AND2x6_ASAP7_75t_L g1290 ( 
.A(n_1202),
.B(n_1195),
.Y(n_1290)
);

AOI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1148),
.A2(n_1144),
.B(n_1176),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1201),
.A2(n_1129),
.B(n_1127),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1187),
.A2(n_1131),
.B(n_1147),
.Y(n_1293)
);

NAND3x1_ASAP7_75t_L g1294 ( 
.A(n_1215),
.B(n_1205),
.C(n_1095),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1121),
.A2(n_1188),
.B(n_1090),
.C(n_1104),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1206),
.A2(n_1120),
.B(n_1107),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1166),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1199),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1194),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1177),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1098),
.A2(n_1174),
.B(n_1170),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1206),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1195),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_SL g1304 ( 
.A1(n_1204),
.A2(n_1197),
.B(n_1136),
.C(n_1132),
.Y(n_1304)
);

AOI221x1_ASAP7_75t_L g1305 ( 
.A1(n_1113),
.A2(n_1178),
.B1(n_1128),
.B2(n_1160),
.C(n_1156),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1153),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1124),
.A2(n_1196),
.B(n_1207),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1186),
.A2(n_1152),
.B(n_1183),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1150),
.B(n_1133),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1152),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1151),
.B(n_1156),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1183),
.A2(n_1151),
.B1(n_1160),
.B2(n_896),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1151),
.A2(n_1149),
.B(n_1074),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1160),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1117),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1189),
.A2(n_1154),
.B(n_1218),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1071),
.A2(n_896),
.B1(n_736),
.B2(n_946),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1071),
.B(n_946),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1149),
.A2(n_1074),
.B(n_1185),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1081),
.A2(n_1024),
.A3(n_988),
.B(n_928),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1081),
.A2(n_1024),
.A3(n_988),
.B(n_928),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1071),
.B(n_946),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1071),
.A2(n_896),
.B(n_908),
.C(n_736),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1189),
.A2(n_1154),
.B(n_1218),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1082),
.B(n_1200),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1081),
.A2(n_1024),
.A3(n_988),
.B(n_928),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1084),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1137),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_SL g1329 ( 
.A1(n_1071),
.A2(n_1149),
.B(n_1075),
.C(n_927),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1209),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1189),
.A2(n_1154),
.B(n_1218),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1071),
.A2(n_896),
.B1(n_736),
.B2(n_946),
.Y(n_1332)
);

AOI211x1_ASAP7_75t_L g1333 ( 
.A1(n_1213),
.A2(n_927),
.B(n_1155),
.C(n_910),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1071),
.B(n_825),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1071),
.A2(n_896),
.B1(n_736),
.B2(n_946),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1082),
.B(n_1200),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1082),
.B(n_1200),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1118),
.A2(n_896),
.B1(n_738),
.B2(n_749),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1081),
.A2(n_1024),
.A3(n_988),
.B(n_928),
.Y(n_1339)
);

NAND3xp33_ASAP7_75t_L g1340 ( 
.A(n_1071),
.B(n_908),
.C(n_736),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1100),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1071),
.B(n_825),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_SL g1343 ( 
.A(n_1100),
.B(n_579),
.Y(n_1343)
);

INVx6_ASAP7_75t_L g1344 ( 
.A(n_1100),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1101),
.B(n_1019),
.Y(n_1345)
);

AOI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1146),
.A2(n_908),
.B(n_749),
.Y(n_1346)
);

AOI221xp5_ASAP7_75t_L g1347 ( 
.A1(n_1071),
.A2(n_637),
.B1(n_527),
.B2(n_749),
.C(n_738),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1073),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1209),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1071),
.B(n_825),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1071),
.A2(n_1125),
.B1(n_1190),
.B2(n_896),
.C(n_950),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1071),
.A2(n_736),
.B(n_896),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1071),
.B(n_825),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1149),
.A2(n_1074),
.B(n_1185),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1083),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1084),
.A2(n_749),
.B1(n_738),
.B2(n_908),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1073),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1189),
.A2(n_1154),
.B(n_1218),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1071),
.A2(n_896),
.B(n_908),
.C(n_736),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1071),
.A2(n_896),
.B1(n_736),
.B2(n_946),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1083),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1071),
.B(n_946),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1071),
.B(n_825),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1081),
.A2(n_1024),
.A3(n_988),
.B(n_928),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1209),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1209),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1071),
.B(n_946),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1110),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1073),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1071),
.B(n_825),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1071),
.B(n_946),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1240),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1338),
.A2(n_1371),
.B1(n_1318),
.B2(n_1322),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1347),
.A2(n_1338),
.B1(n_1346),
.B2(n_1352),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1249),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1285),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1317),
.B(n_1332),
.Y(n_1377)
);

BUFx10_ASAP7_75t_L g1378 ( 
.A(n_1277),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1356),
.A2(n_1359),
.B1(n_1323),
.B2(n_1340),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1231),
.A2(n_1280),
.B1(n_1343),
.B2(n_1335),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1300),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1224),
.Y(n_1382)
);

INVx3_ASAP7_75t_SL g1383 ( 
.A(n_1341),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1314),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1300),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1279),
.B(n_1360),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1239),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1341),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1345),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1248),
.A2(n_1259),
.B1(n_1260),
.B2(n_1265),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1239),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1229),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1334),
.A2(n_1353),
.B1(n_1370),
.B2(n_1363),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1362),
.A2(n_1367),
.B1(n_1342),
.B2(n_1350),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1274),
.A2(n_1283),
.B1(n_1232),
.B2(n_1284),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1299),
.A2(n_1290),
.B1(n_1219),
.B2(n_1298),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1290),
.A2(n_1307),
.B1(n_1287),
.B2(n_1309),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_L g1399 ( 
.A(n_1345),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1300),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1221),
.A2(n_1258),
.B1(n_1254),
.B2(n_1246),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1344),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1223),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1290),
.A2(n_1298),
.B1(n_1237),
.B2(n_1247),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1290),
.A2(n_1247),
.B1(n_1303),
.B2(n_1307),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1368),
.B(n_1267),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1303),
.A2(n_1330),
.B1(n_1366),
.B2(n_1365),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1344),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1245),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1223),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1251),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1243),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1314),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1369),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1325),
.B(n_1336),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1357),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1314),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1306),
.B(n_1325),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1336),
.Y(n_1419)
);

INVx8_ASAP7_75t_L g1420 ( 
.A(n_1271),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1355),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1257),
.A2(n_1319),
.B1(n_1354),
.B2(n_1351),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1348),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1330),
.A2(n_1366),
.B1(n_1365),
.B2(n_1349),
.Y(n_1424)
);

CKINVDCx9p33_ASAP7_75t_R g1425 ( 
.A(n_1278),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1349),
.A2(n_1233),
.B1(n_1315),
.B2(n_1293),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1337),
.B(n_1294),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1333),
.A2(n_1289),
.B1(n_1271),
.B2(n_1337),
.Y(n_1428)
);

INVx4_ASAP7_75t_L g1429 ( 
.A(n_1328),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1220),
.A2(n_1242),
.B1(n_1333),
.B2(n_1234),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1262),
.B(n_1328),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1310),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1295),
.A2(n_1273),
.B1(n_1302),
.B2(n_1304),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1297),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1220),
.A2(n_1242),
.B1(n_1302),
.B2(n_1244),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_R g1436 ( 
.A1(n_1264),
.A2(n_1329),
.B1(n_1255),
.B2(n_1222),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1311),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1310),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1361),
.B(n_1243),
.Y(n_1439)
);

INVx6_ASAP7_75t_L g1440 ( 
.A(n_1361),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1312),
.Y(n_1441)
);

BUFx2_ASAP7_75t_SL g1442 ( 
.A(n_1308),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1225),
.A2(n_1282),
.B1(n_1250),
.B2(n_1227),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1296),
.A2(n_1292),
.B1(n_1269),
.B2(n_1270),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1301),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1313),
.A2(n_1276),
.B1(n_1238),
.B2(n_1253),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1268),
.A2(n_1275),
.B1(n_1241),
.B2(n_1235),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_1305),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1252),
.A2(n_1230),
.B1(n_1236),
.B2(n_1291),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1261),
.A2(n_1263),
.B1(n_1272),
.B2(n_1326),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1263),
.A2(n_1272),
.B1(n_1364),
.B2(n_1326),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1228),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1263),
.A2(n_1272),
.B1(n_1339),
.B2(n_1326),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1288),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1320),
.B(n_1321),
.Y(n_1455)
);

INVx3_ASAP7_75t_SL g1456 ( 
.A(n_1266),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1320),
.A2(n_1364),
.B1(n_1339),
.B2(n_1321),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1364),
.A2(n_1266),
.B1(n_1256),
.B2(n_1358),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1256),
.A2(n_1316),
.B1(n_1324),
.B2(n_1331),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1266),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1226),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1281),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1281),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1338),
.A2(n_1347),
.B1(n_749),
.B2(n_738),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1281),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1338),
.A2(n_1356),
.B1(n_1347),
.B2(n_927),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1231),
.B(n_1327),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1325),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1338),
.A2(n_1356),
.B1(n_1347),
.B2(n_927),
.Y(n_1469)
);

BUFx8_ASAP7_75t_SL g1470 ( 
.A(n_1239),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1281),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1231),
.B(n_1327),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1281),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1347),
.A2(n_867),
.B1(n_900),
.B2(n_623),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1314),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1338),
.A2(n_1356),
.B1(n_1359),
.B2(n_1323),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1347),
.A2(n_867),
.B1(n_900),
.B2(n_623),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1325),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1280),
.A2(n_867),
.B1(n_623),
.B2(n_749),
.Y(n_1479)
);

BUFx8_ASAP7_75t_L g1480 ( 
.A(n_1357),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1347),
.A2(n_867),
.B1(n_900),
.B2(n_623),
.Y(n_1481)
);

BUFx2_ASAP7_75t_SL g1482 ( 
.A(n_1224),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1314),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1249),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1249),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1338),
.A2(n_1356),
.B1(n_1359),
.B2(n_1323),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1347),
.A2(n_867),
.B1(n_900),
.B2(n_623),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1341),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1347),
.A2(n_867),
.B1(n_900),
.B2(n_623),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1300),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1280),
.A2(n_867),
.B1(n_623),
.B2(n_749),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1281),
.Y(n_1492)
);

NAND2xp33_ASAP7_75t_SL g1493 ( 
.A(n_1317),
.B(n_1086),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1341),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1341),
.Y(n_1495)
);

BUFx2_ASAP7_75t_SL g1496 ( 
.A(n_1224),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1290),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1352),
.B(n_1317),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1249),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1251),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1314),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1341),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1249),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1347),
.A2(n_867),
.B1(n_900),
.B2(n_623),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1223),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1338),
.A2(n_1356),
.B1(n_1359),
.B2(n_1323),
.Y(n_1506)
);

OAI22x1_ASAP7_75t_SL g1507 ( 
.A1(n_1249),
.A2(n_741),
.B1(n_767),
.B2(n_579),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1338),
.A2(n_1347),
.B1(n_749),
.B2(n_738),
.Y(n_1508)
);

BUFx8_ASAP7_75t_SL g1509 ( 
.A(n_1239),
.Y(n_1509)
);

AO22x1_ASAP7_75t_L g1510 ( 
.A1(n_1279),
.A2(n_741),
.B1(n_1274),
.B2(n_769),
.Y(n_1510)
);

BUFx4f_ASAP7_75t_SL g1511 ( 
.A(n_1285),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1403),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1445),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1410),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1497),
.B(n_1505),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1505),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1460),
.A2(n_1443),
.B(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1434),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1424),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1390),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1467),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1395),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1452),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1387),
.B(n_1374),
.C(n_1464),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1455),
.B(n_1457),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1497),
.Y(n_1526)
);

CKINVDCx12_ASAP7_75t_R g1527 ( 
.A(n_1373),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1497),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1387),
.B(n_1377),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1407),
.B(n_1461),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1407),
.Y(n_1531)
);

AND2x4_ASAP7_75t_SL g1532 ( 
.A(n_1417),
.B(n_1475),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1468),
.B(n_1478),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1449),
.A2(n_1459),
.B(n_1443),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1459),
.A2(n_1446),
.B(n_1447),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1386),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1394),
.B(n_1498),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1415),
.B(n_1462),
.Y(n_1538)
);

AOI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1510),
.A2(n_1379),
.B(n_1506),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_R g1540 ( 
.A(n_1372),
.B(n_1376),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1463),
.B(n_1465),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1448),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1399),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1411),
.B(n_1500),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1381),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1471),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1473),
.Y(n_1547)
);

INVxp33_ASAP7_75t_L g1548 ( 
.A(n_1470),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1485),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1492),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1394),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1419),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1451),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1454),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1453),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1426),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1380),
.B(n_1441),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1426),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1472),
.B(n_1374),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1456),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1448),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1466),
.B(n_1469),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1422),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1437),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1406),
.Y(n_1565)
);

O2A1O1Ixp5_ASAP7_75t_L g1566 ( 
.A1(n_1476),
.A2(n_1486),
.B(n_1466),
.C(n_1469),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1427),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1383),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1422),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1435),
.B(n_1430),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1458),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1430),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1417),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1418),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1493),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1446),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1442),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1428),
.B(n_1396),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1432),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1405),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1405),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1450),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1398),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1433),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1404),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1479),
.A2(n_1491),
.B1(n_1474),
.B2(n_1481),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1404),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1436),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1444),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1401),
.B(n_1396),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1401),
.B(n_1397),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1475),
.B(n_1483),
.Y(n_1592)
);

BUFx4f_ASAP7_75t_SL g1593 ( 
.A(n_1392),
.Y(n_1593)
);

AOI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1439),
.A2(n_1431),
.B(n_1408),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1388),
.B(n_1507),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1438),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1483),
.B(n_1501),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1509),
.B(n_1399),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1483),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1384),
.B(n_1501),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1508),
.A2(n_1420),
.B(n_1391),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1381),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1397),
.B(n_1391),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1474),
.A2(n_1504),
.B(n_1477),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1383),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1413),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1413),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1425),
.Y(n_1608)
);

NOR2xp67_ASAP7_75t_L g1609 ( 
.A(n_1400),
.B(n_1429),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1389),
.B(n_1502),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1522),
.B(n_1429),
.Y(n_1611)
);

INVx5_ASAP7_75t_L g1612 ( 
.A(n_1526),
.Y(n_1612)
);

OAI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1537),
.A2(n_1524),
.B(n_1539),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1590),
.A2(n_1425),
.B1(n_1481),
.B2(n_1504),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1523),
.B(n_1495),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1593),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1523),
.B(n_1533),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1524),
.A2(n_1489),
.B(n_1477),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1566),
.A2(n_1489),
.B(n_1487),
.C(n_1488),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_SL g1620 ( 
.A1(n_1562),
.A2(n_1375),
.B(n_1503),
.C(n_1416),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1529),
.B(n_1494),
.Y(n_1621)
);

AOI211xp5_ASAP7_75t_L g1622 ( 
.A1(n_1588),
.A2(n_1414),
.B(n_1389),
.C(n_1409),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1529),
.B(n_1402),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1536),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1601),
.A2(n_1487),
.B(n_1482),
.C(n_1496),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1512),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1546),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1539),
.A2(n_1393),
.B(n_1423),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1549),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1605),
.Y(n_1630)
);

NAND2xp33_ASAP7_75t_R g1631 ( 
.A(n_1608),
.B(n_1499),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1538),
.B(n_1402),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1538),
.B(n_1378),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1594),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1546),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1584),
.A2(n_1557),
.B(n_1551),
.C(n_1603),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1559),
.B(n_1421),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1603),
.A2(n_1421),
.B(n_1385),
.C(n_1490),
.Y(n_1638)
);

NOR2x1_ASAP7_75t_SL g1639 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1527),
.A2(n_1385),
.B1(n_1382),
.B2(n_1412),
.Y(n_1640)
);

AO32x2_ASAP7_75t_L g1641 ( 
.A1(n_1545),
.A2(n_1480),
.A3(n_1440),
.B1(n_1412),
.B2(n_1382),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1559),
.B(n_1440),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1527),
.A2(n_1511),
.B1(n_1480),
.B2(n_1440),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1521),
.B(n_1574),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1515),
.B(n_1511),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1534),
.A2(n_1535),
.B(n_1563),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1552),
.B(n_1592),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1561),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1575),
.A2(n_1520),
.B1(n_1608),
.B2(n_1548),
.Y(n_1649)
);

INVx4_ASAP7_75t_L g1650 ( 
.A(n_1605),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1592),
.B(n_1530),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1575),
.A2(n_1591),
.B1(n_1578),
.B2(n_1586),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1578),
.A2(n_1551),
.B1(n_1570),
.B2(n_1576),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1604),
.A2(n_1530),
.B1(n_1570),
.B2(n_1583),
.Y(n_1654)
);

AO32x2_ASAP7_75t_L g1655 ( 
.A1(n_1602),
.A2(n_1525),
.A3(n_1558),
.B1(n_1556),
.B2(n_1580),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1525),
.B(n_1547),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1568),
.A2(n_1595),
.B1(n_1543),
.B2(n_1544),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1518),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1547),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1550),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1561),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1565),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1563),
.A2(n_1569),
.B(n_1535),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1610),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1569),
.B(n_1577),
.C(n_1582),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1541),
.B(n_1550),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1541),
.B(n_1564),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1610),
.B(n_1597),
.Y(n_1668)
);

BUFx4f_ASAP7_75t_SL g1669 ( 
.A(n_1543),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1599),
.B(n_1567),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1589),
.A2(n_1582),
.B1(n_1571),
.B2(n_1556),
.C(n_1558),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1594),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1604),
.A2(n_1570),
.B1(n_1572),
.B2(n_1571),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1589),
.B(n_1607),
.C(n_1606),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1560),
.A2(n_1581),
.B(n_1580),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1600),
.B(n_1573),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1606),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1532),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1609),
.A2(n_1555),
.B(n_1553),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1641),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1624),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1614),
.A2(n_1570),
.B1(n_1572),
.B2(n_1583),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1658),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1658),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1626),
.Y(n_1686)
);

INVxp67_ASAP7_75t_SL g1687 ( 
.A(n_1648),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1666),
.B(n_1519),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1668),
.B(n_1647),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1644),
.B(n_1579),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1613),
.B(n_1579),
.Y(n_1691)
);

INVx5_ASAP7_75t_L g1692 ( 
.A(n_1612),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1630),
.B(n_1616),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1677),
.B(n_1542),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1674),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1651),
.B(n_1513),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1616),
.Y(n_1697)
);

CKINVDCx14_ASAP7_75t_R g1698 ( 
.A(n_1649),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1630),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1617),
.B(n_1513),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1621),
.B(n_1596),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1648),
.Y(n_1702)
);

INVx5_ASAP7_75t_L g1703 ( 
.A(n_1612),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1627),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1635),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1614),
.A2(n_1604),
.B1(n_1555),
.B2(n_1553),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1611),
.B(n_1596),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1618),
.A2(n_1581),
.B1(n_1587),
.B2(n_1585),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1659),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1661),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1660),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1625),
.A2(n_1526),
.B(n_1528),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1631),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1656),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1654),
.A2(n_1587),
.B1(n_1585),
.B2(n_1554),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1611),
.B(n_1531),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1661),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1676),
.Y(n_1719)
);

NAND2x1p5_ASAP7_75t_SL g1720 ( 
.A(n_1679),
.B(n_1602),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1667),
.B(n_1517),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1678),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1663),
.B(n_1517),
.Y(n_1723)
);

NOR4xp25_ASAP7_75t_L g1724 ( 
.A(n_1683),
.B(n_1636),
.C(n_1620),
.D(n_1619),
.Y(n_1724)
);

OAI33xp33_ASAP7_75t_L g1725 ( 
.A1(n_1716),
.A2(n_1652),
.A3(n_1653),
.B1(n_1657),
.B2(n_1623),
.B3(n_1636),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1719),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1712),
.A2(n_1625),
.B(n_1620),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1684),
.Y(n_1728)
);

AOI211xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1713),
.A2(n_1643),
.B(n_1669),
.C(n_1622),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1681),
.A2(n_1671),
.B1(n_1665),
.B2(n_1654),
.C(n_1628),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1681),
.A2(n_1708),
.B1(n_1706),
.B2(n_1715),
.C(n_1688),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1721),
.B(n_1646),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1685),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1681),
.B(n_1634),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1689),
.B(n_1615),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1681),
.A2(n_1691),
.B1(n_1723),
.B2(n_1675),
.C(n_1719),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1723),
.Y(n_1739)
);

AOI33xp33_ASAP7_75t_L g1740 ( 
.A1(n_1717),
.A2(n_1673),
.A3(n_1633),
.B1(n_1632),
.B2(n_1642),
.B3(n_1637),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1692),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1710),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1721),
.B(n_1646),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1685),
.B(n_1646),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1686),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1682),
.B(n_1718),
.Y(n_1746)
);

OAI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1698),
.A2(n_1650),
.B(n_1640),
.C(n_1680),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1670),
.Y(n_1748)
);

NAND4xp25_ASAP7_75t_L g1749 ( 
.A(n_1697),
.B(n_1631),
.C(n_1619),
.D(n_1650),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1694),
.B(n_1655),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1687),
.A2(n_1639),
.B(n_1638),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1700),
.B(n_1655),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1693),
.A2(n_1645),
.B(n_1540),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.B(n_1655),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1720),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1696),
.B(n_1664),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1710),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1717),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1722),
.B(n_1662),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1692),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1722),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1709),
.B(n_1634),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1696),
.B(n_1664),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1704),
.B(n_1607),
.C(n_1676),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1712),
.A2(n_1645),
.B1(n_1669),
.B2(n_1638),
.Y(n_1765)
);

NOR2x1_ASAP7_75t_SL g1766 ( 
.A(n_1765),
.B(n_1692),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1762),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1745),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1726),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1745),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1728),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1730),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1762),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1732),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1730),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1752),
.B(n_1705),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1735),
.B(n_1711),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1754),
.B(n_1701),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1726),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1760),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1760),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1760),
.B(n_1692),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1735),
.B(n_1758),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1725),
.B(n_1697),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1690),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1750),
.B(n_1707),
.Y(n_1786)
);

INVxp33_ASAP7_75t_L g1787 ( 
.A(n_1751),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1736),
.B(n_1692),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1744),
.B(n_1695),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_L g1790 ( 
.A(n_1749),
.B(n_1540),
.C(n_1672),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1744),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1726),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1736),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1734),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1736),
.B(n_1703),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1761),
.B(n_1695),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1742),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1742),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1734),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1741),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1703),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1755),
.B(n_1703),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1739),
.B(n_1720),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1771),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1771),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1769),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1769),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1772),
.Y(n_1811)
);

NAND2x1_ASAP7_75t_L g1812 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1772),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1772),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1786),
.B(n_1793),
.Y(n_1816)
);

AOI32xp33_ASAP7_75t_L g1817 ( 
.A1(n_1787),
.A2(n_1738),
.A3(n_1731),
.B1(n_1733),
.B2(n_1729),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1780),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1775),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1780),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1787),
.A2(n_1724),
.B1(n_1749),
.B2(n_1739),
.C(n_1764),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1775),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1769),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1775),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1786),
.B(n_1756),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1774),
.B(n_1740),
.Y(n_1826)
);

INVxp67_ASAP7_75t_SL g1827 ( 
.A(n_1791),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1777),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1796),
.B(n_1746),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1774),
.B(n_1724),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1777),
.Y(n_1831)
);

NOR2x1p5_ASAP7_75t_L g1832 ( 
.A(n_1800),
.B(n_1699),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1757),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1768),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1786),
.B(n_1756),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1793),
.B(n_1763),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1797),
.B(n_1757),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1768),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1779),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1798),
.B(n_1737),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1768),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1798),
.B(n_1737),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1779),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1796),
.B(n_1748),
.Y(n_1844)
);

AND2x2_ASAP7_75t_SL g1845 ( 
.A(n_1790),
.B(n_1741),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1790),
.A2(n_1727),
.B1(n_1765),
.B2(n_1739),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1766),
.B(n_1741),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1770),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1779),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1783),
.B(n_1789),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1850),
.B(n_1783),
.Y(n_1851)
);

AND2x4_ASAP7_75t_SL g1852 ( 
.A(n_1836),
.B(n_1782),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1793),
.Y(n_1853)
);

AND2x4_ASAP7_75t_SL g1854 ( 
.A(n_1836),
.B(n_1782),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1825),
.B(n_1835),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1835),
.B(n_1788),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1816),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1808),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1830),
.B(n_1778),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1833),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1850),
.B(n_1789),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1813),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1827),
.B(n_1776),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1828),
.B(n_1776),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1820),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1816),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1832),
.B(n_1788),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1826),
.B(n_1778),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1831),
.B(n_1776),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1844),
.B(n_1789),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1805),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1805),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1844),
.B(n_1799),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1806),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1840),
.B(n_1778),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1847),
.B(n_1788),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1829),
.B(n_1799),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1842),
.B(n_1778),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1847),
.B(n_1788),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1847),
.B(n_1795),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1806),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1829),
.B(n_1785),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1817),
.B(n_1785),
.Y(n_1883)
);

AND2x2_ASAP7_75t_SL g1884 ( 
.A(n_1845),
.B(n_1820),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1785),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1845),
.B(n_1795),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1811),
.Y(n_1887)
);

NOR2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1857),
.B(n_1812),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1855),
.B(n_1818),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1883),
.A2(n_1821),
.B(n_1846),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1871),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1871),
.Y(n_1892)
);

NAND3xp33_ASAP7_75t_L g1893 ( 
.A(n_1858),
.B(n_1862),
.C(n_1884),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1853),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1872),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1859),
.A2(n_1791),
.B(n_1818),
.C(n_1729),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1855),
.B(n_1767),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1872),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1874),
.Y(n_1899)
);

NAND2xp33_ASAP7_75t_SL g1900 ( 
.A(n_1857),
.B(n_1812),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1853),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1865),
.B(n_1857),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1868),
.A2(n_1766),
.B1(n_1794),
.B2(n_1801),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1860),
.A2(n_1863),
.B1(n_1801),
.B2(n_1799),
.C(n_1794),
.Y(n_1904)
);

OAI321xp33_ASAP7_75t_L g1905 ( 
.A1(n_1863),
.A2(n_1804),
.A3(n_1747),
.B1(n_1803),
.B2(n_1802),
.C(n_1764),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1874),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1865),
.B(n_1767),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1884),
.A2(n_1804),
.B1(n_1818),
.B2(n_1800),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1884),
.A2(n_1803),
.B(n_1802),
.Y(n_1909)
);

NOR3xp33_ASAP7_75t_L g1910 ( 
.A(n_1866),
.B(n_1809),
.C(n_1807),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1866),
.B(n_1882),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1881),
.Y(n_1912)
);

OAI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1870),
.A2(n_1804),
.B1(n_1861),
.B2(n_1875),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1881),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1866),
.Y(n_1915)
);

A2O1A1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1890),
.A2(n_1861),
.B(n_1870),
.C(n_1886),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1893),
.A2(n_1886),
.B1(n_1854),
.B2(n_1852),
.Y(n_1917)
);

O2A1O1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1905),
.A2(n_1851),
.B(n_1877),
.C(n_1887),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1914),
.Y(n_1919)
);

OAI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1896),
.A2(n_1877),
.B(n_1851),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1894),
.B(n_1901),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1902),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1914),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1901),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1903),
.A2(n_1854),
.B1(n_1852),
.B2(n_1885),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1902),
.B(n_1852),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1913),
.A2(n_1801),
.B1(n_1794),
.B2(n_1887),
.C(n_1864),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1891),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1892),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1895),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1911),
.B(n_1856),
.Y(n_1931)
);

AOI332xp33_ASAP7_75t_L g1932 ( 
.A1(n_1898),
.A2(n_1864),
.A3(n_1869),
.B1(n_1880),
.B2(n_1879),
.B3(n_1876),
.C1(n_1841),
.C2(n_1834),
.Y(n_1932)
);

OAI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1909),
.A2(n_1873),
.B1(n_1878),
.B2(n_1869),
.Y(n_1933)
);

INVxp33_ASAP7_75t_L g1934 ( 
.A(n_1889),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1899),
.Y(n_1935)
);

XNOR2x1_ASAP7_75t_L g1936 ( 
.A(n_1920),
.B(n_1921),
.Y(n_1936)
);

XNOR2x2_ASAP7_75t_L g1937 ( 
.A(n_1926),
.B(n_1908),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1924),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1922),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1916),
.B(n_1889),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1915),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1927),
.A2(n_1910),
.B1(n_1904),
.B2(n_1794),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1919),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1916),
.B(n_1934),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1923),
.Y(n_1945)
);

O2A1O1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1918),
.A2(n_1907),
.B(n_1912),
.C(n_1906),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1931),
.B(n_1897),
.Y(n_1947)
);

AOI322xp5_ASAP7_75t_L g1948 ( 
.A1(n_1933),
.A2(n_1932),
.A3(n_1935),
.B1(n_1930),
.B2(n_1929),
.C1(n_1928),
.C2(n_1926),
.Y(n_1948)
);

OAI321xp33_ASAP7_75t_L g1949 ( 
.A1(n_1946),
.A2(n_1933),
.A3(n_1925),
.B1(n_1917),
.B2(n_1873),
.C(n_1879),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1936),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1939),
.B(n_1854),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1939),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1938),
.Y(n_1953)
);

AOI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1946),
.A2(n_1900),
.B1(n_1823),
.B2(n_1810),
.C(n_1809),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1944),
.B(n_1856),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1943),
.B(n_1888),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1941),
.B(n_1773),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1940),
.B(n_1773),
.Y(n_1958)
);

NOR2x1_ASAP7_75t_L g1959 ( 
.A(n_1945),
.B(n_1947),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1952),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1950),
.A2(n_1942),
.B1(n_1937),
.B2(n_1948),
.C(n_1900),
.Y(n_1961)
);

AOI211xp5_ASAP7_75t_L g1962 ( 
.A1(n_1949),
.A2(n_1876),
.B(n_1880),
.C(n_1867),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_R g1963 ( 
.A(n_1951),
.B(n_1629),
.Y(n_1963)
);

AOI222xp33_ASAP7_75t_L g1964 ( 
.A1(n_1954),
.A2(n_1823),
.B1(n_1849),
.B2(n_1810),
.C1(n_1843),
.C2(n_1807),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1959),
.A2(n_1766),
.B(n_1867),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1960),
.Y(n_1966)
);

AOI221x1_ASAP7_75t_L g1967 ( 
.A1(n_1965),
.A2(n_1953),
.B1(n_1958),
.B2(n_1957),
.C(n_1956),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1963),
.Y(n_1968)
);

AOI222xp33_ASAP7_75t_L g1969 ( 
.A1(n_1961),
.A2(n_1839),
.B1(n_1843),
.B2(n_1849),
.C1(n_1955),
.C2(n_1792),
.Y(n_1969)
);

OAI22xp33_ASAP7_75t_L g1970 ( 
.A1(n_1964),
.A2(n_1839),
.B1(n_1780),
.B2(n_1800),
.Y(n_1970)
);

OAI211xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1962),
.A2(n_1800),
.B(n_1759),
.C(n_1838),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1961),
.A2(n_1848),
.B1(n_1841),
.B2(n_1838),
.C(n_1834),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1968),
.B(n_1811),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1969),
.A2(n_1803),
.B1(n_1802),
.B2(n_1848),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1966),
.Y(n_1975)
);

NAND2x1p5_ASAP7_75t_SL g1976 ( 
.A(n_1967),
.B(n_1781),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1972),
.A2(n_1971),
.B1(n_1970),
.B2(n_1802),
.Y(n_1977)
);

NAND2x1_ASAP7_75t_L g1978 ( 
.A(n_1968),
.B(n_1800),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1975),
.B(n_1780),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1976),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1973),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1979),
.B(n_1978),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1982),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1983),
.Y(n_1984)
);

XOR2xp5_ASAP7_75t_L g1985 ( 
.A(n_1983),
.B(n_1980),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1981),
.B1(n_1977),
.B2(n_1974),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1984),
.Y(n_1987)
);

AOI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1987),
.A2(n_1979),
.B1(n_1779),
.B2(n_1792),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1986),
.B(n_1814),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1989),
.A2(n_1815),
.B(n_1814),
.Y(n_1990)
);

OAI22x1_ASAP7_75t_L g1991 ( 
.A1(n_1988),
.A2(n_1781),
.B1(n_1822),
.B2(n_1819),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1990),
.B(n_1815),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1992),
.Y(n_1993)
);

OAI221xp5_ASAP7_75t_R g1994 ( 
.A1(n_1993),
.A2(n_1991),
.B1(n_1781),
.B2(n_1822),
.C(n_1819),
.Y(n_1994)
);

AOI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1598),
.B(n_1699),
.C(n_1824),
.Y(n_1995)
);


endmodule