module fake_jpeg_15644_n_90 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.C(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_54),
.B(n_56),
.Y(n_62)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_17),
.B(n_29),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_16),
.B(n_28),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_35),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_13),
.B(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_33),
.B1(n_39),
.B2(n_5),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_10),
.B(n_11),
.Y(n_70)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_67),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_73),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_12),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_67),
.B1(n_69),
.B2(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_77),
.B(n_80),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_83),
.CI(n_79),
.CON(n_85),
.SN(n_85)
);

AOI322xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_77),
.A3(n_75),
.B1(n_72),
.B2(n_20),
.C1(n_24),
.C2(n_15),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_18),
.B(n_19),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_66),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_25),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_85),
.Y(n_90)
);


endmodule