module real_jpeg_5242_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_0),
.A2(n_162),
.B1(n_166),
.B2(n_169),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_0),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_0),
.B(n_182),
.C(n_186),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_0),
.B(n_92),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_0),
.B(n_142),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_0),
.B(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_1),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_1),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_1),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_1),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_2),
.A2(n_81),
.B1(n_214),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_2),
.A2(n_81),
.B1(n_100),
.B2(n_222),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_2),
.A2(n_81),
.B1(n_381),
.B2(n_458),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_49),
.B1(n_51),
.B2(n_57),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_3),
.A2(n_57),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_57),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_3),
.A2(n_57),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_4),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_4),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_4),
.Y(n_371)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_4),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_4),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_4),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_5),
.A2(n_74),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_5),
.A2(n_74),
.B1(n_222),
.B2(n_406),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_5),
.A2(n_74),
.B1(n_298),
.B2(n_416),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_6),
.Y(n_551)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_193),
.B1(n_198),
.B2(n_199),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_8),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_8),
.A2(n_162),
.B1(n_198),
.B2(n_267),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_8),
.A2(n_198),
.B1(n_378),
.B2(n_380),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_8),
.A2(n_198),
.B1(n_419),
.B2(n_421),
.Y(n_418)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_9),
.Y(n_547)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_12),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_12),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_12),
.A2(n_173),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_12),
.A2(n_173),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_12),
.A2(n_173),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_13),
.Y(n_216)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_15),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_64),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_15),
.A2(n_64),
.B1(n_244),
.B2(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_15),
.A2(n_64),
.B1(n_385),
.B2(n_426),
.Y(n_425)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_17),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_17),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_17),
.A2(n_224),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_17),
.A2(n_224),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_17),
.A2(n_224),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_18),
.A2(n_286),
.B1(n_290),
.B2(n_291),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_18),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_18),
.A2(n_122),
.B1(n_290),
.B2(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_18),
.A2(n_290),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_L g470 ( 
.A1(n_18),
.A2(n_290),
.B1(n_365),
.B2(n_471),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_546),
.B(n_548),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_58),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_47),
.Y(n_23)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_24),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_24),
.B(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_25),
.B(n_169),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_25),
.A2(n_59),
.B1(n_418),
.B2(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_25)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_26),
.Y(n_344)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_28),
.Y(n_281)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_29),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_30),
.Y(n_318)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_31),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_31),
.Y(n_349)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_31),
.Y(n_379)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_31),
.Y(n_382)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_35),
.A2(n_364),
.B(n_368),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_35),
.B(n_370),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_46),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_58)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_53),
.B(n_169),
.Y(n_350)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_58),
.B(n_69),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_65),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_75),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_59),
.A2(n_369),
.B(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_59),
.A2(n_65),
.B1(n_73),
.B2(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_65),
.A2(n_442),
.B(n_472),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_151),
.B(n_545),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_147),
.C(n_148),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_70),
.A2(n_71),
.B1(n_541),
.B2(n_542),
.Y(n_540)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.C(n_116),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_72),
.B(n_533),
.Y(n_532)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_78),
.Y(n_446)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_82),
.A2(n_116),
.B1(n_117),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_82),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_104),
.B1(n_111),
.B2(n_112),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_83),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_83),
.A2(n_111),
.B1(n_316),
.B2(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_83),
.A2(n_111),
.B1(n_412),
.B2(n_415),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_83),
.A2(n_104),
.B1(n_111),
.B2(n_522),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_86),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_88),
.Y(n_413)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_89),
.Y(n_305)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_92),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

AOI22x1_ASAP7_75t_L g447 ( 
.A1(n_92),
.A2(n_149),
.B1(n_320),
.B2(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_92),
.A2(n_149),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

AO22x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_100),
.B2(n_102),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_98),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_99),
.Y(n_299)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_99),
.Y(n_408)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_105),
.Y(n_273)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_111),
.B(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_111),
.A2(n_316),
.B(n_319),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_113),
.Y(n_414)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_116),
.A2(n_117),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_116),
.B(n_517),
.C(n_520),
.Y(n_528)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_141),
.B(n_143),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_161),
.B(n_170),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_118),
.A2(n_141),
.B1(n_221),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_118),
.A2(n_170),
.B(n_266),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_118),
.A2(n_141),
.B1(n_384),
.B2(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_119),
.B(n_171),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_119),
.A2(n_142),
.B1(n_405),
.B2(n_409),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_119),
.A2(n_142),
.B1(n_409),
.B2(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_119),
.A2(n_142),
.B1(n_425),
.B2(n_461),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_130),
.A2(n_221),
.B(n_227),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_137),
.B2(n_139),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_135),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_138),
.Y(n_245)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_138),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_138),
.Y(n_401)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_141),
.A2(n_227),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_143),
.Y(n_461)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_147),
.B(n_148),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_149),
.A2(n_272),
.B(n_278),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_149),
.B(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_149),
.A2(n_278),
.B(n_485),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_539),
.B(n_544),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_511),
.B(n_536),
.Y(n_152)
);

OAI311xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_389),
.A3(n_487),
.B1(n_505),
.C1(n_506),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_334),
.B(n_388),
.Y(n_154)
);

AO21x1_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_307),
.B(n_333),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_260),
.B(n_306),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_230),
.B(n_259),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_190),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_159),
.B(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_176),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_160),
.A2(n_176),
.B1(n_177),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_160),
.Y(n_257)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx5_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_168),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_169),
.A2(n_202),
.B(n_210),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g272 ( 
.A1(n_169),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_SL g364 ( 
.A1(n_169),
.A2(n_350),
.B(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_189),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_218),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_219),
.C(n_229),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_202),
.B(n_210),
.Y(n_191)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_197),
.Y(n_398)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_201),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_202),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_202),
.A2(n_395),
.B1(n_399),
.B2(n_400),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_202),
.A2(n_400),
.B(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_213),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_203),
.A2(n_211),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_203),
.A2(n_285),
.B1(n_324),
.B2(n_330),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_203),
.A2(n_356),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_206),
.Y(n_331)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_206),
.Y(n_439)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_216),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_228),
.B2(n_229),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g303 ( 
.A(n_225),
.B(n_304),
.Y(n_303)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_252),
.B(n_258),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_240),
.B(n_251),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_236),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_238),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_250),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_250),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_248),
.B(n_249),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_284),
.B(n_294),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_262),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_282),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_270),
.B2(n_271),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_270),
.C(n_282),
.Y(n_308)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI32xp33_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_298),
.A3(n_299),
.B1(n_300),
.B2(n_303),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_297),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_308),
.B(n_309),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_314),
.B2(n_332),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_313),
.C(n_332),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_314),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_322),
.C(n_323),
.Y(n_358)
);

OAI32xp33_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_341),
.A3(n_343),
.B1(n_345),
.B2(n_350),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_335),
.B(n_336),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_361),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_351),
.B2(n_352),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_340),
.B(n_351),
.Y(n_483)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx6_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_358),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_358),
.B(n_359),
.C(n_361),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_375),
.B2(n_387),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_362),
.B(n_376),
.C(n_383),
.Y(n_496)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_367),
.Y(n_471)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_383),
.Y(n_375)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_377),
.Y(n_485)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_473),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_390),
.A2(n_473),
.B(n_507),
.C(n_510),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_449),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_391),
.B(n_449),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_422),
.C(n_432),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g486 ( 
.A(n_392),
.B(n_422),
.CI(n_432),
.CON(n_486),
.SN(n_486)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_410),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_393),
.B(n_411),
.C(n_417),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_404),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_394),
.B(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_395),
.Y(n_437)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

INVx4_ASAP7_75t_SL g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_428),
.B2(n_431),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_428),
.Y(n_465)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_428),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_428),
.A2(n_431),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_428),
.A2(n_465),
.B(n_468),
.Y(n_514)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_440),
.C(n_447),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_433),
.B(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_434),
.B(n_436),
.Y(n_495)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_440),
.A2(n_441),
.B1(n_447),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_453),
.C(n_463),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_463),
.B2(n_464),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_459),
.B(n_462),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_460),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_457),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g513 ( 
.A(n_462),
.B(n_514),
.CI(n_515),
.CON(n_513),
.SN(n_513)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_462),
.B(n_514),
.C(n_515),
.Y(n_535)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_486),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_486),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_479),
.C(n_480),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_475),
.A2(n_476),
.B1(n_479),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_482),
.B1(n_484),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_484),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_486),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_500),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_489),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2x1_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_497),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_497),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.C(n_496),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_503),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_496),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_502),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_525),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_524),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_524),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g554 ( 
.A(n_513),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_519),
.B2(n_523),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_516),
.A2(n_517),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_516),
.B(n_527),
.C(n_531),
.Y(n_543)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_519),
.Y(n_523)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_525),
.A2(n_537),
.B(n_538),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_526),
.B(n_535),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_535),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_543),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_543),
.Y(n_544)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_547),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_551),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);


endmodule