module fake_jpeg_7987_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_18),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_30),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_28),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_35),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_30),
.B1(n_20),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_53),
.B1(n_43),
.B2(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_30),
.B1(n_20),
.B2(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_37),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_20),
.B(n_21),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_41),
.B(n_35),
.C(n_21),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_20),
.C(n_22),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_42),
.C(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_43),
.B1(n_39),
.B2(n_26),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_31),
.B1(n_18),
.B2(n_26),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_70),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_41),
.B(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_80),
.Y(n_116)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_109)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_94),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_42),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_95),
.C(n_50),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_31),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_26),
.B1(n_32),
.B2(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_28),
.B1(n_43),
.B2(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_65),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_33),
.B1(n_34),
.B2(n_17),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_33),
.B1(n_17),
.B2(n_40),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_40),
.B1(n_19),
.B2(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_49),
.B(n_19),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_19),
.B1(n_25),
.B2(n_8),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_63),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_64),
.B1(n_65),
.B2(n_22),
.Y(n_124)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_77),
.B1(n_78),
.B2(n_74),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_53),
.B1(n_51),
.B2(n_48),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_46),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_49),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_73),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_95),
.C(n_94),
.Y(n_150)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_11),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_64),
.B1(n_22),
.B2(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_75),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_22),
.B1(n_27),
.B2(n_65),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_83),
.B(n_79),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_103),
.B(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_73),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_128),
.B(n_71),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_79),
.B(n_71),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_76),
.B(n_27),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_144),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_81),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_150),
.Y(n_166)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_118),
.B1(n_102),
.B2(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_85),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_100),
.B(n_97),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_89),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_78),
.B1(n_113),
.B2(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_82),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_164),
.B(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_110),
.B1(n_109),
.B2(n_108),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_178),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_114),
.B(n_103),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_157),
.A2(n_110),
.B1(n_108),
.B2(n_107),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_107),
.B1(n_114),
.B2(n_84),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_107),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_171),
.C(n_129),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_99),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_177),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_137),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_105),
.B1(n_121),
.B2(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_22),
.B1(n_80),
.B2(n_27),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_27),
.B1(n_9),
.B2(n_16),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_134),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_138),
.A2(n_155),
.B1(n_153),
.B2(n_158),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_133),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_156),
.B1(n_141),
.B2(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_204),
.C(n_209),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_134),
.B1(n_136),
.B2(n_132),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_197),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_131),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_131),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_210),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_137),
.B(n_151),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_206),
.B(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_205),
.B1(n_213),
.B2(n_210),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_145),
.C(n_132),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_144),
.B(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_0),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_80),
.CI(n_1),
.CON(n_211),
.SN(n_211)
);

XOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_174),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_183),
.B1(n_189),
.B2(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_9),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_168),
.B1(n_179),
.B2(n_175),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_199),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_185),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_179),
.B1(n_175),
.B2(n_163),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_224),
.B1(n_227),
.B2(n_226),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_160),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_177),
.B1(n_173),
.B2(n_178),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_199),
.B(n_211),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_174),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_235),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_0),
.C(n_2),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_230),
.C(n_196),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_2),
.C(n_3),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_198),
.A2(n_16),
.B1(n_9),
.B2(n_4),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_213),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_7),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_244),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_197),
.B(n_201),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_248),
.B1(n_193),
.B2(n_194),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_206),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_247),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_205),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_252),
.C(n_229),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_217),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_202),
.C(n_195),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_211),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_231),
.B1(n_225),
.B2(n_207),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_257),
.B1(n_253),
.B2(n_243),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_218),
.B1(n_193),
.B2(n_235),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_263),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_267),
.Y(n_271)
);

NAND2x1_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_6),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_12),
.B1(n_14),
.B2(n_4),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_192),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_252),
.B(n_245),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_266),
.B(n_260),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_237),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_256),
.B(n_13),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_275),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_243),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_255),
.B(n_237),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_12),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_12),
.C(n_13),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_258),
.C(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_283),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_276),
.B(n_275),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_286),
.B(n_277),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_259),
.B(n_261),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_256),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_284),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_290),
.A3(n_291),
.B1(n_278),
.B2(n_13),
.C1(n_15),
.C2(n_3),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_271),
.B(n_269),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_281),
.C(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_296),
.C(n_15),
.Y(n_298)
);

HB1xp67_ASAP7_75t_SL g297 ( 
.A(n_294),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_295),
.C(n_2),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_3),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_297),
.Y(n_301)
);


endmodule