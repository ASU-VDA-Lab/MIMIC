module fake_jpeg_11890_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_SL g6 ( 
.A(n_1),
.Y(n_6)
);

INVx2_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_3),
.B(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_10),
.B1(n_11),
.B2(n_7),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_15),
.B1(n_7),
.B2(n_17),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_4),
.B1(n_0),
.B2(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_20),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_11),
.B1(n_7),
.B2(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_13),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_24),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_29),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_27),
.Y(n_34)
);


endmodule