module fake_jpeg_2284_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_4),
.B(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_4),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_65),
.B1(n_55),
.B2(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_61),
.C(n_64),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_64),
.Y(n_105)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_93),
.Y(n_104)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_66),
.B1(n_65),
.B2(n_63),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_55),
.B(n_52),
.C(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_100),
.Y(n_115)
);

INVx2_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_2),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_75),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_104),
.B1(n_31),
.B2(n_47),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_3),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_9),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_123),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_63),
.B1(n_56),
.B2(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_58),
.B1(n_66),
.B2(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_119),
.B1(n_124),
.B2(n_129),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_58),
.B1(n_52),
.B2(n_6),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_128),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_21),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_19),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_111),
.C(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_138),
.C(n_33),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_110),
.C(n_20),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_48),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_152),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_23),
.B(n_25),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_30),
.B(n_32),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_28),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_125),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_163),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_168),
.B(n_147),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_34),
.Y(n_165)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_35),
.B(n_37),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_163),
.C(n_157),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_136),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_141),
.B1(n_166),
.B2(n_135),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_164),
.B1(n_158),
.B2(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_166),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_185)
);

AOI321xp33_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_160),
.A3(n_139),
.B1(n_146),
.B2(n_149),
.C(n_159),
.Y(n_180)
);

AOI211xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_176),
.B(n_152),
.C(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_38),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_187),
.B1(n_41),
.B2(n_42),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_40),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_43),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_44),
.B1(n_46),
.B2(n_185),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_184),
.Y(n_191)
);


endmodule