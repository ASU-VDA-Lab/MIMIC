module fake_netlist_5_1726_n_1104 (n_137, n_210, n_168, n_260, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1104);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1104;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_785;
wire n_316;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_1020;
wire n_798;
wire n_350;
wire n_662;
wire n_459;
wire n_897;
wire n_646;
wire n_1062;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_425;
wire n_513;
wire n_679;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_870;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_985;
wire n_904;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_92),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_158),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_133),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_163),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_97),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_253),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_266),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_84),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_173),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_64),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_65),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_138),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_195),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_243),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_177),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_11),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_46),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_19),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_29),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_67),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_257),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_0),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_87),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_259),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_164),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_217),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_70),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_4),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_178),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_125),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_225),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_200),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_74),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_245),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_53),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_130),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_21),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_201),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_105),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_210),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_55),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_104),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_149),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_229),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_114),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_83),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_42),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_135),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_118),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_235),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_124),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_R g331 ( 
.A(n_296),
.B(n_0),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_267),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_268),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_269),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_268),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_270),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_283),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_283),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_1),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_271),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_293),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_272),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_272),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_293),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_R g371 ( 
.A(n_311),
.B(n_273),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_311),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_369),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_344),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_371),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_338),
.B(n_353),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_286),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_284),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_337),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_361),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_357),
.A2(n_313),
.B(n_299),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_352),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_313),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_370),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_370),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_335),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_275),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_331),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_372),
.A2(n_279),
.B1(n_281),
.B2(n_280),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_358),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_359),
.B(n_277),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_343),
.B(n_277),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_288),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_340),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_339),
.B(n_294),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_345),
.B(n_295),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_347),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_420),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_375),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_382),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_376),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_403),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_351),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_411),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_301),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_401),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_406),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_303),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_304),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_383),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

OAI221xp5_ASAP7_75t_L g450 ( 
.A1(n_398),
.A2(n_317),
.B1(n_329),
.B2(n_328),
.C(n_307),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_310),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_312),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_277),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_380),
.B(n_277),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_315),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_387),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_287),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_392),
.A2(n_319),
.B(n_324),
.C(n_318),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_397),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_381),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_383),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_407),
.B(n_327),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_405),
.B(n_330),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_410),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_405),
.B(n_287),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_416),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_414),
.B(n_287),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_452),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_480),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_487),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_424),
.Y(n_493)
);

NOR3xp33_ASAP7_75t_SL g494 ( 
.A(n_436),
.B(n_400),
.C(n_399),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_379),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_487),
.Y(n_496)
);

AND2x6_ASAP7_75t_SL g497 ( 
.A(n_426),
.B(n_419),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_482),
.Y(n_498)
);

OAI221xp5_ASAP7_75t_L g499 ( 
.A1(n_442),
.A2(n_383),
.B1(n_395),
.B2(n_394),
.C(n_409),
.Y(n_499)
);

CKINVDCx11_ASAP7_75t_R g500 ( 
.A(n_479),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_423),
.B(n_389),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_439),
.B(n_389),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_429),
.B(n_418),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_439),
.B(n_391),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_391),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_452),
.Y(n_506)
);

AO22x1_ASAP7_75t_L g507 ( 
.A1(n_473),
.A2(n_378),
.B1(n_384),
.B2(n_399),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_432),
.B(n_377),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_400),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_447),
.B(n_287),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_473),
.A2(n_351),
.B1(n_364),
.B2(n_418),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_424),
.A2(n_397),
.B1(n_421),
.B2(n_302),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_456),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_456),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_447),
.B(n_302),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_447),
.B(n_459),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_L g519 ( 
.A(n_450),
.B(n_421),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_424),
.A2(n_481),
.B1(n_484),
.B2(n_472),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_427),
.A2(n_302),
.B1(n_422),
.B2(n_416),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_424),
.B(n_302),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_475),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_472),
.Y(n_527)
);

AND2x4_ASAP7_75t_SL g528 ( 
.A(n_479),
.B(n_422),
.Y(n_528)
);

OAI221xp5_ASAP7_75t_L g529 ( 
.A1(n_464),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_427),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_440),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_431),
.B(n_445),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_478),
.B(n_54),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_481),
.B(n_6),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_433),
.B(n_56),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_478),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_458),
.A2(n_58),
.B1(n_59),
.B2(n_57),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_433),
.B(n_60),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_444),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_444),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_448),
.B(n_451),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_469),
.B(n_265),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_445),
.B(n_10),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_448),
.B(n_61),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_451),
.B(n_463),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_453),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_431),
.B(n_434),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_483),
.A2(n_63),
.B(n_62),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_463),
.A2(n_68),
.B(n_66),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_453),
.B(n_12),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_471),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_434),
.B(n_13),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_454),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_454),
.B(n_69),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_455),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_434),
.B(n_14),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_457),
.B(n_71),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_457),
.B(n_14),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_468),
.B(n_72),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_505),
.B(n_479),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_526),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_558),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_457),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_493),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_490),
.B(n_443),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_509),
.B(n_469),
.C(n_462),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_503),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_498),
.B(n_457),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_553),
.A2(n_488),
.B1(n_462),
.B2(n_428),
.Y(n_576)
);

NOR3xp33_ASAP7_75t_SL g577 ( 
.A(n_512),
.B(n_486),
.C(n_485),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_540),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_527),
.B(n_462),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_492),
.B(n_462),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_530),
.B(n_488),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_540),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_521),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_535),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_561),
.B(n_488),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_545),
.Y(n_590)
);

AO22x1_ASAP7_75t_L g591 ( 
.A1(n_554),
.A2(n_510),
.B1(n_553),
.B2(n_491),
.Y(n_591)
);

NOR3xp33_ASAP7_75t_SL g592 ( 
.A(n_512),
.B(n_474),
.C(n_471),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_496),
.B(n_488),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_495),
.Y(n_594)
);

NOR3xp33_ASAP7_75t_SL g595 ( 
.A(n_534),
.B(n_477),
.C(n_474),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_489),
.B(n_477),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_506),
.B(n_449),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_520),
.B(n_455),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_508),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_525),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_518),
.B(n_425),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_522),
.B(n_449),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_525),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_508),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

AND2x6_ASAP7_75t_SL g606 ( 
.A(n_547),
.B(n_15),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_562),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_559),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_531),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_549),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_555),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_557),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_519),
.B(n_425),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_SL g616 ( 
.A(n_499),
.B(n_536),
.C(n_551),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_502),
.B(n_461),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_500),
.B(n_465),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_523),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_538),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_562),
.Y(n_624)
);

BUFx4f_ASAP7_75t_L g625 ( 
.A(n_562),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_539),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_504),
.B(n_428),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_542),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_SL g629 ( 
.A(n_536),
.B(n_470),
.C(n_466),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_615),
.A2(n_563),
.B(n_548),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_601),
.A2(n_552),
.B(n_438),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_587),
.A2(n_514),
.B1(n_546),
.B2(n_543),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_617),
.A2(n_438),
.B(n_430),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_587),
.A2(n_544),
.B1(n_532),
.B2(n_501),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_586),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_574),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_570),
.A2(n_467),
.B(n_455),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_617),
.A2(n_446),
.B(n_430),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_574),
.B(n_528),
.Y(n_640)
);

OAI21x1_ASAP7_75t_SL g641 ( 
.A1(n_573),
.A2(n_624),
.B(n_541),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_587),
.A2(n_494),
.B1(n_529),
.B2(n_556),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_588),
.A2(n_560),
.B1(n_547),
.B2(n_550),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_590),
.B(n_551),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_620),
.A2(n_446),
.B(n_461),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_575),
.A2(n_467),
.B(n_455),
.Y(n_646)
);

AO21x2_ASAP7_75t_L g647 ( 
.A1(n_629),
.A2(n_470),
.B(n_466),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_594),
.A2(n_547),
.B1(n_435),
.B2(n_467),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_614),
.A2(n_467),
.B(n_465),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_623),
.B(n_507),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_620),
.A2(n_465),
.B(n_435),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_619),
.A2(n_467),
.B(n_435),
.Y(n_652)
);

AOI21x1_ASAP7_75t_SL g653 ( 
.A1(n_582),
.A2(n_497),
.B(n_435),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_579),
.B(n_73),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_628),
.A2(n_76),
.B(n_75),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_573),
.B(n_77),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_598),
.A2(n_610),
.B(n_578),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_599),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_627),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_611),
.B(n_612),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_598),
.A2(n_79),
.B(n_78),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_572),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_611),
.B(n_15),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_595),
.A2(n_592),
.B(n_616),
.C(n_612),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_618),
.B(n_16),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_567),
.B(n_16),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_610),
.A2(n_81),
.B(n_80),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_579),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_567),
.A2(n_153),
.B1(n_263),
.B2(n_262),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_578),
.A2(n_85),
.B(n_82),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_608),
.A2(n_88),
.B(n_86),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_567),
.B(n_573),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_591),
.B(n_581),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_585),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_564),
.B(n_17),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_576),
.A2(n_90),
.B(n_89),
.Y(n_676)
);

AO21x1_ASAP7_75t_L g677 ( 
.A1(n_564),
.A2(n_17),
.B(n_18),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_605),
.Y(n_678)
);

NOR2x1_ASAP7_75t_SL g679 ( 
.A(n_600),
.B(n_264),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_577),
.B(n_18),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_613),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_608),
.A2(n_93),
.B(n_91),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_607),
.A2(n_19),
.B(n_20),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_568),
.B(n_20),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_565),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_568),
.B(n_21),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_589),
.Y(n_687)
);

AO31x2_ASAP7_75t_L g688 ( 
.A1(n_628),
.A2(n_22),
.A3(n_23),
.B(n_24),
.Y(n_688)
);

BUFx8_ASAP7_75t_SL g689 ( 
.A(n_599),
.Y(n_689)
);

BUFx4_ASAP7_75t_SL g690 ( 
.A(n_604),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_R g691 ( 
.A1(n_606),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_691)
);

AOI211x1_ASAP7_75t_L g692 ( 
.A1(n_660),
.A2(n_593),
.B(n_566),
.C(n_571),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_678),
.Y(n_693)
);

OA21x2_ASAP7_75t_L g694 ( 
.A1(n_631),
.A2(n_576),
.B(n_605),
.Y(n_694)
);

AOI221xp5_ASAP7_75t_L g695 ( 
.A1(n_643),
.A2(n_624),
.B1(n_625),
.B2(n_627),
.C(n_621),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_657),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_645),
.A2(n_639),
.B(n_633),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_636),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_662),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_674),
.Y(n_700)
);

AOI221x1_ASAP7_75t_L g701 ( 
.A1(n_673),
.A2(n_626),
.B1(n_602),
.B2(n_596),
.C(n_622),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_635),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_672),
.B(n_569),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_672),
.B(n_569),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_659),
.B(n_568),
.Y(n_705)
);

AO21x2_ASAP7_75t_L g706 ( 
.A1(n_652),
.A2(n_584),
.B(n_589),
.Y(n_706)
);

NOR2x1_ASAP7_75t_L g707 ( 
.A(n_644),
.B(n_608),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_661),
.B(n_569),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_681),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_675),
.A2(n_625),
.B1(n_589),
.B2(n_583),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_659),
.B(n_597),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_637),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_664),
.A2(n_626),
.A3(n_625),
.B(n_597),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_636),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_637),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_666),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_685),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_676),
.B(n_626),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_665),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_651),
.A2(n_603),
.B(n_626),
.Y(n_721)
);

AOI221xp5_ASAP7_75t_SL g722 ( 
.A1(n_664),
.A2(n_600),
.B1(n_609),
.B2(n_597),
.C(n_580),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_636),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_583),
.B(n_580),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_650),
.B(n_580),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_684),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_675),
.A2(n_583),
.B1(n_621),
.B2(n_600),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_647),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_652),
.A2(n_649),
.B(n_646),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_687),
.B(n_600),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_647),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_634),
.A2(n_609),
.B1(n_604),
.B2(n_27),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_668),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_649),
.A2(n_609),
.B(n_95),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_642),
.A2(n_609),
.B1(n_26),
.B2(n_27),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_687),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_680),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_663),
.B(n_30),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_638),
.A2(n_96),
.B(n_94),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_689),
.Y(n_740)
);

AO21x2_ASAP7_75t_L g741 ( 
.A1(n_646),
.A2(n_99),
.B(n_98),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_668),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_630),
.A2(n_30),
.B(n_31),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_686),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_689),
.Y(n_745)
);

AOI211xp5_ASAP7_75t_L g746 ( 
.A1(n_732),
.A2(n_683),
.B(n_677),
.C(n_669),
.Y(n_746)
);

AO22x1_ASAP7_75t_L g747 ( 
.A1(n_736),
.A2(n_640),
.B1(n_654),
.B2(n_691),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_737),
.A2(n_656),
.B1(n_655),
.B2(n_641),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_720),
.B(n_654),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_720),
.B(n_648),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_716),
.B(n_656),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_735),
.A2(n_656),
.B1(n_655),
.B2(n_658),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_709),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_SL g754 ( 
.A1(n_719),
.A2(n_679),
.B1(n_658),
.B2(n_682),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_SL g755 ( 
.A1(n_719),
.A2(n_671),
.B1(n_667),
.B2(n_670),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_699),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_726),
.B(n_688),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

CKINVDCx6p67_ASAP7_75t_R g759 ( 
.A(n_733),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_719),
.A2(n_638),
.B1(n_653),
.B2(n_690),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_695),
.B(n_653),
.C(n_690),
.Y(n_761)
);

OAI21xp33_ASAP7_75t_SL g762 ( 
.A1(n_719),
.A2(n_688),
.B(n_101),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_727),
.B(n_688),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_698),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_SL g765 ( 
.A(n_744),
.B(n_688),
.C(n_32),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_719),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_SL g767 ( 
.A(n_710),
.B(n_34),
.C(n_35),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_738),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_700),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_725),
.B(n_36),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_715),
.B(n_100),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_705),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_702),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_SL g774 ( 
.A(n_712),
.B(n_39),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_711),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_700),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_717),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_713),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_724),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_712),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_697),
.A2(n_103),
.B(n_102),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_715),
.B(n_106),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_740),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_717),
.A2(n_741),
.B1(n_693),
.B2(n_707),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_693),
.Y(n_785)
);

OAI211xp5_ASAP7_75t_L g786 ( 
.A1(n_692),
.A2(n_701),
.B(n_739),
.C(n_707),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_701),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_740),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_715),
.B(n_107),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_714),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_714),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_714),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_703),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_741),
.A2(n_743),
.B1(n_703),
.B2(n_704),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_741),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_795)
);

AOI221x1_ASAP7_75t_SL g796 ( 
.A1(n_730),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.C(n_50),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_743),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_703),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_729),
.A2(n_51),
.B(n_52),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_742),
.B(n_108),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_703),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_R g803 ( 
.A(n_745),
.B(n_112),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_698),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_733),
.B(n_113),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_713),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_722),
.A2(n_115),
.B(n_116),
.C(n_117),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_758),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_779),
.A2(n_704),
.B1(n_733),
.B2(n_706),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_756),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_778),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_749),
.B(n_692),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_787),
.A2(n_706),
.B(n_729),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_776),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_779),
.A2(n_743),
.B1(n_704),
.B2(n_731),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_781),
.A2(n_697),
.B(n_734),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_769),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_773),
.B(n_713),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_787),
.A2(n_743),
.B1(n_722),
.B2(n_745),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_757),
.B(n_713),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_767),
.A2(n_731),
.B1(n_728),
.B2(n_698),
.Y(n_822)
);

AO21x2_ASAP7_75t_L g823 ( 
.A1(n_800),
.A2(n_696),
.B(n_728),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_752),
.A2(n_704),
.B1(n_706),
.B2(n_718),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_752),
.A2(n_734),
.B(n_721),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_766),
.A2(n_698),
.B1(n_718),
.B2(n_694),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_764),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_807),
.A2(n_694),
.B(n_721),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_777),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_793),
.B(n_713),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_770),
.B(n_698),
.Y(n_831)
);

OAI221xp5_ASAP7_75t_L g832 ( 
.A1(n_768),
.A2(n_708),
.B1(n_696),
.B2(n_723),
.C(n_694),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_753),
.B(n_694),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_768),
.A2(n_723),
.B1(n_708),
.B2(n_121),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_772),
.A2(n_708),
.B1(n_120),
.B2(n_122),
.Y(n_835)
);

OA21x2_ASAP7_75t_L g836 ( 
.A1(n_784),
.A2(n_119),
.B(n_123),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_796),
.A2(n_775),
.B1(n_772),
.B2(n_795),
.C(n_799),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_838)
);

AOI222xp33_ASAP7_75t_L g839 ( 
.A1(n_747),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.C1(n_136),
.C2(n_139),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_774),
.A2(n_795),
.B1(n_765),
.B2(n_748),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_759),
.Y(n_841)
);

OAI211xp5_ASAP7_75t_L g842 ( 
.A1(n_797),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_842)
);

OAI211xp5_ASAP7_75t_L g843 ( 
.A1(n_797),
.A2(n_143),
.B(n_144),
.C(n_145),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_750),
.A2(n_261),
.B1(n_147),
.B2(n_150),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_761),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_751),
.A2(n_258),
.B1(n_155),
.B2(n_156),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_763),
.A2(n_154),
.B1(n_159),
.B2(n_160),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_760),
.A2(n_161),
.B1(n_162),
.B2(n_165),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_794),
.A2(n_166),
.B(n_167),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_785),
.B(n_168),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_783),
.B(n_169),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_790),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_791),
.Y(n_853)
);

OAI221xp5_ASAP7_75t_L g854 ( 
.A1(n_746),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.C(n_174),
.Y(n_854)
);

OAI211xp5_ASAP7_75t_L g855 ( 
.A1(n_762),
.A2(n_175),
.B(n_176),
.C(n_179),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_789),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_856)
);

AOI222xp33_ASAP7_75t_L g857 ( 
.A1(n_802),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C1(n_187),
.C2(n_188),
.Y(n_857)
);

OAI211xp5_ASAP7_75t_L g858 ( 
.A1(n_803),
.A2(n_189),
.B(n_190),
.C(n_191),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_794),
.A2(n_784),
.B(n_798),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_808),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_837),
.A2(n_754),
.B1(n_771),
.B2(n_782),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_815),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_833),
.Y(n_864)
);

AOI21x1_ASAP7_75t_L g865 ( 
.A1(n_814),
.A2(n_786),
.B(n_806),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_821),
.B(n_778),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_852),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_818),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_840),
.A2(n_771),
.B1(n_782),
.B2(n_806),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_829),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_859),
.B(n_755),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_811),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_811),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_819),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_840),
.A2(n_834),
.B1(n_835),
.B2(n_854),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_812),
.B(n_792),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_853),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_827),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_830),
.B(n_804),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_823),
.B(n_804),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_804),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_820),
.B(n_801),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_817),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_836),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_836),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_825),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_816),
.B(n_804),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_827),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_832),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_849),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_826),
.B(n_764),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_826),
.B(n_764),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_SL g894 ( 
.A1(n_834),
.A2(n_788),
.B1(n_805),
.B2(n_764),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_841),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_831),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_822),
.B(n_805),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_828),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_820),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_816),
.B(n_824),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_850),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_809),
.B(n_193),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_822),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_847),
.B(n_194),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_841),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_855),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_838),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_847),
.B(n_196),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_835),
.B(n_256),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_844),
.B(n_197),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_844),
.B(n_198),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_846),
.B(n_199),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_845),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_860),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_860),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_885),
.A2(n_842),
.B(n_843),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_860),
.Y(n_917)
);

INVxp67_ASAP7_75t_SL g918 ( 
.A(n_873),
.Y(n_918)
);

AOI21xp33_ASAP7_75t_L g919 ( 
.A1(n_883),
.A2(n_839),
.B(n_857),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_867),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_867),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_867),
.Y(n_922)
);

AOI221xp5_ASAP7_75t_L g923 ( 
.A1(n_883),
.A2(n_846),
.B1(n_858),
.B2(n_851),
.C(n_848),
.Y(n_923)
);

AOI222xp33_ASAP7_75t_L g924 ( 
.A1(n_875),
.A2(n_856),
.B1(n_203),
.B2(n_204),
.C1(n_205),
.C2(n_206),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_875),
.A2(n_202),
.B1(n_207),
.B2(n_208),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_909),
.A2(n_209),
.B(n_211),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_866),
.B(n_212),
.Y(n_927)
);

OAI221xp5_ASAP7_75t_L g928 ( 
.A1(n_861),
.A2(n_909),
.B1(n_894),
.B2(n_887),
.C(n_913),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_872),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_866),
.B(n_213),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_907),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_881),
.B(n_218),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_907),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_861),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_862),
.Y(n_935)
);

OAI221xp5_ASAP7_75t_L g936 ( 
.A1(n_909),
.A2(n_227),
.B1(n_228),
.B2(n_231),
.C(n_232),
.Y(n_936)
);

AOI33xp33_ASAP7_75t_L g937 ( 
.A1(n_899),
.A2(n_887),
.A3(n_906),
.B1(n_890),
.B2(n_900),
.B3(n_871),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_868),
.Y(n_938)
);

OA21x2_ASAP7_75t_L g939 ( 
.A1(n_885),
.A2(n_234),
.B(n_236),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_896),
.B(n_237),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_862),
.Y(n_941)
);

OAI31xp33_ASAP7_75t_L g942 ( 
.A1(n_912),
.A2(n_238),
.A3(n_240),
.B(n_242),
.Y(n_942)
);

OAI211xp5_ASAP7_75t_L g943 ( 
.A1(n_903),
.A2(n_244),
.B(n_246),
.C(n_247),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_877),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_907),
.B(n_248),
.C(n_249),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_937),
.B(n_896),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_932),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_914),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_914),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_914),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_929),
.B(n_871),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_915),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_929),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_918),
.B(n_896),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_915),
.B(n_871),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_915),
.B(n_866),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_921),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_921),
.B(n_874),
.Y(n_958)
);

AND2x2_ASAP7_75t_SL g959 ( 
.A(n_939),
.B(n_898),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_935),
.B(n_874),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_940),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_935),
.B(n_863),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_921),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_941),
.B(n_863),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_920),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_917),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_944),
.B(n_864),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_941),
.B(n_863),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_919),
.A2(n_894),
.B1(n_911),
.B2(n_910),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_917),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_944),
.B(n_890),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_949),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_966),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_SL g974 ( 
.A1(n_959),
.A2(n_903),
.B(n_942),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_966),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_970),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_970),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_960),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_949),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_954),
.B(n_922),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_969),
.A2(n_926),
.B(n_942),
.C(n_928),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_949),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_971),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_946),
.B(n_890),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_955),
.B(n_920),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_949),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_956),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_957),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_955),
.B(n_938),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_961),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_987),
.B(n_951),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_973),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_951),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_981),
.B(n_926),
.C(n_945),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_978),
.B(n_962),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_985),
.B(n_947),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_980),
.B(n_964),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_972),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_989),
.B(n_947),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_989),
.B(n_947),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_983),
.B(n_947),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_994),
.A2(n_974),
.B1(n_981),
.B2(n_959),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_992),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_997),
.B(n_968),
.Y(n_1004)
);

OAI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_994),
.A2(n_898),
.B1(n_899),
.B2(n_945),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_996),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_995),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_990),
.B(n_958),
.Y(n_1008)
);

OAI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_990),
.A2(n_923),
.B1(n_936),
.B2(n_925),
.C(n_924),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_959),
.C(n_943),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1005),
.A2(n_1001),
.B(n_934),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_SL g1012 ( 
.A1(n_1009),
.A2(n_895),
.B(n_939),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1003),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1007),
.B(n_993),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1013),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1014),
.B(n_1006),
.Y(n_1016)
);

XNOR2xp5_ASAP7_75t_L g1017 ( 
.A(n_1010),
.B(n_1011),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1012),
.B(n_1008),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1014),
.B(n_999),
.Y(n_1019)
);

OAI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1018),
.A2(n_1004),
.B1(n_988),
.B2(n_895),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1016),
.B(n_991),
.Y(n_1021)
);

NOR4xp25_ASAP7_75t_L g1022 ( 
.A(n_1015),
.B(n_1018),
.C(n_1017),
.D(n_1019),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_1000),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_SL g1024 ( 
.A1(n_1017),
.A2(n_912),
.B(n_911),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1017),
.A2(n_988),
.B1(n_895),
.B2(n_953),
.Y(n_1025)
);

AOI211x1_ASAP7_75t_L g1026 ( 
.A1(n_1018),
.A2(n_975),
.B(n_976),
.C(n_977),
.Y(n_1026)
);

AOI211xp5_ASAP7_75t_L g1027 ( 
.A1(n_1022),
.A2(n_912),
.B(n_910),
.C(n_911),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1021),
.B(n_998),
.Y(n_1028)
);

AOI321xp33_ASAP7_75t_L g1029 ( 
.A1(n_1020),
.A2(n_910),
.A3(n_908),
.B1(n_904),
.B2(n_902),
.C(n_932),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1025),
.B(n_998),
.Y(n_1030)
);

NOR2x1_ASAP7_75t_L g1031 ( 
.A(n_1024),
.B(n_939),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1026),
.B(n_972),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_1030),
.B(n_1031),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1029),
.B(n_1023),
.Y(n_1034)
);

OAI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1028),
.A2(n_913),
.B1(n_905),
.B2(n_979),
.Y(n_1035)
);

OAI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1032),
.A2(n_905),
.B1(n_913),
.B2(n_931),
.C(n_933),
.Y(n_1036)
);

XNOR2x1_ASAP7_75t_L g1037 ( 
.A(n_1028),
.B(n_908),
.Y(n_1037)
);

AOI311xp33_ASAP7_75t_L g1038 ( 
.A1(n_1027),
.A2(n_906),
.A3(n_948),
.B(n_952),
.C(n_963),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1027),
.A2(n_905),
.B1(n_932),
.B2(n_904),
.Y(n_1039)
);

AOI221xp5_ASAP7_75t_L g1040 ( 
.A1(n_1027),
.A2(n_904),
.B1(n_908),
.B2(n_902),
.C(n_932),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1037),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1034),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1033),
.A2(n_939),
.B(n_902),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1039),
.B(n_986),
.Y(n_1044)
);

AOI211xp5_ASAP7_75t_SL g1045 ( 
.A1(n_1035),
.A2(n_927),
.B(n_930),
.C(n_869),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_1038),
.B(n_927),
.C(n_930),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1036),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_1040),
.A2(n_869),
.B1(n_897),
.B2(n_900),
.C(n_986),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_1034),
.B(n_982),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_1034),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_1034),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_1033),
.B(n_897),
.C(n_876),
.Y(n_1052)
);

NAND4xp75_ASAP7_75t_L g1053 ( 
.A(n_1033),
.B(n_916),
.C(n_958),
.D(n_979),
.Y(n_1053)
);

CKINVDCx6p67_ASAP7_75t_R g1054 ( 
.A(n_1034),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_1034),
.B(n_901),
.C(n_876),
.Y(n_1055)
);

NAND4xp25_ASAP7_75t_L g1056 ( 
.A(n_1042),
.B(n_900),
.C(n_901),
.D(n_888),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_1049),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1054),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_1051),
.B(n_982),
.C(n_901),
.Y(n_1059)
);

AOI211xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1047),
.A2(n_893),
.B(n_892),
.C(n_873),
.Y(n_1060)
);

OAI211xp5_ASAP7_75t_SL g1061 ( 
.A1(n_1041),
.A2(n_893),
.B(n_892),
.C(n_878),
.Y(n_1061)
);

AOI222xp33_ASAP7_75t_L g1062 ( 
.A1(n_1050),
.A2(n_1048),
.B1(n_1046),
.B2(n_1043),
.C1(n_1055),
.C2(n_1052),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_1044),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1046),
.B(n_965),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_L g1065 ( 
.A(n_1053),
.B(n_891),
.C(n_878),
.Y(n_1065)
);

NAND5xp2_ASAP7_75t_L g1066 ( 
.A(n_1045),
.B(n_888),
.C(n_865),
.D(n_881),
.E(n_882),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1042),
.A2(n_965),
.B1(n_957),
.B2(n_950),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_L g1068 ( 
.A(n_1042),
.B(n_891),
.C(n_889),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1054),
.B(n_956),
.Y(n_1069)
);

NOR4xp25_ASAP7_75t_L g1070 ( 
.A(n_1042),
.B(n_963),
.C(n_952),
.D(n_948),
.Y(n_1070)
);

OAI211xp5_ASAP7_75t_SL g1071 ( 
.A1(n_1042),
.A2(n_892),
.B(n_893),
.C(n_891),
.Y(n_1071)
);

OAI311xp33_ASAP7_75t_L g1072 ( 
.A1(n_1049),
.A2(n_967),
.A3(n_880),
.B1(n_888),
.C1(n_882),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_1057),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1058),
.A2(n_886),
.B1(n_965),
.B2(n_950),
.C(n_889),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1069),
.B(n_967),
.Y(n_1075)
);

CKINVDCx16_ASAP7_75t_R g1076 ( 
.A(n_1059),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1063),
.B(n_916),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1067),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1056),
.B(n_916),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_1070),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_1062),
.B(n_916),
.C(n_889),
.Y(n_1081)
);

NOR4xp25_ASAP7_75t_L g1082 ( 
.A(n_1071),
.B(n_922),
.C(n_886),
.D(n_868),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1073),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1080),
.Y(n_1084)
);

XNOR2xp5_ASAP7_75t_L g1085 ( 
.A(n_1078),
.B(n_1068),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1076),
.Y(n_1086)
);

OR3x2_ASAP7_75t_L g1087 ( 
.A(n_1081),
.B(n_1066),
.C(n_1060),
.Y(n_1087)
);

AO22x1_ASAP7_75t_L g1088 ( 
.A1(n_1077),
.A2(n_1065),
.B1(n_1064),
.B2(n_1072),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1075),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1086),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1087),
.A2(n_1079),
.B1(n_1074),
.B2(n_1061),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_1084),
.A2(n_1082),
.B(n_938),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_1085),
.A2(n_886),
.B(n_884),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1090),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_1091),
.Y(n_1095)
);

AOI221xp5_ASAP7_75t_L g1096 ( 
.A1(n_1094),
.A2(n_1083),
.B1(n_1088),
.B2(n_1089),
.C(n_1092),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1095),
.A2(n_1093),
.B(n_884),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1094),
.A2(n_879),
.B(n_868),
.C(n_870),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_SL g1099 ( 
.A1(n_1097),
.A2(n_879),
.B1(n_881),
.B2(n_882),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_SL g1100 ( 
.A1(n_1096),
.A2(n_879),
.B1(n_872),
.B2(n_870),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1100),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1102),
.A2(n_1101),
.B1(n_1098),
.B2(n_870),
.C(n_884),
.Y(n_1103)
);

AOI211xp5_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_250),
.B(n_251),
.C(n_252),
.Y(n_1104)
);


endmodule