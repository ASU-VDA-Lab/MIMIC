module fake_jpeg_10192_n_193 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_193);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_31),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_23),
.B1(n_24),
.B2(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_44),
.B1(n_18),
.B2(n_12),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_23),
.B1(n_12),
.B2(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_18),
.B1(n_6),
.B2(n_11),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_53),
.B1(n_6),
.B2(n_11),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_34),
.B1(n_38),
.B2(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_11),
.B(n_10),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_5),
.B1(n_7),
.B2(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_37),
.B1(n_35),
.B2(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_12),
.B1(n_22),
.B2(n_13),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_59),
.B1(n_63),
.B2(n_27),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_43),
.B1(n_44),
.B2(n_19),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_42),
.B1(n_33),
.B2(n_32),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_27),
.B(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_89),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_64),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_98),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_55),
.A3(n_59),
.B1(n_49),
.B2(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_51),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_69),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_65),
.Y(n_106)
);

NOR2x1_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_89),
.C(n_84),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_93),
.C(n_90),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_114),
.B(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_111),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_66),
.B1(n_81),
.B2(n_76),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_76),
.B1(n_68),
.B2(n_96),
.Y(n_124)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_74),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_132),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_90),
.B1(n_87),
.B2(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_104),
.B1(n_110),
.B2(n_105),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_125),
.C(n_128),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_93),
.B(n_86),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_130),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_86),
.C(n_71),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_70),
.C(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

XOR2x1_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_95),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_75),
.B(n_2),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_100),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_145),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_140),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_115),
.B1(n_108),
.B2(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_115),
.B1(n_107),
.B2(n_110),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_143),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_152),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_122),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_153),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_123),
.C(n_131),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_128),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_99),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_135),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_136),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_162),
.C(n_111),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_133),
.B(n_121),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_132),
.C(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_105),
.B1(n_118),
.B2(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_166),
.B1(n_7),
.B2(n_3),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_111),
.B1(n_60),
.B2(n_3),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_155),
.B(n_149),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_170),
.B1(n_159),
.B2(n_158),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_148),
.B(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_158),
.C(n_30),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_3),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_178),
.C(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_1),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_30),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_30),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_180),
.B(n_183),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_167),
.B(n_27),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_60),
.B1(n_58),
.B2(n_2),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_179),
.Y(n_185)
);

AOI21x1_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_182),
.B(n_1),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_182),
.B(n_2),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_189),
.B(n_187),
.C(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_1),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_27),
.Y(n_193)
);


endmodule