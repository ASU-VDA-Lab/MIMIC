module fake_netlist_6_868_n_789 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_789);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_789;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_772;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_719;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_49),
.Y(n_147)
);

BUFx10_ASAP7_75t_L g148 ( 
.A(n_19),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_14),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_32),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_31),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_28),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_107),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_23),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_73),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_56),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_54),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_88),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_97),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_3),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_48),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_55),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_70),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_46),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_71),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_106),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_34),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_115),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_36),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_66),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_2),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_138),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_7),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_30),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_42),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_67),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_68),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_38),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_25),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_146),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_149),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_179),
.B(n_0),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_148),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_0),
.Y(n_215)
);

CKINVDCx6p67_ASAP7_75t_R g216 ( 
.A(n_160),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_1),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_1),
.B(n_2),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_162),
.B(n_3),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_16),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

OAI22x1_ASAP7_75t_SL g230 ( 
.A1(n_166),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_17),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_190),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_157),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g239 ( 
.A(n_152),
.B(n_18),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_20),
.Y(n_241)
);

BUFx8_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_163),
.B(n_21),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_164),
.Y(n_244)
);

BUFx8_ASAP7_75t_SL g245 ( 
.A(n_165),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_203),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_203),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_R g254 ( 
.A(n_238),
.B(n_168),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_212),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_205),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_242),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_236),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_236),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_172),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_173),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_237),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_219),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_219),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_219),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_238),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_234),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_234),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_240),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_214),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_240),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_244),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_202),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_246),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_246),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_214),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_214),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_227),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_211),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_241),
.Y(n_304)
);

BUFx8_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_267),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_241),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_241),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_243),
.Y(n_310)
);

OR2x6_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_225),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_225),
.B(n_227),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_295),
.B(n_243),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_243),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_226),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_276),
.B(n_211),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_286),
.Y(n_321)
);

BUFx6f_ASAP7_75t_SL g322 ( 
.A(n_283),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_286),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_262),
.A2(n_231),
.B(n_227),
.C(n_218),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_278),
.B(n_226),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_265),
.B(n_231),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_279),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_266),
.B(n_231),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_254),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_269),
.B(n_223),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_273),
.B(n_232),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_223),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_281),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g336 ( 
.A(n_274),
.B(n_215),
.C(n_208),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_233),
.C(n_207),
.Y(n_337)
);

NAND2x1_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_239),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_283),
.B(n_175),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_232),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_294),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_207),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_259),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_257),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_261),
.B(n_239),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_263),
.B(n_208),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_253),
.B(n_223),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_247),
.B(n_228),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_250),
.B(n_177),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_252),
.B(n_204),
.Y(n_354)
);

BUFx8_ASAP7_75t_L g355 ( 
.A(n_255),
.Y(n_355)
);

AOI221xp5_ASAP7_75t_L g356 ( 
.A1(n_262),
.A2(n_230),
.B1(n_204),
.B2(n_228),
.C(n_187),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_287),
.B(n_178),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_258),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_248),
.B(n_228),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_260),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_300),
.B(n_182),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

AOI22x1_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_239),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_239),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_239),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_300),
.A2(n_239),
.B1(n_201),
.B2(n_199),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_222),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_304),
.B(n_185),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_316),
.B(n_206),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_311),
.A2(n_229),
.B1(n_224),
.B2(n_222),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_224),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_320),
.B(n_189),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_193),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_224),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

AOI21x1_ASAP7_75t_L g381 ( 
.A1(n_299),
.A2(n_209),
.B(n_210),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_327),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_302),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_334),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_327),
.B(n_224),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_329),
.A2(n_310),
.B1(n_313),
.B2(n_314),
.Y(n_389)
);

AND2x6_ASAP7_75t_SL g390 ( 
.A(n_354),
.B(n_4),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_332),
.B(n_194),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_328),
.B(n_195),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_303),
.B(n_196),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_347),
.B(n_197),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_329),
.A2(n_198),
.B1(n_224),
.B2(n_229),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_299),
.B(n_229),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_349),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

NOR3xp33_ASAP7_75t_SL g401 ( 
.A(n_356),
.B(n_5),
.C(n_6),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_349),
.B(n_229),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_343),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_229),
.B1(n_220),
.B2(n_217),
.Y(n_404)
);

BUFx12f_ASAP7_75t_L g405 ( 
.A(n_305),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_297),
.Y(n_406)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_220),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_309),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_326),
.B(n_350),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_312),
.B(n_217),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_361),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_SL g416 ( 
.A(n_336),
.B(n_8),
.C(n_9),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_337),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_321),
.B(n_22),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_311),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_301),
.Y(n_420)
);

AND2x6_ASAP7_75t_SL g421 ( 
.A(n_348),
.B(n_11),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_301),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_306),
.B(n_24),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_339),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_312),
.B(n_26),
.Y(n_425)
);

NAND2x1p5_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_27),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_12),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_346),
.B(n_13),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_351),
.B(n_14),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_R g430 ( 
.A(n_322),
.B(n_305),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

O2A1O1Ixp5_ASAP7_75t_SL g432 ( 
.A1(n_402),
.A2(n_311),
.B(n_318),
.C(n_315),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_353),
.B(n_361),
.Y(n_433)
);

O2A1O1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_15),
.B(n_361),
.C(n_301),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_15),
.B(n_29),
.C(n_33),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_35),
.B(n_37),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_387),
.A2(n_39),
.B(n_40),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

AO21x2_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_41),
.B(n_43),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_412),
.Y(n_441)
);

BUFx12f_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_397),
.B(n_355),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_400),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_355),
.B1(n_45),
.B2(n_47),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_44),
.C(n_50),
.Y(n_447)
);

INVx8_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_363),
.B(n_51),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_386),
.Y(n_450)
);

NOR3xp33_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_52),
.C(n_53),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_372),
.A2(n_57),
.B(n_59),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

O2A1O1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_417),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_382),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_458)
);

O2A1O1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_403),
.A2(n_69),
.B(n_72),
.C(n_75),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_76),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_374),
.B(n_77),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_393),
.B(n_78),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_376),
.A2(n_79),
.B(n_80),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_388),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_368),
.B(n_86),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_389),
.B(n_87),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_415),
.Y(n_469)
);

NAND2x1p5_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_89),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_362),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_422),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_409),
.B(n_429),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_379),
.B(n_90),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_414),
.B(n_92),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_409),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_377),
.B(n_93),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_413),
.A2(n_94),
.B(n_95),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_430),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_98),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_371),
.B(n_99),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_375),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_487)
);

CKINVDCx8_ASAP7_75t_R g488 ( 
.A(n_390),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_396),
.B(n_105),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_391),
.B(n_109),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_438),
.Y(n_491)
);

AOI22x1_ASAP7_75t_L g492 ( 
.A1(n_433),
.A2(n_426),
.B1(n_431),
.B2(n_369),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_475),
.Y(n_493)
);

AO21x2_ASAP7_75t_L g494 ( 
.A1(n_433),
.A2(n_425),
.B(n_413),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_439),
.B(n_409),
.Y(n_495)
);

OAI21x1_ASAP7_75t_SL g496 ( 
.A1(n_457),
.A2(n_423),
.B(n_418),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_401),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_461),
.A2(n_370),
.B(n_394),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_448),
.Y(n_499)
);

AO21x2_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_489),
.B(n_484),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_432),
.A2(n_426),
.B(n_367),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_486),
.A2(n_404),
.B(n_395),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_392),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_445),
.B(n_429),
.Y(n_506)
);

BUFx2_ASAP7_75t_SL g507 ( 
.A(n_450),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_448),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_444),
.B(n_364),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

BUFx12f_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

AOI22x1_ASAP7_75t_L g512 ( 
.A1(n_481),
.A2(n_394),
.B1(n_373),
.B2(n_378),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_463),
.B(n_428),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_477),
.A2(n_112),
.B(n_113),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_114),
.Y(n_516)
);

AOI21x1_ASAP7_75t_L g517 ( 
.A1(n_480),
.A2(n_449),
.B(n_485),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_453),
.Y(n_518)
);

INVx8_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_490),
.A2(n_116),
.B(n_117),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_482),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_456),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_454),
.B(n_472),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_476),
.B(n_462),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_118),
.Y(n_527)
);

BUFx2_ASAP7_75t_SL g528 ( 
.A(n_479),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_460),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_434),
.A2(n_120),
.B(n_121),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_483),
.Y(n_532)
);

OA21x2_ASAP7_75t_L g533 ( 
.A1(n_435),
.A2(n_436),
.B(n_437),
.Y(n_533)
);

AOI22x1_ASAP7_75t_L g534 ( 
.A1(n_454),
.A2(n_421),
.B1(n_123),
.B2(n_124),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_472),
.Y(n_535)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_452),
.A2(n_122),
.B(n_125),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_465),
.A2(n_127),
.B(n_128),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_510),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_515),
.Y(n_539)
);

AO21x1_ASAP7_75t_L g540 ( 
.A1(n_513),
.A2(n_487),
.B(n_459),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_498),
.A2(n_517),
.B(n_496),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_505),
.Y(n_542)
);

AOI21x1_ASAP7_75t_L g543 ( 
.A1(n_496),
.A2(n_487),
.B(n_446),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_505),
.Y(n_544)
);

OA21x2_ASAP7_75t_L g545 ( 
.A1(n_502),
.A2(n_451),
.B(n_458),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_501),
.Y(n_546)
);

AO21x1_ASAP7_75t_SL g547 ( 
.A1(n_522),
.A2(n_458),
.B(n_466),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_518),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_491),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_493),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_521),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_491),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

BUFx8_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_497),
.B(n_506),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_535),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_535),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_493),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_524),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_446),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_502),
.A2(n_478),
.B(n_470),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_506),
.B(n_469),
.Y(n_562)
);

CKINVDCx11_ASAP7_75t_R g563 ( 
.A(n_511),
.Y(n_563)
);

INVx6_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_497),
.A2(n_447),
.B1(n_483),
.B2(n_443),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_492),
.A2(n_467),
.B(n_440),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_494),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_494),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_503),
.Y(n_570)
);

AO21x1_ASAP7_75t_SL g571 ( 
.A1(n_504),
.A2(n_130),
.B(n_132),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_495),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_495),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_495),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g575 ( 
.A(n_523),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

BUFx2_ASAP7_75t_SL g577 ( 
.A(n_501),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_525),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_576),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_555),
.B(n_527),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_R g581 ( 
.A(n_560),
.B(n_520),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_564),
.Y(n_582)
);

OR2x2_ASAP7_75t_SL g583 ( 
.A(n_558),
.B(n_499),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_575),
.B(n_523),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_576),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_547),
.A2(n_534),
.B1(n_516),
.B2(n_529),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_559),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_538),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_541),
.A2(n_537),
.B(n_514),
.Y(n_589)
);

AO32x2_ASAP7_75t_L g590 ( 
.A1(n_550),
.A2(n_531),
.A3(n_530),
.B1(n_514),
.B2(n_533),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_555),
.B(n_528),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_542),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_539),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_550),
.B(n_499),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_549),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_547),
.A2(n_516),
.B1(n_529),
.B2(n_512),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g597 ( 
.A1(n_567),
.A2(n_541),
.B(n_570),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_544),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_563),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_559),
.B(n_499),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_542),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_499),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_553),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_562),
.A2(n_516),
.B1(n_519),
.B2(n_488),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_553),
.B(n_531),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_575),
.B(n_508),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_519),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_554),
.A2(n_516),
.B1(n_531),
.B2(n_507),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_R g609 ( 
.A(n_563),
.B(n_508),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_527),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_564),
.Y(n_612)
);

CKINVDCx8_ASAP7_75t_R g613 ( 
.A(n_577),
.Y(n_613)
);

NOR3xp33_ASAP7_75t_SL g614 ( 
.A(n_574),
.B(n_578),
.C(n_551),
.Y(n_614)
);

CKINVDCx11_ASAP7_75t_R g615 ( 
.A(n_554),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_546),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_565),
.B(n_526),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_557),
.B(n_526),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_554),
.Y(n_623)
);

AND2x4_ASAP7_75t_SL g624 ( 
.A(n_546),
.B(n_508),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_566),
.Y(n_627)
);

INVxp33_ASAP7_75t_SL g628 ( 
.A(n_568),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_588),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_519),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_625),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_569),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_595),
.B(n_519),
.Y(n_633)
);

NAND2x1_ASAP7_75t_L g634 ( 
.A(n_614),
.B(n_546),
.Y(n_634)
);

BUFx2_ASAP7_75t_SL g635 ( 
.A(n_613),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_627),
.B(n_569),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_621),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_593),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_619),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_598),
.B(n_568),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_579),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_592),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_612),
.B(n_508),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_605),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_579),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_585),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_587),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_585),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_590),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_605),
.B(n_571),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_620),
.B(n_571),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_595),
.B(n_526),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_545),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_603),
.B(n_545),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_591),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_611),
.B(n_545),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_597),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_610),
.B(n_618),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_612),
.B(n_501),
.Y(n_659)
);

OA21x2_ASAP7_75t_L g660 ( 
.A1(n_589),
.A2(n_567),
.B(n_543),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_590),
.B(n_530),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_582),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_590),
.Y(n_663)
);

INVx4_ASAP7_75t_R g664 ( 
.A(n_615),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_616),
.B(n_532),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_586),
.A2(n_533),
.B1(n_532),
.B2(n_524),
.C(n_536),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_587),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_597),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_614),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_656),
.B(n_608),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_656),
.B(n_608),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_655),
.B(n_628),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_644),
.B(n_596),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_641),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_644),
.B(n_530),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_650),
.B(n_622),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_631),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_648),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_669),
.A2(n_604),
.B1(n_540),
.B2(n_602),
.C(n_584),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_658),
.B(n_583),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_646),
.B(n_607),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_645),
.B(n_622),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_665),
.B(n_582),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_638),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_649),
.B(n_663),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_631),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_639),
.B(n_587),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_668),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_640),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_640),
.Y(n_693)
);

AOI211xp5_ASAP7_75t_L g694 ( 
.A1(n_666),
.A2(n_540),
.B(n_606),
.C(n_609),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_650),
.B(n_561),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_637),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_674),
.B(n_632),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_680),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_685),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_678),
.B(n_661),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_679),
.A2(n_581),
.B1(n_651),
.B2(n_635),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_670),
.B(n_661),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_691),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_676),
.B(n_651),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_696),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_694),
.B(n_633),
.C(n_652),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_676),
.B(n_653),
.Y(n_707)
);

BUFx12f_ASAP7_75t_L g708 ( 
.A(n_681),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_670),
.B(n_649),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_677),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_671),
.B(n_654),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_677),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_698),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_700),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_710),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_699),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_701),
.A2(n_708),
.B1(n_706),
.B2(n_673),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_712),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_711),
.B(n_673),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_708),
.A2(n_671),
.B1(n_635),
.B2(n_695),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_705),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_704),
.B(n_686),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_703),
.Y(n_723)
);

XOR2xp5_ASAP7_75t_L g724 ( 
.A(n_717),
.B(n_599),
.Y(n_724)
);

NOR2x1_ASAP7_75t_L g725 ( 
.A(n_721),
.B(n_684),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_718),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_L g727 ( 
.A1(n_720),
.A2(n_697),
.B(n_690),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_L g728 ( 
.A1(n_713),
.A2(n_672),
.B1(n_709),
.B2(n_697),
.C(n_683),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_716),
.B(n_682),
.C(n_695),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_724),
.A2(n_722),
.B1(n_719),
.B2(n_714),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_725),
.A2(n_634),
.B(n_714),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_727),
.B(n_709),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_726),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_729),
.A2(n_722),
.B1(n_702),
.B2(n_634),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_L g735 ( 
.A1(n_728),
.A2(n_715),
.B(n_723),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_733),
.Y(n_736)
);

XOR2x2_ASAP7_75t_L g737 ( 
.A(n_730),
.B(n_664),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_734),
.B(n_630),
.C(n_667),
.Y(n_738)
);

OAI21xp33_ASAP7_75t_SL g739 ( 
.A1(n_732),
.A2(n_702),
.B(n_707),
.Y(n_739)
);

AOI31xp33_ASAP7_75t_L g740 ( 
.A1(n_738),
.A2(n_623),
.A3(n_731),
.B(n_735),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_736),
.B(n_667),
.C(n_617),
.Y(n_741)
);

AOI221xp5_ASAP7_75t_L g742 ( 
.A1(n_740),
.A2(n_739),
.B1(n_737),
.B2(n_703),
.C(n_693),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_741),
.A2(n_647),
.B(n_594),
.C(n_600),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_740),
.B(n_501),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_744),
.B(n_647),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_643),
.B1(n_600),
.B2(n_662),
.Y(n_746)
);

INVx5_ASAP7_75t_L g747 ( 
.A(n_743),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_744),
.B(n_643),
.Y(n_748)
);

AND3x4_ASAP7_75t_L g749 ( 
.A(n_744),
.B(n_643),
.C(n_594),
.Y(n_749)
);

NOR2x1_ASAP7_75t_L g750 ( 
.A(n_744),
.B(n_662),
.Y(n_750)
);

NAND4xp75_ASAP7_75t_L g751 ( 
.A(n_750),
.B(n_533),
.C(n_675),
.D(n_692),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_745),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_749),
.B(n_662),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_747),
.B(n_662),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_L g755 ( 
.A1(n_746),
.A2(n_662),
.B1(n_688),
.B2(n_689),
.C(n_687),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_748),
.B(n_688),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_747),
.B(n_687),
.Y(n_757)
);

NOR2x1_ASAP7_75t_L g758 ( 
.A(n_754),
.B(n_602),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_752),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_757),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_753),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_756),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_755),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_759),
.A2(n_751),
.B1(n_659),
.B2(n_624),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

NOR2x2_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_689),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_760),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_763),
.A2(n_659),
.B1(n_687),
.B2(n_564),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_758),
.Y(n_769)
);

OA22x2_ASAP7_75t_L g770 ( 
.A1(n_761),
.A2(n_659),
.B1(n_642),
.B2(n_691),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_759),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_766),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_771),
.A2(n_663),
.B1(n_657),
.B2(n_642),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_765),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_764),
.A2(n_657),
.B1(n_636),
.B2(n_668),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_767),
.A2(n_675),
.B1(n_654),
.B2(n_653),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_769),
.A2(n_660),
.B1(n_537),
.B2(n_632),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_768),
.A2(n_636),
.B1(n_660),
.B2(n_525),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_770),
.A2(n_660),
.B1(n_536),
.B2(n_135),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_774),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_772),
.B(n_133),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_775),
.Y(n_782)
);

XOR2x2_ASAP7_75t_L g783 ( 
.A(n_779),
.B(n_134),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_783),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_780),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_781),
.B(n_782),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_SL g787 ( 
.A1(n_786),
.A2(n_784),
.B1(n_773),
.B2(n_778),
.Y(n_787)
);

AOI221x1_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_777),
.B1(n_776),
.B2(n_139),
.C(n_141),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_500),
.B1(n_561),
.B2(n_503),
.Y(n_789)
);


endmodule