module fake_jpeg_26466_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_45),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_33),
.B(n_19),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_42),
.Y(n_65)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_23),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_61),
.B(n_62),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_41),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_64),
.B1(n_43),
.B2(n_37),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_40),
.B1(n_29),
.B2(n_33),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_65),
.A2(n_27),
.B1(n_32),
.B2(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_84),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_19),
.B1(n_21),
.B2(n_24),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_68),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_73),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_92),
.B1(n_101),
.B2(n_59),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_75),
.Y(n_125)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_59),
.B1(n_51),
.B2(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_39),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_91),
.C(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_39),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_43),
.B1(n_36),
.B2(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_52),
.B(n_29),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_25),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_43),
.B1(n_20),
.B2(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_18),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_42),
.C(n_2),
.Y(n_129)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_20),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_73),
.B1(n_94),
.B2(n_87),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_129),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_115),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_59),
.B1(n_51),
.B2(n_28),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_22),
.B1(n_42),
.B2(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_22),
.B1(n_42),
.B2(n_17),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_130),
.B1(n_86),
.B2(n_97),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_77),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_103),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_134),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_88),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_90),
.B(n_80),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_139),
.B(n_117),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_75),
.B1(n_81),
.B2(n_100),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_153),
.B1(n_108),
.B2(n_104),
.Y(n_176)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_69),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_151),
.B1(n_156),
.B2(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_72),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_70),
.Y(n_149)
);

XOR2x2_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_120),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_102),
.B1(n_92),
.B2(n_11),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_101),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_142),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_0),
.Y(n_159)
);

XNOR2x2_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_8),
.C(n_14),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_130),
.C(n_129),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_105),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_168),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_119),
.B1(n_125),
.B2(n_109),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_187),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_126),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_179),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_132),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_185),
.B(n_191),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_142),
.A2(n_111),
.B1(n_105),
.B2(n_9),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_179),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_111),
.B1(n_4),
.B2(n_5),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_197),
.B1(n_148),
.B2(n_160),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_133),
.A2(n_0),
.B(n_4),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_5),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_133),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_156),
.B1(n_151),
.B2(n_158),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_187),
.B1(n_177),
.B2(n_169),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_197)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_149),
.A3(n_144),
.B1(n_145),
.B2(n_134),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_199),
.B(n_220),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_222),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_196),
.B1(n_165),
.B2(n_180),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_172),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_217),
.B1(n_152),
.B2(n_157),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_215),
.B1(n_171),
.B2(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_214),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_182),
.B(n_162),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_166),
.B(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_164),
.A2(n_148),
.B1(n_135),
.B2(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_174),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_188),
.B(n_171),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_135),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_135),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_188),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_157),
.Y(n_225)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_167),
.B(n_139),
.C(n_15),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_226),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_229),
.A2(n_6),
.B1(n_227),
.B2(n_236),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_6),
.B1(n_244),
.B2(n_229),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_193),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_207),
.B1(n_221),
.B2(n_205),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_189),
.B(n_173),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_210),
.B(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_244),
.Y(n_251)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_198),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_178),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_172),
.C(n_150),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_245),
.C(n_218),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_263),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_205),
.CI(n_222),
.CON(n_254),
.SN(n_254)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_228),
.C(n_239),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_239),
.C(n_233),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_261),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_268),
.B(n_255),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_209),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_201),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_202),
.B(n_150),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_267),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_237),
.B1(n_241),
.B2(n_231),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_280),
.B(n_260),
.Y(n_290)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_266),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_256),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_246),
.C(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_258),
.C(n_264),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_242),
.B(n_230),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_286),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_260),
.A2(n_6),
.B1(n_237),
.B2(n_270),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_285),
.A2(n_251),
.B1(n_265),
.B2(n_263),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_296),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_293),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_286),
.B1(n_283),
.B2(n_254),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_261),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_264),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_275),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_300),
.A2(n_274),
.B1(n_265),
.B2(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_280),
.B(n_282),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_291),
.B(n_254),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_251),
.B1(n_282),
.B2(n_276),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_292),
.B1(n_294),
.B2(n_291),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_311),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_279),
.B(n_278),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_297),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_307),
.B1(n_302),
.B2(n_306),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_277),
.B1(n_293),
.B2(n_304),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_277),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_322),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_318),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_324),
.B1(n_319),
.B2(n_321),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_325),
.C(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_318),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_307),
.Y(n_331)
);


endmodule