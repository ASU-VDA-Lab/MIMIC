module real_jpeg_15764_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_360),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_0),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_2),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_2),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_2),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_2),
.B(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

NAND2x1_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_3),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_5),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_5),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_8),
.Y(n_361)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_10),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_10),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_10),
.B(n_194),
.Y(n_193)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_10),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_10),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_10),
.B(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g243 ( 
.A(n_12),
.Y(n_243)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_177),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_175),
.Y(n_16)
);

INVxp67_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_151),
.Y(n_18)
);

AND2x4_ASAP7_75t_SL g176 ( 
.A(n_19),
.B(n_151),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_91),
.C(n_115),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_20),
.B(n_91),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_21),
.B(n_64),
.C(n_75),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.C(n_45),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_22),
.B(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_23),
.A2(n_33),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.Y(n_23)
);

NAND2x1p5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_24),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_24),
.A2(n_66),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_24),
.B(n_94),
.C(n_99),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_24),
.A2(n_66),
.B1(n_143),
.B2(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_27),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_37),
.B(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_31),
.C(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_28),
.A2(n_37),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_28),
.A2(n_120),
.B1(n_240),
.B2(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_30),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_30),
.B(n_31),
.C(n_213),
.Y(n_290)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_31),
.A2(n_34),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_31),
.A2(n_34),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_33),
.A2(n_187),
.B(n_193),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_34),
.B(n_82),
.C(n_107),
.Y(n_169)
);

XOR2x1_ASAP7_75t_L g333 ( 
.A(n_35),
.B(n_45),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_36),
.Y(n_277)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_37),
.A2(n_121),
.B1(n_188),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_37),
.A2(n_78),
.B1(n_121),
.B2(n_135),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_37),
.B(n_78),
.C(n_226),
.Y(n_314)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_41),
.B(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_58),
.Y(n_45)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_47),
.A2(n_48),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_47),
.A2(n_48),
.B1(n_99),
.B2(n_100),
.Y(n_221)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_53),
.C(n_114),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_48),
.A2(n_100),
.B(n_198),
.C(n_252),
.Y(n_276)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_58),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_58),
.B(n_134),
.C(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_58),
.A2(n_85),
.B1(n_114),
.B2(n_134),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_58),
.A2(n_114),
.B1(n_213),
.B2(n_216),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_95),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_59),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_75),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_65),
.B(n_68),
.C(n_71),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_66),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_68),
.A2(n_74),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_68),
.A2(n_74),
.B1(n_173),
.B2(n_174),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_68),
.B(n_100),
.C(n_129),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_76),
.C(n_89),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_70),
.A2(n_71),
.B1(n_137),
.B2(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_137),
.C(n_139),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_71),
.B(n_89),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_71),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_71),
.B(n_82),
.C(n_226),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_76),
.A2(n_77),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_78),
.A2(n_85),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_82),
.A2(n_106),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_123),
.B(n_131),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_85),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_85),
.B(n_124),
.Y(n_303)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_89),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_140),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_92),
.B(n_103),
.C(n_113),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_94),
.A2(n_285),
.B(n_289),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_94),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_99),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_99),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_99),
.B(n_259),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_114),
.B(n_216),
.C(n_299),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_115),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_136),
.C(n_147),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_116),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_132),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_122),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_125),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_128),
.A2(n_129),
.B1(n_193),
.B2(n_195),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_128),
.A2(n_129),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_R g249 ( 
.A1(n_129),
.A2(n_193),
.B(n_250),
.C(n_252),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_129),
.B(n_193),
.Y(n_252)
);

XOR2x2_ASAP7_75t_L g345 ( 
.A(n_132),
.B(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_136),
.A2(n_147),
.B1(n_148),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_136),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_137),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_139),
.B(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_140),
.A2(n_143),
.B1(n_229),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_140),
.Y(n_311)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_143),
.Y(n_229)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_145),
.Y(n_288)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_166),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI321xp33_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_317),
.A3(n_348),
.B1(n_353),
.B2(n_354),
.C(n_359),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_292),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_269),
.B(n_291),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_230),
.B(n_268),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_208),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_184),
.B(n_208),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.C(n_201),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_196),
.A2(n_201),
.B1(n_202),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_198),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_198),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_205),
.A2(n_226),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_217),
.B2(n_218),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_217),
.C(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_224),
.C(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_229),
.A2(n_239),
.B(n_240),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_247),
.B(n_267),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_235),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_244),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_244),
.B1(n_245),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_256),
.B(n_266),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_253),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_263),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_265),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_260),
.B(n_261),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_271),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_274),
.C(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_278),
.C(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_284),
.C(n_290),
.Y(n_316)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_294),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_307),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_295),
.B(n_308),
.C(n_316),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_305),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_301),
.C(n_305),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_316),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_314),
.C(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_336),
.Y(n_317)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_334),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_334),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.C(n_331),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_332),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.C(n_327),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI31xp67_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_349),
.A3(n_355),
.B(n_358),
.Y(n_354)
);

NAND2x1p5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_339),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.C(n_345),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_345),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_352),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);


endmodule