module fake_jpeg_14971_n_359 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_SL g18 ( 
.A(n_16),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_SL g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_22),
.B(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_29),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_61),
.Y(n_93)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_19),
.B1(n_23),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_19),
.B1(n_56),
.B2(n_29),
.Y(n_81)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_81),
.A2(n_65),
.B1(n_71),
.B2(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

NOR5xp2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_43),
.C(n_34),
.D(n_24),
.E(n_21),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_115),
.B(n_37),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_92),
.B1(n_116),
.B2(n_28),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_94),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_98),
.B(n_100),
.Y(n_149)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_40),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_105),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_40),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_108),
.Y(n_145)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_21),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_59),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_112),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_35),
.B(n_41),
.C(n_20),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_58),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_120),
.B1(n_58),
.B2(n_61),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_26),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_60),
.A2(n_35),
.B1(n_28),
.B2(n_39),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_46),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_80),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_141),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_45),
.B(n_44),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_142),
.B1(n_151),
.B2(n_88),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_146),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_45),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_107),
.B(n_65),
.C(n_93),
.Y(n_146)
);

AO22x2_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_52),
.B1(n_58),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_148),
.A2(n_150),
.B1(n_88),
.B2(n_76),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_154),
.Y(n_198)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_163),
.B1(n_174),
.B2(n_143),
.Y(n_199)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_168),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_98),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_170),
.B(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_85),
.C(n_94),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_130),
.C(n_136),
.Y(n_194)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_97),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_95),
.B1(n_84),
.B2(n_82),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_111),
.B1(n_131),
.B2(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_104),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_172),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_120),
.B1(n_119),
.B2(n_117),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_99),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_134),
.B1(n_142),
.B2(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_193),
.B1(n_208),
.B2(n_174),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_133),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_194),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_125),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_190),
.B(n_169),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_146),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_199),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_142),
.B1(n_144),
.B2(n_143),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_149),
.C(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_160),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_39),
.B1(n_121),
.B2(n_37),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_144),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_106),
.C(n_26),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_83),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_209),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_210),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_109),
.B1(n_96),
.B2(n_135),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_121),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_217),
.B1(n_238),
.B2(n_181),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_223),
.B1(n_31),
.B2(n_33),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_163),
.B1(n_158),
.B2(n_155),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_216),
.A2(n_218),
.B1(n_224),
.B2(n_226),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_168),
.B1(n_159),
.B2(n_165),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_227),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_193),
.B1(n_188),
.B2(n_183),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_152),
.B1(n_156),
.B2(n_135),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_140),
.B1(n_177),
.B2(n_178),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_167),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_172),
.A3(n_166),
.B1(n_20),
.B2(n_28),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_39),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_236),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_36),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_192),
.A2(n_137),
.B1(n_53),
.B2(n_54),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_235),
.A2(n_240),
.B1(n_241),
.B2(n_38),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_194),
.A2(n_173),
.B1(n_103),
.B2(n_38),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_173),
.B1(n_103),
.B2(n_38),
.Y(n_241)
);

A2O1A1O1Ixp25_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_189),
.B(n_205),
.C(n_202),
.D(n_209),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_212),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_195),
.B(n_184),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_251),
.B1(n_222),
.B2(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_190),
.B(n_201),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_196),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_201),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_0),
.B(n_1),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_233),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_38),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_26),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_264),
.C(n_220),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_26),
.C(n_36),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_265),
.A2(n_214),
.B1(n_217),
.B2(n_234),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_215),
.B1(n_216),
.B2(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_286),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_220),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_277),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_212),
.B1(n_237),
.B2(n_232),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_284),
.B1(n_261),
.B2(n_257),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_259),
.C(n_256),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_248),
.B(n_218),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_226),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.C(n_282),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_242),
.Y(n_282)
);

AO21x2_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_240),
.B(n_1),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_R g286 ( 
.A(n_250),
.B(n_18),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_36),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_258),
.C(n_255),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_8),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_8),
.B(n_17),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_274),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_254),
.B(n_247),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_253),
.C(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_297),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_296),
.B(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_249),
.C(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_298),
.B(n_302),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_260),
.C(n_33),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_306),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_33),
.C(n_31),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_284),
.B1(n_275),
.B2(n_288),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_301),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_299),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_322),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_290),
.C(n_302),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_284),
.B(n_282),
.C(n_280),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_317),
.B(n_321),
.Y(n_329)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_289),
.A2(n_278),
.B1(n_287),
.B2(n_2),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_313),
.A2(n_31),
.B1(n_14),
.B2(n_11),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_33),
.B1(n_31),
.B2(n_8),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_314),
.B(n_11),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_291),
.A2(n_7),
.B(n_17),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_297),
.A2(n_7),
.B(n_17),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_326),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_294),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_330),
.C(n_332),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_309),
.C(n_303),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_10),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_292),
.C(n_296),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_313),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_319),
.B(n_316),
.Y(n_334)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_316),
.B(n_320),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_323),
.B(n_3),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_336),
.A2(n_342),
.B1(n_9),
.B2(n_1),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_310),
.B(n_14),
.C(n_11),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_337),
.A2(n_0),
.B(n_2),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_342),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_18),
.C(n_10),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_327),
.Y(n_344)
);

OR2x6_ASAP7_75t_SL g342 ( 
.A(n_332),
.B(n_9),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_344),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_346),
.C(n_347),
.Y(n_351)
);

OAI31xp67_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_338),
.A3(n_323),
.B(n_339),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_0),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_349),
.A2(n_338),
.B(n_345),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_353),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_350),
.B(n_351),
.Y(n_355)
);

AOI322xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_353),
.C2(n_352),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_3),
.B(n_4),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_3),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_5),
.B(n_6),
.Y(n_359)
);


endmodule