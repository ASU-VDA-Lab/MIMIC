module fake_jpeg_23863_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_30),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_9),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_65),
.B1(n_72),
.B2(n_28),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_56),
.B1(n_59),
.B2(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_24),
.B1(n_17),
.B2(n_29),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_59)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_33),
.B1(n_28),
.B2(n_21),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_42),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_35),
.B1(n_21),
.B2(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_44),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_85),
.B(n_90),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_83),
.B1(n_95),
.B2(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_89),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_66),
.B(n_25),
.Y(n_125)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_18),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_91),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_44),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_89),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_0),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_35),
.B1(n_23),
.B2(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_32),
.B(n_50),
.C(n_46),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_55),
.B1(n_66),
.B2(n_20),
.Y(n_132)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_32),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_20),
.B1(n_31),
.B2(n_25),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_63),
.B1(n_59),
.B2(n_65),
.Y(n_121)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_104),
.B1(n_71),
.B2(n_64),
.Y(n_128)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_105),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_0),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_25),
.C(n_15),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_118),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_77),
.B1(n_75),
.B2(n_53),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_121),
.B1(n_122),
.B2(n_134),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_123),
.Y(n_165)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_77),
.A2(n_71),
.B1(n_58),
.B2(n_64),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_132),
.B1(n_133),
.B2(n_101),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_103),
.Y(n_161)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_84),
.Y(n_146)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_104),
.B1(n_73),
.B2(n_87),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_105),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_81),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_75),
.A2(n_20),
.B1(n_49),
.B2(n_46),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_50),
.B1(n_49),
.B2(n_31),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_138),
.B(n_142),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_81),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_82),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_119),
.B(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_98),
.B1(n_74),
.B2(n_79),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_149),
.B1(n_132),
.B2(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_136),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_31),
.B(n_25),
.C(n_96),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_154),
.B(n_120),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_155),
.B1(n_164),
.B2(n_123),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_25),
.B(n_91),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_20),
.B1(n_25),
.B2(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_103),
.C(n_2),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_112),
.C(n_3),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_113),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_162),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_169),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_114),
.CI(n_125),
.CON(n_170),
.SN(n_170)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_170),
.B(n_177),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_180),
.B1(n_185),
.B2(n_137),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_176),
.B(n_196),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_151),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_179),
.A2(n_183),
.B1(n_192),
.B2(n_152),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_182),
.B(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_137),
.A2(n_117),
.B1(n_109),
.B2(n_119),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_127),
.B1(n_126),
.B2(n_118),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_115),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_115),
.B1(n_127),
.B2(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_195),
.C(n_164),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_112),
.C(n_130),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_2),
.B(n_4),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_152),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_203),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_208),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_207),
.B1(n_221),
.B2(n_198),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_166),
.B1(n_152),
.B2(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_181),
.C(n_182),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_10),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_184),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_187),
.A2(n_172),
.B1(n_180),
.B2(n_174),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_225),
.C(n_6),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_152),
.C(n_130),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_230),
.B1(n_178),
.B2(n_169),
.Y(n_235)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_184),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_248),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_203),
.B(n_206),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_201),
.B(n_220),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_241),
.B1(n_254),
.B2(n_219),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_250),
.B(n_210),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_198),
.B1(n_170),
.B2(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_199),
.B1(n_168),
.B2(n_170),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_130),
.B1(n_4),
.B2(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_11),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_6),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_214),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_222),
.C(n_214),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_201),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_275),
.C(n_16),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_255),
.B(n_8),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_208),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_202),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_269),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_231),
.CI(n_216),
.CON(n_266),
.SN(n_266)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_266),
.B(n_9),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_267),
.B(n_270),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_243),
.B1(n_234),
.B2(n_248),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_206),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_202),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_217),
.C(n_204),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_211),
.Y(n_277)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_233),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_291),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_257),
.B1(n_250),
.B2(n_245),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_285),
.A2(n_286),
.B1(n_295),
.B2(n_261),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_245),
.B1(n_238),
.B2(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_294),
.B(n_276),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_265),
.B1(n_271),
.B2(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_285),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_258),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_268),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_295),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_305),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_269),
.B(n_273),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_269),
.B(n_266),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_309),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_311),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_267),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_278),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_323),
.B(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_291),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_324),
.C(n_296),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_281),
.C(n_283),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_289),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_333),
.B(n_330),
.Y(n_338)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_289),
.B1(n_286),
.B2(n_283),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_313),
.B1(n_317),
.B2(n_263),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_331),
.B(n_12),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_284),
.B1(n_259),
.B2(n_298),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_314),
.A2(n_266),
.B(n_280),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_336),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_10),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_337),
.A2(n_338),
.B(n_339),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_325),
.A2(n_326),
.B(n_329),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_SL g343 ( 
.A(n_340),
.B(n_12),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_343),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_341),
.A2(n_334),
.B(n_335),
.Y(n_345)
);

AOI211xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_342),
.B(n_14),
.C(n_15),
.Y(n_346)
);

OAI21x1_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_344),
.B(n_13),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_13),
.C(n_14),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_13),
.Y(n_349)
);


endmodule