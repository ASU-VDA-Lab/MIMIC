module fake_jpeg_28037_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_46),
.B1(n_41),
.B2(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_82),
.B1(n_84),
.B2(n_45),
.Y(n_88)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_50),
.B1(n_54),
.B2(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_55),
.B1(n_52),
.B2(n_42),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_62),
.B1(n_57),
.B2(n_63),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_48),
.B1(n_51),
.B2(n_49),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_91),
.B(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_61),
.C(n_49),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_95),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_2),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_0),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_1),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_88),
.B1(n_86),
.B2(n_93),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_114),
.B1(n_119),
.B2(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_4),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_110),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_5),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_123),
.B(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

CKINVDCx9p33_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_6),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_131),
.B1(n_94),
.B2(n_7),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_133),
.C(n_123),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_141),
.A2(n_142),
.B1(n_137),
.B2(n_132),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_134),
.B(n_140),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_139),
.C(n_125),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_138),
.B(n_131),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_136),
.B(n_24),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_22),
.C(n_37),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_39),
.C(n_16),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_15),
.C(n_34),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_14),
.B(n_32),
.C(n_8),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_151),
.Y(n_152)
);


endmodule