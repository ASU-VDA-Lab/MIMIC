module fake_jpeg_31235_n_473 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_50),
.Y(n_149)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_68),
.Y(n_107)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_15),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_17),
.Y(n_142)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_102),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_49),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_52),
.A2(n_42),
.B1(n_23),
.B2(n_20),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_105),
.A2(n_136),
.B1(n_82),
.B2(n_95),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_143),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_58),
.A2(n_33),
.B1(n_45),
.B2(n_43),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_114),
.A2(n_120),
.B1(n_70),
.B2(n_72),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_45),
.B1(n_39),
.B2(n_43),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_83),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_20),
.B1(n_41),
.B2(n_21),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_69),
.B(n_21),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_60),
.B(n_41),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_25),
.Y(n_184)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_151),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_40),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_191),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_74),
.B1(n_66),
.B2(n_91),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_180),
.B1(n_199),
.B2(n_145),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_108),
.A2(n_33),
.B1(n_28),
.B2(n_32),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_158),
.A2(n_176),
.B(n_194),
.Y(n_221)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_169),
.Y(n_205)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_175),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_100),
.A2(n_36),
.B1(n_32),
.B2(n_92),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_178),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_36),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_181),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g181 ( 
.A(n_112),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_127),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_182),
.A2(n_190),
.B1(n_31),
.B2(n_30),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_186),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_118),
.B(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_59),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_185),
.B(n_187),
.Y(n_226)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_101),
.B(n_22),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_79),
.C(n_90),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_47),
.C(n_31),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_133),
.A2(n_56),
.B1(n_80),
.B2(n_86),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_195),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_124),
.A2(n_76),
.B1(n_65),
.B2(n_71),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_120),
.B1(n_124),
.B2(n_97),
.Y(n_202)
);

NAND2x1_ASAP7_75t_SL g194 ( 
.A(n_147),
.B(n_18),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

BUFx6f_ASAP7_75t_SL g196 ( 
.A(n_122),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_200),
.B1(n_80),
.B2(n_86),
.Y(n_217)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_198),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_114),
.A2(n_64),
.B1(n_89),
.B2(n_67),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_208),
.B1(n_218),
.B2(n_228),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_167),
.B1(n_176),
.B2(n_188),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_198),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_157),
.A2(n_97),
.B1(n_145),
.B2(n_130),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_103),
.B1(n_99),
.B2(n_117),
.Y(n_211)
);

OA21x2_ASAP7_75t_SL g275 ( 
.A1(n_212),
.A2(n_30),
.B(n_25),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_236),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_130),
.B1(n_117),
.B2(n_103),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_156),
.B(n_132),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_181),
.C(n_196),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_153),
.B(n_47),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_230),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_163),
.A2(n_106),
.B1(n_112),
.B2(n_39),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_154),
.B(n_47),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_47),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_162),
.B(n_47),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_174),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_25),
.B1(n_18),
.B2(n_3),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_183),
.B(n_160),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_243),
.A2(n_258),
.B(n_262),
.Y(n_291)
);

INVx4_ASAP7_75t_SL g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_245),
.B(n_255),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_236),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_256),
.B1(n_271),
.B2(n_202),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_206),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_209),
.A2(n_191),
.B1(n_186),
.B2(n_195),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_181),
.B(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_260),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_220),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_261),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_165),
.B(n_164),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_265),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_172),
.B(n_168),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_201),
.B(n_159),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_1),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_278),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_231),
.A2(n_177),
.B(n_175),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_201),
.B(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_274),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_31),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_270),
.B(n_272),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_208),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_233),
.B(n_30),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_22),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_232),
.B1(n_240),
.B2(n_215),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_205),
.B(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_203),
.B1(n_207),
.B2(n_222),
.Y(n_296)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_280),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_281),
.A2(n_296),
.B1(n_307),
.B2(n_314),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_282),
.A2(n_277),
.B1(n_271),
.B2(n_255),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_288),
.B(n_22),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_244),
.A2(n_215),
.B1(n_240),
.B2(n_229),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_217),
.A3(n_230),
.B1(n_223),
.B2(n_237),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_244),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_217),
.B1(n_228),
.B2(n_214),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_301),
.A2(n_303),
.B1(n_279),
.B2(n_261),
.Y(n_326)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_302),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_217),
.B1(n_214),
.B2(n_219),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_247),
.A2(n_217),
.B1(n_204),
.B2(n_207),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_266),
.B(n_242),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_311),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_247),
.A2(n_204),
.B1(n_216),
.B2(n_222),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_235),
.C(n_241),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_272),
.C(n_263),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_270),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_325),
.C(n_337),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_268),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_326),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_252),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_333),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_262),
.B(n_264),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_323),
.A2(n_331),
.B(n_340),
.Y(n_368)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_257),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_243),
.B1(n_256),
.B2(n_253),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_327),
.A2(n_346),
.B1(n_300),
.B2(n_297),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_299),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_342),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_245),
.B1(n_249),
.B2(n_260),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_339),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_257),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_330),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_311),
.A2(n_267),
.B(n_265),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_332),
.A2(n_344),
.B1(n_341),
.B2(n_302),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_273),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_290),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_345),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_250),
.Y(n_335)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_336),
.A2(n_297),
.B1(n_310),
.B2(n_284),
.Y(n_352)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_294),
.A2(n_259),
.B1(n_251),
.B2(n_235),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_294),
.A2(n_241),
.B(n_2),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_18),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_306),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_301),
.A2(n_18),
.B1(n_2),
.B2(n_4),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_345),
.B(n_298),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_350),
.B(n_364),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_352),
.B1(n_326),
.B2(n_330),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_317),
.A2(n_287),
.B1(n_310),
.B2(n_308),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_354),
.A2(n_330),
.B1(n_340),
.B2(n_287),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_321),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_355),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_339),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_357),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_305),
.C(n_284),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_347),
.C(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_319),
.B1(n_327),
.B2(n_317),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_334),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_370),
.Y(n_380)
);

BUFx4f_ASAP7_75t_SL g367 ( 
.A(n_341),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_367),
.Y(n_384)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_295),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_283),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_4),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_322),
.Y(n_372)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_343),
.A2(n_306),
.B(n_309),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_373),
.A2(n_369),
.B(n_358),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_386),
.B1(n_387),
.B2(n_389),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_351),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_378),
.B1(n_375),
.B2(n_358),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_318),
.B1(n_319),
.B2(n_325),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_378),
.A2(n_373),
.B1(n_359),
.B2(n_371),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_379),
.B(n_368),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_318),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_385),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_370),
.B(n_337),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_366),
.A2(n_331),
.B1(n_346),
.B2(n_283),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_366),
.A2(n_293),
.B1(n_286),
.B2(n_296),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_349),
.A2(n_286),
.B1(n_293),
.B2(n_312),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_363),
.A2(n_312),
.B1(n_304),
.B2(n_7),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_348),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_358),
.A2(n_312),
.B1(n_304),
.B2(n_7),
.Y(n_394)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_394),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_395),
.Y(n_410)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_356),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_399),
.B(n_379),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_406),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_377),
.A2(n_368),
.B1(n_371),
.B2(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_413),
.C(n_380),
.Y(n_417)
);

FAx1_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_371),
.CI(n_364),
.CON(n_408),
.SN(n_408)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_409),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_350),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_353),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_412),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_367),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_362),
.C(n_367),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_414),
.A2(n_396),
.B(n_388),
.Y(n_415)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_418),
.C(n_428),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_380),
.C(n_383),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_428),
.C(n_400),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_382),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_422),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_398),
.A2(n_375),
.B1(n_381),
.B2(n_374),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_429),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_SL g426 ( 
.A(n_413),
.B(n_382),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_408),
.B(n_404),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_386),
.C(n_389),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_398),
.A2(n_381),
.B1(n_387),
.B2(n_384),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_403),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_432),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_22),
.Y(n_450)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_399),
.C(n_412),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_438),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_411),
.Y(n_435)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_435),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_440),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_408),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_388),
.Y(n_441)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_405),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_8),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_439),
.A2(n_427),
.B1(n_402),
.B2(n_410),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_447),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g446 ( 
.A1(n_435),
.A2(n_422),
.B(n_420),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_429),
.B1(n_423),
.B2(n_10),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_450),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_8),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_436),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_436),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_454),
.A2(n_455),
.B(n_450),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_452),
.A2(n_433),
.B(n_440),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_460),
.Y(n_463)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_457),
.B(n_453),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_462),
.B(n_9),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_456),
.A2(n_451),
.B(n_448),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_464),
.A2(n_454),
.B(n_459),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_465),
.A2(n_466),
.B(n_467),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_463),
.A2(n_448),
.B(n_433),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_465),
.A2(n_14),
.B(n_11),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_14),
.B(n_11),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_470),
.A2(n_468),
.B(n_13),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_11),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_13),
.Y(n_473)
);


endmodule