module fake_jpeg_21057_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_25),
.B1(n_20),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_58),
.B1(n_27),
.B2(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_32),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_21),
.B(n_31),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_36),
.B(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_25),
.B1(n_20),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_40),
.B1(n_15),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_25),
.B1(n_20),
.B2(n_18),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_17),
.B1(n_28),
.B2(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_68),
.B(n_75),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_47),
.B1(n_44),
.B2(n_46),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_32),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_21),
.B(n_15),
.C(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_74),
.B1(n_76),
.B2(n_46),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_37),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_57),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_15),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_38),
.B1(n_39),
.B2(n_26),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_15),
.B1(n_26),
.B2(n_27),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_38),
.B1(n_39),
.B2(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_26),
.B1(n_30),
.B2(n_22),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_75),
.B1(n_77),
.B2(n_76),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_84),
.B(n_101),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_53),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_93),
.B1(n_103),
.B2(n_99),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_94),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_52),
.B1(n_42),
.B2(n_43),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_22),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_69),
.B(n_59),
.C(n_78),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_68),
.B(n_69),
.Y(n_107)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_12),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_39),
.B1(n_38),
.B2(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_119),
.B1(n_120),
.B2(n_89),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_113),
.B(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_68),
.B1(n_78),
.B2(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_98),
.B1(n_92),
.B2(n_52),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_72),
.CI(n_68),
.CON(n_110),
.SN(n_110)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_114),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_3),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_1),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_70),
.B1(n_81),
.B2(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_85),
.B1(n_105),
.B2(n_99),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_48),
.C(n_64),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

OAI22x1_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_30),
.B1(n_48),
.B2(n_53),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_52),
.B1(n_97),
.B2(n_90),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_53),
.B(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_126),
.A2(n_90),
.B(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_29),
.C(n_24),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_5),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_139),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_136),
.B(n_146),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_104),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_140),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_89),
.B1(n_29),
.B2(n_0),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_29),
.B1(n_7),
.B2(n_2),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_117),
.B1(n_129),
.B2(n_121),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_29),
.B1(n_1),
.B2(n_0),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_1),
.B(n_2),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_131),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_120),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_168),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_110),
.C(n_122),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_165),
.C(n_171),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_162),
.B1(n_142),
.B2(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_152),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_114),
.C(n_111),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_119),
.C(n_123),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_135),
.B1(n_145),
.B2(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_186),
.B1(n_187),
.B2(n_173),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_181),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_134),
.C(n_136),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_134),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_146),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_163),
.C(n_154),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_160),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_140),
.B1(n_149),
.B2(n_150),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_137),
.B1(n_140),
.B2(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_157),
.B(n_163),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_158),
.B(n_126),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_162),
.CI(n_126),
.CON(n_190),
.SN(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_185),
.A2(n_166),
.B(n_153),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_186),
.B(n_183),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_192),
.A2(n_181),
.B(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_153),
.B(n_159),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_160),
.B1(n_170),
.B2(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_174),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_6),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_172),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_108),
.C(n_116),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_116),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_196),
.B1(n_108),
.B2(n_9),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_208),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_188),
.B1(n_190),
.B2(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_216),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_8),
.B(n_9),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_8),
.B(n_10),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_206),
.B1(n_219),
.B2(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_203),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_222),
.A2(n_201),
.B(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_215),
.B1(n_216),
.B2(n_210),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_227),
.A2(n_12),
.B(n_13),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_229),
.C(n_13),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_231),
.Y(n_233)
);


endmodule