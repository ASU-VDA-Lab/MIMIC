module fake_jpeg_11367_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_55),
.Y(n_87)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_11),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_58),
.B1(n_18),
.B2(n_14),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_2),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_63),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_23),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_66),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_73),
.Y(n_77)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_72),
.Y(n_90)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_9),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_4),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_16),
.B1(n_31),
.B2(n_34),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_62),
.B1(n_70),
.B2(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_34),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_108),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_19),
.B1(n_30),
.B2(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_8),
.B1(n_9),
.B2(n_118),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_19),
.B1(n_17),
.B2(n_30),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_98),
.B1(n_107),
.B2(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_102),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_19),
.C(n_17),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_100),
.C(n_122),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_44),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_43),
.B(n_36),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_113),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_51),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_4),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_40),
.A2(n_31),
.B1(n_15),
.B2(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_15),
.B1(n_38),
.B2(n_37),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_37),
.B1(n_29),
.B2(n_27),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_78),
.B1(n_122),
.B2(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_27),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_25),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_18),
.B1(n_25),
.B2(n_5),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_3),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_4),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_129),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_87),
.B(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_130),
.B(n_132),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_51),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_152),
.B(n_162),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_133),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_134),
.B(n_144),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_148),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_77),
.A2(n_4),
.B(n_6),
.C(n_8),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_93),
.B1(n_147),
.B2(n_153),
.Y(n_167)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_8),
.B1(n_77),
.B2(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_164),
.B1(n_154),
.B2(n_162),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_81),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_83),
.B1(n_115),
.B2(n_116),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_91),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_150),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_92),
.Y(n_152)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_120),
.B1(n_105),
.B2(n_112),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_160),
.B1(n_135),
.B2(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_74),
.B(n_89),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_112),
.B1(n_86),
.B2(n_88),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_76),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_163),
.C(n_141),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_93),
.B(n_78),
.C(n_121),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_99),
.A2(n_76),
.B1(n_86),
.B2(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_167),
.B1(n_188),
.B2(n_194),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_147),
.B1(n_153),
.B2(n_163),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_189),
.B(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_173),
.C(n_187),
.Y(n_203)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_133),
.A3(n_126),
.B1(n_134),
.B2(n_129),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_192),
.B(n_200),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_152),
.B(n_158),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_125),
.B1(n_161),
.B2(n_160),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_128),
.A2(n_150),
.B1(n_136),
.B2(n_123),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_130),
.A2(n_156),
.B(n_151),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_146),
.B1(n_138),
.B2(n_140),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_157),
.B1(n_149),
.B2(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_129),
.A2(n_134),
.B(n_144),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_203),
.B(n_204),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_200),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_167),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_193),
.C(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_207),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_184),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_180),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_169),
.A2(n_190),
.B1(n_198),
.B2(n_188),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_183),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_194),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_175),
.C(n_174),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_169),
.B1(n_191),
.B2(n_175),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_180),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_227),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_176),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_228),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_176),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_172),
.B(n_177),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_243),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_197),
.B1(n_182),
.B2(n_170),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_239),
.B1(n_253),
.B2(n_221),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_170),
.B(n_199),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_238),
.B(n_240),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_182),
.B(n_197),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_217),
.B1(n_205),
.B2(n_218),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_177),
.B(n_221),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_216),
.B(n_203),
.Y(n_243)
);

OAI211xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_221),
.B(n_204),
.C(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_227),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_206),
.B1(n_214),
.B2(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_255),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_222),
.B1(n_228),
.B2(n_223),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_263),
.Y(n_283)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_267),
.C(n_268),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_232),
.B1(n_235),
.B2(n_231),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_266),
.B1(n_269),
.B2(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_207),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_225),
.B1(n_213),
.B2(n_211),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_238),
.B(n_240),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_226),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_230),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_213),
.C(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_236),
.Y(n_279)
);

OAI322xp33_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_242),
.A3(n_235),
.B1(n_232),
.B2(n_249),
.C1(n_248),
.C2(n_243),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_242),
.C(n_248),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_279),
.B(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_250),
.C(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.C(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_252),
.C(n_249),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_233),
.B1(n_241),
.B2(n_247),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_292),
.B1(n_274),
.B2(n_278),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.C(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_264),
.B1(n_259),
.B2(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_283),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_269),
.B(n_246),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_290),
.B(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_246),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_303),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_284),
.B1(n_276),
.B2(n_275),
.Y(n_300)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_300),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_273),
.B1(n_279),
.B2(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_297),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

NAND4xp25_ASAP7_75t_SL g311 ( 
.A(n_305),
.B(n_301),
.C(n_302),
.D(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_301),
.C(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_307),
.C(n_297),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_313),
.Y(n_318)
);


endmodule