module fake_jpeg_28842_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_SL g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_3),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_1),
.C(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_16),
.B1(n_17),
.B2(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_45),
.B1(n_53),
.B2(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_16),
.B1(n_12),
.B2(n_15),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_12),
.B(n_21),
.C(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_57),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_16),
.B1(n_12),
.B2(n_15),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_52),
.B1(n_59),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_24),
.B1(n_25),
.B2(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_30),
.A2(n_24),
.B(n_25),
.C(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_72),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_11),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_62),
.C(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_70),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_68),
.B1(n_75),
.B2(n_76),
.Y(n_87)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_44),
.B1(n_41),
.B2(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_51),
.B1(n_54),
.B2(n_50),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_64),
.B1(n_69),
.B2(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_59),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_38),
.B1(n_17),
.B2(n_13),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_76),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_78),
.B(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_87),
.C(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_90),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_90),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_103),
.B(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_98),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_94),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_108),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_107),
.Y(n_114)
);


endmodule