module real_jpeg_31347_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_92),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_5),
.B(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_8),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_9),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_72),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_51),
.B(n_71),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_39),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_15),
.B1(n_26),
.B2(n_27),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_21),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_21),
.C(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_62),
.B(n_70),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_100),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp67_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_77),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_86),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_96),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);


endmodule