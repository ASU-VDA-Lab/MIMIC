module fake_jpeg_3476_n_432 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_47),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_15),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_60),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_16),
.B(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_75),
.B(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx9p33_ASAP7_75t_R g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_77),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_79),
.Y(n_122)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_82),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_33),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_92),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_29),
.A2(n_8),
.B1(n_13),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_35),
.B1(n_44),
.B2(n_26),
.Y(n_126)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_15),
.B(n_9),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_31),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_45),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_48),
.A2(n_28),
.B1(n_27),
.B2(n_45),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_106),
.A2(n_125),
.B1(n_136),
.B2(n_139),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_59),
.A2(n_43),
.B(n_23),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_0),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_144),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_31),
.B1(n_20),
.B2(n_43),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_123),
.A2(n_21),
.B1(n_1),
.B2(n_0),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_20),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_124),
.B(n_129),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_128),
.B1(n_153),
.B2(n_84),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_49),
.A2(n_26),
.B1(n_44),
.B2(n_42),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_38),
.Y(n_129)
);

CKINVDCx12_ASAP7_75t_R g131 ( 
.A(n_80),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_45),
.B1(n_23),
.B2(n_34),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_89),
.B(n_42),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_92),
.B(n_40),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_51),
.B(n_38),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_157),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_100),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_167),
.Y(n_230)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_105),
.B1(n_134),
.B2(n_113),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_163),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_21),
.B(n_14),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_169),
.B(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_83),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_119),
.B(n_77),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_170),
.B(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_105),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_76),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_118),
.A2(n_99),
.B1(n_123),
.B2(n_103),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_98),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_73),
.B1(n_67),
.B2(n_66),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_99),
.A2(n_63),
.B1(n_62),
.B2(n_54),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_196),
.B1(n_121),
.B2(n_145),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_103),
.B(n_9),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_13),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_105),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_105),
.A2(n_152),
.B1(n_154),
.B2(n_107),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_107),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_118),
.A2(n_7),
.B(n_10),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_114),
.C(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_195),
.Y(n_221)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_98),
.A2(n_1),
.B1(n_11),
.B2(n_12),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_117),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_1),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_110),
.A2(n_1),
.B1(n_13),
.B2(n_101),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_133),
.B(n_109),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_220),
.B1(n_177),
.B2(n_160),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_203),
.B(n_181),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_114),
.B(n_149),
.C(n_117),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_183),
.B(n_157),
.C(n_192),
.D(n_193),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_212),
.B1(n_172),
.B2(n_170),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_211),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_121),
.B1(n_145),
.B2(n_138),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_196),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_133),
.B(n_149),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_161),
.B(n_169),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_171),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_150),
.B1(n_115),
.B2(n_111),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_229),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_115),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_155),
.B(n_109),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_112),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_179),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_172),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_159),
.B(n_164),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_237),
.B(n_244),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_194),
.B(n_156),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_261),
.B1(n_203),
.B2(n_215),
.Y(n_273)
);

OAI22x1_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_244),
.B1(n_258),
.B2(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_209),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_169),
.B(n_171),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_252),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_216),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_246),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_247),
.B(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_254),
.B1(n_263),
.B2(n_220),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_219),
.B(n_215),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_200),
.A2(n_181),
.B1(n_158),
.B2(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_181),
.B1(n_158),
.B2(n_156),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_181),
.B1(n_197),
.B2(n_189),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_184),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_264),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_209),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_202),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_212),
.B1(n_205),
.B2(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_174),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_267),
.B1(n_269),
.B2(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_276),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_215),
.B1(n_233),
.B2(n_213),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_201),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_215),
.B1(n_201),
.B2(n_222),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_258),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_270),
.A2(n_261),
.B(n_202),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_236),
.B1(n_254),
.B2(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_277),
.B(n_283),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_215),
.B1(n_228),
.B2(n_235),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_250),
.B1(n_239),
.B2(n_252),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_229),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_248),
.B(n_214),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_256),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_288),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_235),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_298),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_266),
.B1(n_269),
.B2(n_272),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_246),
.C(n_243),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_305),
.Y(n_321)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_289),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_243),
.B1(n_253),
.B2(n_241),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_267),
.A2(n_240),
.B1(n_264),
.B2(n_237),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_245),
.C(n_231),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_286),
.A2(n_239),
.B1(n_247),
.B2(n_208),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_288),
.B1(n_290),
.B2(n_234),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_310),
.B(n_282),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_287),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_309),
.B(n_277),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_282),
.A2(n_260),
.B(n_232),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_232),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_276),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_298),
.Y(n_318)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_329),
.B(n_334),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_280),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_322),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_288),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_325),
.A2(n_328),
.B1(n_331),
.B2(n_332),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_285),
.Y(n_326)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_327),
.A2(n_336),
.B1(n_309),
.B2(n_295),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_272),
.B1(n_265),
.B2(n_274),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_266),
.B(n_270),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_302),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_333),
.B(n_193),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_268),
.B(n_272),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_283),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_190),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_301),
.B1(n_299),
.B2(n_294),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_339),
.A2(n_318),
.B1(n_317),
.B2(n_325),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_357),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_296),
.C(n_305),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_346),
.C(n_352),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_310),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_347),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_308),
.C(n_306),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_307),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_312),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_359),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_311),
.C(n_304),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_225),
.C(n_223),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_329),
.C(n_323),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_259),
.B1(n_218),
.B2(n_223),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_259),
.B1(n_218),
.B2(n_226),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_323),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_315),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_360),
.B(n_363),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_352),
.Y(n_366)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_367),
.Y(n_385)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_371),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_334),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_338),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_374),
.Y(n_390)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_319),
.C(n_315),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_335),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_376),
.A2(n_340),
.B1(n_349),
.B2(n_356),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_351),
.B(n_345),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_377),
.A2(n_378),
.B(n_379),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_376),
.A2(n_345),
.B(n_355),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_339),
.B(n_347),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_380),
.A2(n_365),
.B1(n_369),
.B2(n_316),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_317),
.Y(n_381)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_SL g384 ( 
.A1(n_361),
.A2(n_359),
.A3(n_357),
.B1(n_353),
.B2(n_335),
.C1(n_316),
.C2(n_358),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_373),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_391),
.A2(n_397),
.B(n_396),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_378),
.A2(n_377),
.B(n_379),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_392),
.A2(n_162),
.B(n_168),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_361),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_394),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_383),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_371),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_397),
.C(n_401),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_372),
.C(n_369),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_400),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_226),
.B1(n_180),
.B2(n_224),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_206),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_402),
.B(n_224),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_385),
.Y(n_403)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_403),
.Y(n_416)
);

AOI322xp5_ASAP7_75t_L g404 ( 
.A1(n_395),
.A2(n_382),
.A3(n_380),
.B1(n_386),
.B2(n_206),
.C1(n_224),
.C2(n_149),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_408),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_R g405 ( 
.A(n_392),
.B(n_226),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_405),
.A2(n_409),
.B(n_210),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_395),
.A2(n_398),
.B(n_400),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_401),
.B1(n_162),
.B2(n_168),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_112),
.Y(n_417)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

AOI21x1_ASAP7_75t_SL g424 ( 
.A1(n_414),
.A2(n_102),
.B(n_137),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_411),
.B(n_406),
.Y(n_415)
);

AOI31xp33_ASAP7_75t_L g421 ( 
.A1(n_415),
.A2(n_420),
.A3(n_191),
.B(n_195),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_137),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_404),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_419),
.A2(n_166),
.B(n_149),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_210),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_422),
.Y(n_428)
);

OAI21x1_ASAP7_75t_SL g427 ( 
.A1(n_423),
.A2(n_424),
.B(n_138),
.Y(n_427)
);

AOI321xp33_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_416),
.A3(n_419),
.B1(n_418),
.B2(n_417),
.C(n_102),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_426),
.A2(n_13),
.B1(n_102),
.B2(n_428),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_427),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_429),
.Y(n_431)
);

XNOR2x2_ASAP7_75t_SL g432 ( 
.A(n_431),
.B(n_430),
.Y(n_432)
);


endmodule