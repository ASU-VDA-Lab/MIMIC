module fake_ariane_1844_n_787 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_787);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_787;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_664;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_785;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_34),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_29),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_28),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_148),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_112),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_22),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_23),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_60),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_54),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_88),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_13),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_8),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_133),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_84),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_113),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_59),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_53),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_66),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_116),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_62),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_48),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_41),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_30),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_47),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_50),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_51),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_92),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_160),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_73),
.B(n_153),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_0),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_0),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

AOI22x1_ASAP7_75t_SL g227 ( 
.A1(n_163),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_200),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_162),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_158),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_167),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_170),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_159),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_161),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_5),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_5),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_244),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_169),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_175),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_R g263 ( 
.A(n_214),
.B(n_172),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

CKINVDCx6p67_ASAP7_75t_R g268 ( 
.A(n_219),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_245),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_176),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_221),
.A2(n_170),
.B1(n_177),
.B2(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_220),
.B(n_178),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_240),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_249),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_219),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_218),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_218),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_195),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_R g288 ( 
.A(n_232),
.B(n_183),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_227),
.B(n_177),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_185),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_226),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_237),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_246),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_246),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_228),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_236),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_282),
.B(n_223),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_216),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_236),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_231),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_225),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_252),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_253),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_217),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_257),
.B(n_251),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_222),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_243),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_217),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_271),
.B(n_288),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_258),
.B(n_250),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_250),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_254),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_230),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_254),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_243),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_243),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_275),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_248),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_288),
.B(n_248),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_225),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_263),
.B(n_248),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_274),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_278),
.B(n_230),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_263),
.B(n_230),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_248),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_269),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_273),
.B(n_255),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_230),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_260),
.B(n_234),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_261),
.B(n_234),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_279),
.B(n_255),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_289),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_270),
.B(n_255),
.Y(n_364)
);

NOR3xp33_ASAP7_75t_L g365 ( 
.A(n_292),
.B(n_180),
.C(n_215),
.Y(n_365)
);

AO21x2_ASAP7_75t_L g366 ( 
.A1(n_288),
.A2(n_238),
.B(n_234),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_255),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_285),
.B(n_234),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_290),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_275),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_238),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_341),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_238),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_238),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_188),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_347),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_320),
.A2(n_211),
.B1(n_205),
.B2(n_204),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_320),
.B(n_189),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

NAND2x1p5_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_6),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_328),
.B(n_337),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

NOR2x1p5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_190),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_193),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_315),
.B(n_198),
.Y(n_393)
);

BUFx8_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_201),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_312),
.B(n_7),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_309),
.A2(n_203),
.B(n_76),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_360),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_360),
.B(n_7),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_8),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_363),
.B(n_9),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_332),
.B(n_9),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

AO22x1_ASAP7_75t_L g408 ( 
.A1(n_356),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_307),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

NOR2x1_ASAP7_75t_R g414 ( 
.A(n_310),
.B(n_10),
.Y(n_414)
);

AND2x6_ASAP7_75t_SL g415 ( 
.A(n_316),
.B(n_11),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_317),
.B(n_12),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_311),
.Y(n_418)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_313),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_359),
.B(n_13),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_354),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_362),
.B(n_14),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_342),
.B(n_14),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_309),
.B(n_16),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_17),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_348),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

A2O1A1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_365),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_358),
.B(n_21),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_338),
.B(n_24),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_390),
.A2(n_352),
.B1(n_370),
.B2(n_344),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_322),
.B1(n_353),
.B2(n_334),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

NOR2x1_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_353),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_389),
.B(n_338),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_431),
.A2(n_346),
.B(n_338),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_SL g449 ( 
.A(n_379),
.B(n_349),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_383),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_SL g452 ( 
.A1(n_397),
.A2(n_349),
.B(n_338),
.C(n_27),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_338),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_431),
.A2(n_349),
.B(n_26),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_396),
.A2(n_349),
.B1(n_31),
.B2(n_32),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_373),
.B(n_25),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_416),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

O2A1O1Ixp33_ASAP7_75t_SL g461 ( 
.A1(n_437),
.A2(n_349),
.B(n_35),
.C(n_36),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_429),
.A2(n_33),
.B(n_37),
.C(n_38),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_39),
.C(n_42),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_374),
.A2(n_43),
.B(n_44),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_388),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_378),
.A2(n_55),
.B(n_56),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_393),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_400),
.B(n_63),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_R g473 ( 
.A(n_420),
.B(n_64),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_407),
.B(n_65),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_432),
.A2(n_67),
.B(n_68),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_380),
.B(n_156),
.Y(n_478)
);

AO21x1_ASAP7_75t_L g479 ( 
.A1(n_377),
.A2(n_69),
.B(n_70),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_430),
.A2(n_71),
.B(n_72),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

OAI22x1_ASAP7_75t_L g483 ( 
.A1(n_395),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_413),
.B(n_80),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_405),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_384),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_430),
.A2(n_93),
.B(n_94),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_95),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_372),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_406),
.A2(n_417),
.B(n_385),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_424),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_426),
.B(n_96),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_384),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_419),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_428),
.B(n_102),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_424),
.B(n_103),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_418),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_447),
.A2(n_440),
.B(n_402),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_448),
.A2(n_440),
.B(n_377),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_455),
.A2(n_438),
.B(n_382),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_445),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_481),
.A2(n_404),
.B(n_382),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_487),
.A2(n_404),
.B(n_434),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_477),
.A2(n_436),
.B(n_409),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_474),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_485),
.A2(n_403),
.B1(n_375),
.B2(n_391),
.Y(n_510)
);

BUFx2_ASAP7_75t_SL g511 ( 
.A(n_464),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_450),
.Y(n_512)
);

OA21x2_ASAP7_75t_L g513 ( 
.A1(n_453),
.A2(n_392),
.B(n_375),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_433),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_479),
.A2(n_408),
.B(n_425),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_409),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_474),
.Y(n_517)
);

INVx8_ASAP7_75t_L g518 ( 
.A(n_458),
.Y(n_518)
);

NAND2x1p5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_425),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_494),
.A2(n_414),
.B(n_387),
.Y(n_521)
);

AOI21x1_ASAP7_75t_L g522 ( 
.A1(n_472),
.A2(n_415),
.B(n_106),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_496),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_466),
.A2(n_104),
.B(n_111),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_469),
.A2(n_114),
.B(n_115),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_458),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_473),
.Y(n_528)
);

OA21x2_ASAP7_75t_L g529 ( 
.A1(n_462),
.A2(n_488),
.B(n_486),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_459),
.B(n_415),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_499),
.A2(n_117),
.B(n_118),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

BUFx8_ASAP7_75t_SL g533 ( 
.A(n_468),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_452),
.A2(n_497),
.B(n_461),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_476),
.B(n_119),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_121),
.Y(n_537)
);

AO21x2_ASAP7_75t_L g538 ( 
.A1(n_475),
.A2(n_123),
.B(n_125),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_454),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_446),
.B(n_126),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_492),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_492),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_492),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_483),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_498),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_498),
.Y(n_548)
);

AO21x1_ASAP7_75t_SL g549 ( 
.A1(n_510),
.A2(n_484),
.B(n_491),
.Y(n_549)
);

CKINVDCx6p67_ASAP7_75t_R g550 ( 
.A(n_504),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_507),
.Y(n_551)
);

AOI21x1_ASAP7_75t_L g552 ( 
.A1(n_529),
.A2(n_449),
.B(n_456),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_546),
.A2(n_478),
.B1(n_465),
.B2(n_443),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_520),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_539),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_509),
.Y(n_556)
);

CKINVDCx11_ASAP7_75t_R g557 ( 
.A(n_504),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_500),
.B(n_471),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_539),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_544),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_510),
.A2(n_444),
.B1(n_495),
.B2(n_467),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_518),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_546),
.A2(n_457),
.B1(n_470),
.B2(n_498),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_523),
.Y(n_565)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_509),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g567 ( 
.A1(n_529),
.A2(n_128),
.B(n_129),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_534),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_540),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_512),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_544),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_514),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_529),
.A2(n_130),
.B(n_131),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_530),
.B(n_149),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_506),
.A2(n_132),
.B(n_134),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_532),
.B(n_135),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_506),
.A2(n_136),
.B(n_138),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_513),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_502),
.A2(n_139),
.B(n_140),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_542),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_518),
.Y(n_584)
);

INVx6_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_536),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_536),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_536),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_501),
.A2(n_146),
.B1(n_147),
.B2(n_537),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_551),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_R g593 ( 
.A(n_574),
.B(n_528),
.Y(n_593)
);

AO31x2_ASAP7_75t_L g594 ( 
.A1(n_577),
.A2(n_541),
.A3(n_502),
.B(n_515),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_570),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_566),
.B(n_528),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_590),
.B(n_548),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_579),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_563),
.B(n_548),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_569),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_532),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_557),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_572),
.B(n_517),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_561),
.A2(n_521),
.B1(n_515),
.B2(n_531),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_565),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_568),
.B(n_527),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_R g607 ( 
.A(n_566),
.B(n_524),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_511),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_556),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_553),
.B(n_527),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_557),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_550),
.B(n_518),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_522),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_554),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_515),
.C(n_531),
.Y(n_616)
);

BUFx12f_ASAP7_75t_L g617 ( 
.A(n_585),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_585),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_571),
.Y(n_619)
);

CKINVDCx12_ASAP7_75t_R g620 ( 
.A(n_554),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_585),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_555),
.Y(n_622)
);

AOI221xp5_ASAP7_75t_L g623 ( 
.A1(n_589),
.A2(n_521),
.B1(n_535),
.B2(n_538),
.C(n_547),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_588),
.B(n_519),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_583),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_558),
.B(n_576),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_559),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_SL g629 ( 
.A(n_591),
.B(n_516),
.C(n_519),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_549),
.A2(n_531),
.B1(n_538),
.B2(n_535),
.Y(n_630)
);

NOR2x1_ASAP7_75t_L g631 ( 
.A(n_589),
.B(n_547),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_560),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_588),
.B(n_547),
.Y(n_633)
);

AO31x2_ASAP7_75t_L g634 ( 
.A1(n_577),
.A2(n_503),
.A3(n_525),
.B(n_526),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_583),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_576),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_562),
.B(n_542),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_626),
.A2(n_578),
.B1(n_562),
.B2(n_581),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_592),
.B(n_605),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_581),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_637),
.B(n_578),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_598),
.B(n_586),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_617),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_600),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_622),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_L g646 ( 
.A(n_616),
.B(n_584),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_613),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_586),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_627),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_628),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_636),
.B(n_576),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_632),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_606),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_625),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_609),
.B(n_533),
.Y(n_656)
);

INVx5_ASAP7_75t_SL g657 ( 
.A(n_608),
.Y(n_657)
);

OAI211xp5_ASAP7_75t_L g658 ( 
.A1(n_623),
.A2(n_552),
.B(n_567),
.C(n_573),
.Y(n_658)
);

OAI221xp5_ASAP7_75t_L g659 ( 
.A1(n_623),
.A2(n_516),
.B1(n_542),
.B2(n_533),
.C(n_525),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_594),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_606),
.B(n_575),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_635),
.B(n_575),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_594),
.B(n_580),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_580),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_582),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

AO21x2_ASAP7_75t_L g667 ( 
.A1(n_616),
.A2(n_582),
.B(n_526),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_634),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g669 ( 
.A1(n_610),
.A2(n_505),
.B(n_503),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_610),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_634),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_597),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_620),
.Y(n_674)
);

NAND4xp25_ASAP7_75t_L g675 ( 
.A(n_654),
.B(n_614),
.C(n_603),
.D(n_593),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_647),
.B(n_595),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_653),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_656),
.A2(n_631),
.B(n_630),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_639),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_670),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_672),
.B(n_599),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_655),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_642),
.B(n_607),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_645),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_642),
.B(n_608),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_661),
.B(n_608),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_640),
.B(n_611),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_644),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_640),
.B(n_641),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_661),
.B(n_648),
.Y(n_691)
);

NAND2x1_ASAP7_75t_L g692 ( 
.A(n_654),
.B(n_633),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_643),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_SL g694 ( 
.A(n_651),
.B(n_596),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_648),
.B(n_633),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_649),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_641),
.B(n_633),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_673),
.B(n_638),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_649),
.B(n_599),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_650),
.B(n_601),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_646),
.B(n_624),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_691),
.B(n_665),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_691),
.B(n_665),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_680),
.B(n_652),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_687),
.B(n_662),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_696),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_679),
.B(n_663),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_694),
.B(n_657),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_696),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_690),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_677),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_686),
.B(n_663),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_684),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_684),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_682),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_687),
.B(n_664),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_698),
.B(n_652),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_689),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_683),
.B(n_657),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_685),
.B(n_664),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_655),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_713),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_704),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_702),
.B(n_683),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_711),
.B(n_676),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_710),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_709),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_718),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_702),
.B(n_688),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_713),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_706),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_726),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_724),
.B(n_703),
.Y(n_733)
);

AOI21xp33_ASAP7_75t_SL g734 ( 
.A1(n_729),
.A2(n_602),
.B(n_708),
.Y(n_734)
);

OAI21xp33_ASAP7_75t_L g735 ( 
.A1(n_723),
.A2(n_725),
.B(n_728),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_727),
.A2(n_678),
.B1(n_675),
.B2(n_694),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_732),
.B(n_693),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_735),
.B(n_728),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_736),
.B(n_708),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_733),
.B(n_725),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_734),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_735),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_739),
.B(n_693),
.Y(n_743)
);

OAI322xp33_ASAP7_75t_L g744 ( 
.A1(n_742),
.A2(n_717),
.A3(n_699),
.B1(n_700),
.B2(n_681),
.C1(n_659),
.C2(n_692),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_712),
.Y(n_745)
);

AO22x1_ASAP7_75t_SL g746 ( 
.A1(n_743),
.A2(n_741),
.B1(n_738),
.B2(n_737),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_719),
.B(n_731),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_R g748 ( 
.A(n_746),
.B(n_612),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_747),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_747),
.B(n_745),
.C(n_643),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_749),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_750),
.A2(n_701),
.B1(n_674),
.B2(n_703),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_749),
.Y(n_754)
);

NOR4xp25_ASAP7_75t_L g755 ( 
.A(n_749),
.B(n_658),
.C(n_715),
.D(n_629),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_749),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_753),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_R g758 ( 
.A(n_751),
.B(n_715),
.Y(n_758)
);

OAI211xp5_ASAP7_75t_SL g759 ( 
.A1(n_754),
.A2(n_715),
.B(n_674),
.C(n_682),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_756),
.A2(n_716),
.B(n_701),
.C(n_731),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_752),
.A2(n_701),
.B1(n_716),
.B2(n_720),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_SL g762 ( 
.A(n_755),
.B(n_657),
.C(n_668),
.Y(n_762)
);

NOR4xp75_ASAP7_75t_L g763 ( 
.A(n_753),
.B(n_712),
.C(n_707),
.D(n_721),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_757),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_758),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_705),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_761),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_763),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_760),
.B(n_705),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_768),
.A2(n_759),
.B1(n_705),
.B2(n_657),
.Y(n_770)
);

AOI22x1_ASAP7_75t_L g771 ( 
.A1(n_765),
.A2(n_542),
.B1(n_601),
.B2(n_682),
.Y(n_771)
);

AO22x2_ASAP7_75t_L g772 ( 
.A1(n_764),
.A2(n_730),
.B1(n_722),
.B2(n_621),
.Y(n_772)
);

AND4x1_ASAP7_75t_L g773 ( 
.A(n_764),
.B(n_707),
.C(n_721),
.D(n_720),
.Y(n_773)
);

AOI22x1_ASAP7_75t_L g774 ( 
.A1(n_767),
.A2(n_662),
.B1(n_697),
.B2(n_706),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_766),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_769),
.B(n_618),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_L g777 ( 
.A1(n_775),
.A2(n_655),
.B1(n_714),
.B2(n_668),
.Y(n_777)
);

AOI31xp33_ASAP7_75t_L g778 ( 
.A1(n_776),
.A2(n_697),
.A3(n_695),
.B(n_651),
.Y(n_778)
);

AO22x2_ASAP7_75t_L g779 ( 
.A1(n_770),
.A2(n_772),
.B1(n_771),
.B2(n_773),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_SL g780 ( 
.A1(n_774),
.A2(n_671),
.B(n_714),
.C(n_650),
.Y(n_780)
);

OR3x2_ASAP7_75t_L g781 ( 
.A(n_779),
.B(n_667),
.C(n_666),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_SL g783 ( 
.A1(n_782),
.A2(n_780),
.B1(n_777),
.B2(n_624),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_783),
.A2(n_781),
.B1(n_624),
.B2(n_660),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_784),
.A2(n_667),
.B1(n_660),
.B2(n_671),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_667),
.B(n_505),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_786),
.A2(n_651),
.B1(n_669),
.B2(n_695),
.Y(n_787)
);


endmodule