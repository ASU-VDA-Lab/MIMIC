module real_jpeg_29635_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_54),
.B(n_55),
.C(n_59),
.D(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_1),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_1),
.A2(n_79),
.B(n_83),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_1),
.A2(n_24),
.B(n_117),
.C(n_118),
.D(n_122),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_1),
.B(n_24),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_2),
.B(n_23),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_101),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_64),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_64),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_4),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_4),
.A2(n_53),
.B1(n_55),
.B2(n_150),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_150),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_150),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_53),
.B1(n_55),
.B2(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_75),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_75),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_75),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_7),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_53),
.B1(n_55),
.B2(n_167),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_167),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_167),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_8),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_8),
.A2(n_53),
.B1(n_55),
.B2(n_132),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_132),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_10),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_53),
.B1(n_55),
.B2(n_82),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_82),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_82),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_11),
.A2(n_34),
.B1(n_53),
.B2(n_55),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_291)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_12),
.A2(n_55),
.B(n_60),
.C(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_12),
.B(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_30),
.B1(n_49),
.B2(n_50),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_13),
.A2(n_30),
.B1(n_53),
.B2(n_55),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_311)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_53),
.B1(n_55),
.B2(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_29),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_21),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_21),
.A2(n_25),
.B1(n_200),
.B2(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_21),
.A2(n_25),
.B1(n_33),
.B2(n_327),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_22),
.A2(n_27),
.B(n_101),
.C(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_23),
.A2(n_24),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_23),
.A2(n_55),
.A3(n_117),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_25),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_25),
.B(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_25),
.Y(n_241)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_32),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_32),
.B(n_333),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_332),
.B(n_334),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_320),
.B(n_331),
.Y(n_38)
);

OAI321xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_284),
.A3(n_313),
.B1(n_318),
.B2(n_319),
.C(n_336),
.Y(n_39)
);

AOI321xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_234),
.A3(n_273),
.B1(n_278),
.B2(n_283),
.C(n_337),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_187),
.C(n_230),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_158),
.B(n_186),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_137),
.B(n_157),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_112),
.B(n_136),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_88),
.B(n_111),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_66),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_47),
.B(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_58),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_58),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.A3(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_49),
.B(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_57),
.Y(n_56)
);

NAND2x1_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_53),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_59),
.A2(n_61),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_59),
.A2(n_61),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_59),
.A2(n_61),
.B1(n_250),
.B2(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_74),
.B(n_76),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_65),
.A2(n_76),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_65),
.A2(n_154),
.B1(n_185),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_65),
.A2(n_154),
.B1(n_208),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_65),
.A2(n_154),
.B(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_78),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_73),
.C(n_78),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_70),
.A2(n_118),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_70),
.A2(n_118),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_70),
.A2(n_118),
.B1(n_262),
.B2(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_70),
.A2(n_118),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_74),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_79),
.A2(n_96),
.B1(n_131),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_79),
.A2(n_96),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_79),
.A2(n_206),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_79),
.A2(n_223),
.B(n_224),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_86),
.A2(n_93),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx5_ASAP7_75t_SL g223 ( 
.A(n_86),
.Y(n_223)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_101),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_98),
.B(n_110),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_96),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_104),
.B(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_105),
.B(n_109),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_114),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_128),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_125),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_125),
.C(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_124),
.A2(n_143),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_124),
.A2(n_195),
.B1(n_220),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_124),
.A2(n_195),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_133),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_139),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_151),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_152),
.C(n_153),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_146),
.C(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_199),
.B(n_201),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_147),
.A2(n_201),
.B(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_147),
.A2(n_241),
.B1(n_269),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_147),
.A2(n_241),
.B1(n_296),
.B2(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_160),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_172),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_163),
.C(n_172),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_166),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_171),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_180),
.C(n_183),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_176),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_182),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_188),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_210),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_189),
.B(n_210),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_203),
.C(n_209),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_193),
.C(n_202),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_198),
.B2(n_202),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B(n_197),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_209),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_221),
.C(n_229),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_216),
.C(n_218),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_225),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_254),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_254),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_246),
.C(n_253),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_246),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_245),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_243),
.C(n_245),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_252),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_252),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_267),
.B(n_270),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_264),
.B1(n_265),
.B2(n_271),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_260),
.B(n_263),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_263),
.A2(n_286),
.B1(n_287),
.B2(n_298),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_271),
.C(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_279),
.B(n_282),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_301),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_301),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.C(n_299),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_297),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_290),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_294),
.C(n_295),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_294),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_305),
.C(n_309),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_304),
.C(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_300),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_312),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_306),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_311),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_322),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_326),
.B1(n_328),
.B2(n_329),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_324),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_326),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_329),
.C(n_330),
.Y(n_333)
);


endmodule