module fake_jpeg_5820_n_298 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_121;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_46),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx9p33_ASAP7_75t_R g88 ( 
.A(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_36),
.B(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_11),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_16),
.B(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_23),
.B1(n_30),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_73),
.B1(n_76),
.B2(n_91),
.Y(n_117)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_61),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_18),
.B1(n_29),
.B2(n_13),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_63),
.B1(n_94),
.B2(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_30),
.B1(n_13),
.B2(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_79),
.B1(n_81),
.B2(n_86),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_78),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_25),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_14),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_14),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_89),
.Y(n_102)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_93),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_37),
.A2(n_27),
.B1(n_20),
.B2(n_15),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_43),
.A2(n_27),
.B1(n_20),
.B2(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_7),
.B(n_11),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_26),
.C(n_28),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_26),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_67),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_108),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_104),
.A2(n_112),
.B1(n_115),
.B2(n_92),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_21),
.B1(n_28),
.B2(n_10),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_56),
.A2(n_28),
.B1(n_16),
.B2(n_2),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_51),
.B1(n_91),
.B2(n_81),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_0),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_10),
.B(n_8),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_132),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_48),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_124),
.C(n_125),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_59),
.B1(n_92),
.B2(n_74),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_157),
.B1(n_160),
.B2(n_116),
.Y(n_163)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_55),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_100),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_89),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_102),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_54),
.Y(n_140)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_65),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_102),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_64),
.B(n_87),
.C(n_79),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_110),
.B(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_52),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_148),
.Y(n_176)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_109),
.B(n_72),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_152),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_105),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_153),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_86),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_118),
.B(n_59),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_156),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_66),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_104),
.A2(n_88),
.B1(n_16),
.B2(n_53),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_53),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_163),
.A2(n_177),
.B1(n_186),
.B2(n_144),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_126),
.B1(n_122),
.B2(n_133),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_180),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_179),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_173),
.B(n_75),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_137),
.B1(n_147),
.B2(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_193),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_100),
.B(n_114),
.Y(n_179)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_108),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_145),
.C(n_7),
.D(n_3),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_114),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_138),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_122),
.B1(n_106),
.B2(n_119),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_187),
.B(n_191),
.Y(n_205)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_66),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_204),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_211),
.B1(n_218),
.B2(n_194),
.Y(n_219)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_134),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_148),
.B1(n_153),
.B2(n_161),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_207),
.B1(n_209),
.B2(n_191),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_139),
.B1(n_152),
.B2(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_214),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_135),
.B1(n_150),
.B2(n_161),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_213),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_194),
.B1(n_178),
.B2(n_186),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_176),
.B(n_182),
.Y(n_237)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_126),
.A3(n_106),
.B1(n_129),
.B2(n_4),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_175),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_221),
.B1(n_201),
.B2(n_205),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_184),
.B1(n_187),
.B2(n_172),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_169),
.B(n_184),
.C(n_179),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_237),
.B(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_171),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.C(n_238),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_206),
.B(n_203),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_184),
.C(n_172),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_163),
.C(n_164),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_254),
.B1(n_228),
.B2(n_164),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_247),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_224),
.B1(n_220),
.B2(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_246),
.B(n_231),
.Y(n_264)
);

OAI321xp33_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_222),
.A3(n_224),
.B1(n_223),
.B2(n_210),
.C(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_196),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_217),
.C(n_212),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_243),
.C(n_254),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_200),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_228),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_230),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_235),
.B1(n_230),
.B2(n_218),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_237),
.B1(n_205),
.B2(n_238),
.Y(n_254)
);

AOI321xp33_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_222),
.A3(n_227),
.B1(n_232),
.B2(n_236),
.C(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_243),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_264),
.B(n_242),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_180),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_249),
.C(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_167),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_266),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_239),
.A2(n_231),
.B1(n_170),
.B2(n_197),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_274),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_252),
.B1(n_244),
.B2(n_248),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_257),
.A3(n_256),
.B1(n_264),
.B2(n_266),
.C1(n_255),
.C2(n_174),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_255),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_272),
.C(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_246),
.Y(n_272)
);

NAND4xp25_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_198),
.C(n_189),
.D(n_128),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_242),
.C(n_170),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_279),
.B(n_273),
.Y(n_287)
);

OAI211xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_280),
.B(n_121),
.C(n_165),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_174),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_121),
.C(n_129),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_121),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_276),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_273),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_269),
.B1(n_270),
.B2(n_267),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_289),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_165),
.B(n_180),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_296)
);

AOI321xp33_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_121),
.A3(n_128),
.B1(n_75),
.B2(n_4),
.C(n_5),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_293),
.B(n_291),
.Y(n_298)
);


endmodule