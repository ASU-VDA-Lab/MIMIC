module fake_ariane_1369_n_1661 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1661);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1661;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_57),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_26),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_74),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_22),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_52),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_87),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_10),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_47),
.Y(n_160)
);

INVxp33_ASAP7_75t_R g161 ( 
.A(n_99),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_25),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_79),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_34),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_59),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_89),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_7),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_111),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_8),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_119),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_2),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

BUFx8_ASAP7_75t_SL g187 ( 
.A(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_44),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_30),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_42),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_30),
.Y(n_193)
);

BUFx2_ASAP7_75t_SL g194 ( 
.A(n_124),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_127),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_68),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_46),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_49),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_71),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_86),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_54),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_23),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_24),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_113),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_26),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_48),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_56),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_27),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_115),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_6),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_131),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_37),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_73),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_38),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_11),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_19),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_19),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_93),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_36),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_34),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_32),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_3),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_82),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_67),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_17),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_64),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_22),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_41),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_83),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_28),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_122),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_97),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_69),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_78),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_0),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_109),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_28),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_62),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_39),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_51),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_43),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_6),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_13),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_27),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_76),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_123),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_16),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_14),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_108),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_94),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_8),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_91),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_37),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_66),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_25),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_21),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_60),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_120),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_65),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_5),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_39),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_110),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_20),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_4),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_183),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_187),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_187),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_169),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_178),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_178),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_149),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_153),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_147),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_196),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_159),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_196),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_144),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_159),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_153),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_144),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_205),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_152),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_162),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_179),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_162),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_189),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_173),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_205),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_208),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_197),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_208),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_230),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_211),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_181),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_209),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_215),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_209),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_175),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_218),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_188),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_213),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_185),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_190),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_221),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_204),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_230),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_251),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_212),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_163),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_225),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_189),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_237),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_226),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_173),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_227),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_228),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_234),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_231),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_232),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_149),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_242),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_239),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_244),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_163),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_261),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_262),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_275),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_282),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_155),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_308),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g366 ( 
.A1(n_308),
.A2(n_150),
.B(n_141),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_290),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_287),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_329),
.B(n_155),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_288),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_315),
.B(n_342),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

OAI21x1_ASAP7_75t_L g376 ( 
.A1(n_316),
.A2(n_166),
.B(n_157),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_297),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_298),
.B(n_250),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_186),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_229),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_289),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_329),
.B(n_189),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_146),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_319),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_293),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_302),
.B(n_250),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_349),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_294),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_291),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_293),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_325),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_298),
.B(n_216),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_307),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_361),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_295),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_295),
.Y(n_404)
);

AND3x2_ASAP7_75t_L g405 ( 
.A(n_292),
.B(n_161),
.C(n_156),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_296),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_296),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_355),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_299),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_299),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_326),
.B(n_214),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_301),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_301),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_304),
.B(n_274),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_320),
.B(n_274),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_335),
.B(n_220),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_300),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_216),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_328),
.B(n_284),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_331),
.B(n_284),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_219),
.Y(n_424)
);

BUFx8_ASAP7_75t_L g425 ( 
.A(n_314),
.Y(n_425)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_331),
.B(n_194),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_303),
.B(n_219),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_313),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_336),
.A2(n_180),
.B(n_170),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_336),
.B(n_182),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_428),
.B(n_335),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_377),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

OR2x6_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_343),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

CKINVDCx6p67_ASAP7_75t_R g440 ( 
.A(n_392),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_339),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_425),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_428),
.B(n_322),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_310),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_343),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_400),
.B(n_312),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

CKINVDCx6p67_ASAP7_75t_R g465 ( 
.A(n_391),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

BUFx4f_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_344),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_400),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_318),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_398),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_403),
.B(n_408),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_412),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_426),
.B(n_344),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_417),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_429),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_362),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_362),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_395),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_364),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_364),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_401),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_364),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_371),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_431),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_363),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_371),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_371),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_365),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_371),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_400),
.B(n_321),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_372),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_400),
.B(n_324),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_400),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_408),
.B(n_327),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_365),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_R g513 ( 
.A(n_367),
.B(n_306),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_427),
.B(n_346),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_368),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_368),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_371),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_369),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_366),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_372),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_369),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_370),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_370),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_311),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_408),
.B(n_337),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_371),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_431),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_424),
.A2(n_356),
.B1(n_172),
.B2(n_191),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_371),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_380),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_373),
.Y(n_532)
);

CKINVDCx6p67_ASAP7_75t_R g533 ( 
.A(n_385),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_373),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_373),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_373),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_393),
.B(n_332),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_430),
.B(n_346),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_373),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_373),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_380),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_373),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_383),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_409),
.B(n_338),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_421),
.B(n_341),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_404),
.Y(n_548)
);

AND3x2_ASAP7_75t_L g549 ( 
.A(n_390),
.B(n_347),
.C(n_340),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_383),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_430),
.B(n_348),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_409),
.B(n_345),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_387),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_409),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_387),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_394),
.Y(n_557)
);

AND3x2_ASAP7_75t_L g558 ( 
.A(n_390),
.B(n_350),
.C(n_348),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_404),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_385),
.B(n_352),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_394),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_390),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_379),
.B(n_330),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_406),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_397),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_374),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_406),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_406),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_399),
.B(n_350),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_397),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_366),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_422),
.B(n_351),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_407),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_399),
.B(n_351),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_424),
.B(n_154),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_407),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_407),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_366),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_411),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_422),
.B(n_354),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_366),
.Y(n_581)
);

CKINVDCx11_ASAP7_75t_R g582 ( 
.A(n_435),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_449),
.B(n_412),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_466),
.B(n_424),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_546),
.B(n_416),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_416),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_564),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_529),
.A2(n_255),
.B1(n_193),
.B2(n_233),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_560),
.B(n_419),
.C(n_418),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_564),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_493),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_562),
.A2(n_171),
.B1(n_172),
.B2(n_191),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_526),
.B(n_416),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_562),
.A2(n_376),
.B(n_424),
.C(n_432),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_433),
.B(n_447),
.C(n_547),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_564),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_566),
.B(n_418),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_466),
.B(n_418),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_548),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_548),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_466),
.B(n_379),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_566),
.B(n_425),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_425),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_437),
.A2(n_488),
.B1(n_456),
.B2(n_468),
.Y(n_606)
);

OAI221xp5_ASAP7_75t_L g607 ( 
.A1(n_569),
.A2(n_223),
.B1(n_259),
.B2(n_386),
.C(n_381),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_425),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_425),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_466),
.B(n_432),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_511),
.B(n_381),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_488),
.B(n_374),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_452),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_563),
.B(n_452),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_553),
.B(n_386),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_444),
.B(n_171),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_437),
.A2(n_198),
.B1(n_378),
.B2(n_193),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_378),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_422),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_543),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_437),
.A2(n_198),
.B1(n_378),
.B2(n_185),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_467),
.B(n_376),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_494),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_468),
.B(n_378),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_514),
.B(n_423),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_467),
.B(n_376),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_514),
.B(n_423),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_474),
.B(n_423),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_559),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_538),
.B(n_388),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_538),
.B(n_552),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_502),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_552),
.B(n_388),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_475),
.B(n_402),
.Y(n_637)
);

INVx8_ASAP7_75t_L g638 ( 
.A(n_443),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_440),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_444),
.B(n_154),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_437),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_571),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_475),
.B(n_402),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_475),
.B(n_410),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_572),
.B(n_410),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_543),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_533),
.B(n_413),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_467),
.A2(n_431),
.B1(n_233),
.B2(n_255),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_572),
.B(n_413),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_580),
.B(n_437),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_505),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_537),
.B(n_270),
.C(n_240),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_505),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_533),
.B(n_414),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_SL g657 ( 
.A(n_580),
.B(n_270),
.C(n_253),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_512),
.B(n_515),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_414),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_465),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_558),
.B(n_508),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_515),
.B(n_411),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_442),
.B(n_252),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_519),
.B(n_160),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_471),
.B(n_405),
.Y(n_667)
);

AO21x2_ASAP7_75t_L g668 ( 
.A1(n_571),
.A2(n_199),
.B(n_201),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_490),
.A2(n_411),
.B1(n_357),
.B2(n_354),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_549),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_440),
.B(n_444),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_578),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_518),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_518),
.B(n_148),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_519),
.A2(n_220),
.B1(n_257),
.B2(n_246),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_521),
.B(n_158),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_575),
.B(n_260),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_459),
.B(n_412),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_462),
.B(n_265),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_519),
.A2(n_581),
.B1(n_578),
.B2(n_523),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_444),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_471),
.B(n_160),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_521),
.B(n_202),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_523),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_524),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_513),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_498),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_524),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_568),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_476),
.A2(n_271),
.B1(n_278),
.B2(n_164),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_510),
.B(n_520),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_531),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_531),
.Y(n_694)
);

AND2x4_ASAP7_75t_SL g695 ( 
.A(n_510),
.B(n_272),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_541),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_568),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_507),
.B(n_266),
.Y(n_699)
);

BUFx6f_ASAP7_75t_SL g700 ( 
.A(n_544),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_544),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_459),
.B(n_460),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_550),
.A2(n_360),
.B(n_359),
.C(n_358),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_509),
.B(n_279),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_581),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_550),
.B(n_249),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_554),
.B(n_254),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_554),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_556),
.B(n_269),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_573),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_556),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_557),
.B(n_164),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_557),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_561),
.A2(n_271),
.B1(n_278),
.B2(n_222),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_576),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_576),
.Y(n_717)
);

AND2x4_ASAP7_75t_SL g718 ( 
.A(n_561),
.B(n_272),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_565),
.B(n_222),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_565),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_357),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_577),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_460),
.B(n_358),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_470),
.B(n_203),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_470),
.B(n_359),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_472),
.B(n_280),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_543),
.Y(n_727)
);

BUFx6f_ASAP7_75t_SL g728 ( 
.A(n_487),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_472),
.B(n_285),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_477),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_477),
.B(n_286),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_478),
.B(n_142),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_577),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_464),
.A2(n_220),
.B1(n_246),
.B2(n_257),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_579),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_478),
.B(n_483),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_483),
.B(n_143),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_555),
.B(n_145),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_464),
.B(n_206),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_487),
.B(n_151),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_489),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_SL g742 ( 
.A(n_489),
.B(n_165),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_458),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_492),
.B(n_167),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_492),
.B(n_168),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_612),
.B(n_585),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_650),
.A2(n_501),
.B1(n_522),
.B2(n_528),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_638),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_612),
.B(n_464),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_603),
.B(n_586),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_622),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_582),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_709),
.A2(n_439),
.B1(n_464),
.B2(n_501),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_600),
.B(n_458),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_603),
.B(n_405),
.Y(n_755)
);

NOR2x1p5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_439),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_601),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_592),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_642),
.B(n_661),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_599),
.B(n_600),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_706),
.B(n_439),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_687),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_696),
.B(n_481),
.Y(n_763)
);

NOR2x1p5_ASAP7_75t_L g764 ( 
.A(n_590),
.B(n_501),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_595),
.B(n_501),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_709),
.B(n_643),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_522),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_634),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_622),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_625),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_650),
.A2(n_528),
.B1(n_522),
.B2(n_441),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_SL g773 ( 
.A(n_657),
.B(n_248),
.C(n_174),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_642),
.B(n_522),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_622),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_616),
.B(n_528),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_615),
.B(n_272),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_633),
.B(n_479),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_638),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_602),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_434),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_596),
.A2(n_436),
.B(n_457),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_611),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_636),
.B(n_434),
.Y(n_784)
);

NAND2x1p5_ASAP7_75t_L g785 ( 
.A(n_701),
.B(n_481),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_647),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_627),
.B(n_441),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_614),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_635),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_617),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_634),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_661),
.B(n_504),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_SL g793 ( 
.A(n_691),
.B(n_192),
.C(n_268),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_629),
.B(n_446),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_743),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_621),
.B(n_446),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_639),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_653),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_655),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_663),
.A2(n_453),
.B(n_454),
.C(n_457),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_672),
.B(n_450),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_672),
.B(n_450),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_664),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_673),
.B(n_461),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_685),
.B(n_461),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_686),
.B(n_463),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_727),
.B(n_458),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_689),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_743),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_SL g810 ( 
.A(n_657),
.B(n_238),
.C(n_176),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_630),
.B(n_594),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_693),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_606),
.B(n_458),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_613),
.B(n_463),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_694),
.B(n_698),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_647),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_712),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_681),
.B(n_458),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_714),
.B(n_469),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_720),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_631),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_658),
.B(n_469),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_652),
.B(n_473),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_646),
.A2(n_453),
.B1(n_454),
.B2(n_445),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_638),
.B(n_671),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_692),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_649),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_624),
.A2(n_445),
.B(n_438),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_730),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_743),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_688),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_640),
.B(n_473),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_665),
.B(n_480),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_624),
.A2(n_436),
.B(n_438),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_637),
.B(n_644),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_637),
.B(n_480),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_743),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_644),
.B(n_482),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_684),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_741),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_718),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_628),
.A2(n_496),
.B(n_497),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_690),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_700),
.B(n_588),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_692),
.B(n_504),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_659),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_593),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_660),
.B(n_545),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_597),
.B(n_527),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_587),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_670),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_665),
.B(n_482),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_700),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_597),
.B(n_527),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_651),
.A2(n_451),
.B1(n_455),
.B2(n_448),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_591),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_697),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_619),
.B(n_484),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_598),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_728),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_722),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_674),
.B(n_484),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_667),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_626),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_645),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_702),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_667),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_728),
.Y(n_868)
);

INVx5_ASAP7_75t_L g869 ( 
.A(n_711),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_620),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_618),
.B(n_485),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_SL g872 ( 
.A1(n_623),
.A2(n_236),
.B1(n_245),
.B2(n_247),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_589),
.B(n_504),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_695),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_648),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_676),
.B(n_485),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_648),
.B(n_532),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_683),
.B(n_707),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_716),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_609),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_723),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_725),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_669),
.B(n_527),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_656),
.B(n_486),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_656),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_679),
.A2(n_542),
.B1(n_532),
.B2(n_455),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_669),
.B(n_527),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_679),
.A2(n_542),
.B1(n_532),
.B2(n_455),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_708),
.B(n_486),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_717),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_721),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_608),
.B(n_527),
.Y(n_892)
);

OAI21xp33_ASAP7_75t_L g893 ( 
.A1(n_715),
.A2(n_448),
.B(n_451),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_710),
.B(n_491),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_733),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_680),
.A2(n_448),
.B1(n_455),
.B2(n_451),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_610),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_L g898 ( 
.A(n_706),
.B(n_530),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_735),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_662),
.Y(n_900)
);

AND2x2_ASAP7_75t_SL g901 ( 
.A(n_675),
.B(n_256),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_SL g902 ( 
.A(n_641),
.B(n_195),
.C(n_281),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_699),
.A2(n_542),
.B1(n_451),
.B2(n_448),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_654),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_729),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_742),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_604),
.B(n_530),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_703),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_605),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_584),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_706),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_699),
.B(n_530),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_682),
.B(n_491),
.Y(n_913)
);

INVxp33_ASAP7_75t_SL g914 ( 
.A(n_705),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_703),
.Y(n_915)
);

BUFx4f_ASAP7_75t_L g916 ( 
.A(n_704),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_706),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_736),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_736),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_706),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_706),
.B(n_495),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_705),
.A2(n_506),
.B1(n_540),
.B2(n_496),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_724),
.B(n_481),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_724),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_726),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_678),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_731),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_713),
.B(n_530),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_677),
.B(n_495),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_777),
.B(n_677),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_758),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_914),
.B(n_607),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_759),
.B(n_719),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_892),
.A2(n_666),
.B(n_928),
.C(n_754),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_746),
.B(n_675),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_752),
.B(n_732),
.C(n_737),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_746),
.A2(n_666),
.B(n_745),
.C(n_740),
.Y(n_937)
);

BUFx10_ASAP7_75t_L g938 ( 
.A(n_755),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_842),
.A2(n_628),
.B(n_739),
.Y(n_939)
);

AND3x1_ASAP7_75t_SL g940 ( 
.A(n_756),
.B(n_264),
.C(n_273),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_875),
.B(n_738),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_750),
.A2(n_744),
.B(n_739),
.C(n_583),
.Y(n_942)
);

AOI22x1_ASAP7_75t_L g943 ( 
.A1(n_764),
.A2(n_497),
.B1(n_499),
.B2(n_500),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_795),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_767),
.A2(n_734),
.B1(n_499),
.B2(n_540),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_885),
.B(n_668),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_878),
.B(n_668),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_749),
.A2(n_500),
.B(n_506),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_846),
.B(n_503),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_835),
.A2(n_503),
.B(n_536),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_774),
.Y(n_951)
);

INVx6_ASAP7_75t_L g952 ( 
.A(n_851),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_759),
.B(n_517),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_835),
.A2(n_517),
.B(n_535),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_811),
.B(n_246),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_891),
.B(n_534),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_795),
.Y(n_957)
);

INVx3_ASAP7_75t_SL g958 ( 
.A(n_860),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_767),
.B(n_539),
.Y(n_959)
);

CKINVDCx14_ASAP7_75t_R g960 ( 
.A(n_762),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_760),
.A2(n_539),
.B(n_243),
.C(n_235),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_864),
.B(n_3),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_877),
.A2(n_224),
.B(n_177),
.C(n_184),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_749),
.A2(n_815),
.B1(n_768),
.B2(n_917),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_831),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_868),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_791),
.B(n_257),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_916),
.A2(n_4),
.B(n_9),
.C(n_12),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_769),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_872),
.B(n_200),
.Y(n_970)
);

O2A1O1Ixp5_ASAP7_75t_L g971 ( 
.A1(n_916),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_788),
.B(n_15),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_863),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_925),
.A2(n_263),
.B(n_210),
.C(n_217),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_795),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_927),
.A2(n_258),
.B(n_214),
.C(n_545),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_768),
.A2(n_258),
.B(n_214),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_826),
.B(n_18),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_907),
.A2(n_276),
.B(n_207),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_861),
.B(n_545),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_757),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_826),
.B(n_18),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_881),
.B(n_20),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_771),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_921),
.A2(n_258),
.B(n_214),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_809),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_921),
.A2(n_545),
.B(n_481),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_861),
.B(n_545),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_897),
.A2(n_21),
.B(n_29),
.C(n_31),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_873),
.A2(n_481),
.B(n_276),
.C(n_207),
.Y(n_990)
);

BUFx4f_ASAP7_75t_L g991 ( 
.A(n_847),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_882),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_792),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_748),
.B(n_779),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_858),
.B(n_33),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_780),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_792),
.B(n_35),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_833),
.A2(n_852),
.B(n_900),
.C(n_910),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_836),
.A2(n_481),
.B(n_98),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_865),
.A2(n_36),
.B(n_40),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_836),
.A2(n_100),
.B(n_45),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_849),
.A2(n_41),
.B(n_276),
.C(n_207),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_838),
.A2(n_50),
.B(n_53),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_841),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_775),
.Y(n_1005)
);

AO22x1_ASAP7_75t_L g1006 ( 
.A1(n_853),
.A2(n_412),
.B1(n_276),
.B2(n_207),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_R g1007 ( 
.A(n_748),
.B(n_276),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_884),
.B(n_412),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_880),
.B(n_276),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_775),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_838),
.A2(n_58),
.B(n_80),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_779),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_867),
.B(n_412),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_825),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_793),
.A2(n_778),
.B(n_776),
.C(n_910),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_917),
.A2(n_412),
.B1(n_276),
.B2(n_207),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_840),
.A2(n_207),
.B(n_95),
.C(n_96),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_789),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_870),
.B(n_207),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_797),
.B(n_798),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_918),
.B(n_917),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_766),
.A2(n_126),
.B(n_133),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_799),
.B(n_136),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_929),
.A2(n_138),
.B(n_140),
.C(n_908),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_870),
.B(n_832),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_874),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_766),
.A2(n_822),
.B(n_801),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_854),
.A2(n_829),
.B(n_808),
.C(n_820),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_822),
.A2(n_801),
.B(n_802),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_783),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_774),
.Y(n_1031)
);

INVx3_ASAP7_75t_SL g1032 ( 
.A(n_905),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_845),
.B(n_751),
.Y(n_1033)
);

INVx6_ASAP7_75t_L g1034 ( 
.A(n_845),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_803),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_812),
.A2(n_817),
.B1(n_802),
.B2(n_919),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_904),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_SL g1038 ( 
.A(n_818),
.B(n_855),
.C(n_807),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_906),
.B(n_871),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_L g1040 ( 
.A(n_883),
.B(n_887),
.C(n_824),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_848),
.B(n_918),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_790),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_751),
.B(n_765),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_782),
.A2(n_834),
.B(n_828),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_915),
.A2(n_893),
.B(n_924),
.C(n_781),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_796),
.A2(n_800),
.B(n_824),
.C(n_773),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_784),
.B(n_823),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_844),
.B(n_909),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_828),
.A2(n_834),
.B(n_753),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_753),
.A2(n_920),
.B(n_911),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_775),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_909),
.B(n_816),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_810),
.B(n_902),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_850),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_782),
.A2(n_787),
.B(n_794),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_821),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_848),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_850),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_786),
.B(n_850),
.Y(n_1059)
);

AO32x1_ASAP7_75t_L g1060 ( 
.A1(n_855),
.A2(n_896),
.A3(n_827),
.B1(n_843),
.B2(n_866),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_964),
.A2(n_896),
.A3(n_814),
.B(n_862),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_939),
.A2(n_806),
.B(n_819),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_930),
.B(n_889),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_952),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_L g1065 ( 
.A(n_1051),
.B(n_765),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_932),
.B(n_894),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_SL g1067 ( 
.A1(n_998),
.A2(n_813),
.B(n_876),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_985),
.A2(n_805),
.B(n_804),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1034),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1050),
.A2(n_805),
.B(n_804),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_969),
.B(n_879),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_977),
.A2(n_954),
.B(n_950),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_1057),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_955),
.B(n_890),
.Y(n_1074)
);

AOI211x1_ASAP7_75t_L g1075 ( 
.A1(n_935),
.A2(n_912),
.B(n_913),
.C(n_903),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_931),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_933),
.B(n_913),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1025),
.B(n_890),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_SL g1079 ( 
.A1(n_992),
.A2(n_747),
.B1(n_772),
.B2(n_859),
.C(n_856),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_966),
.Y(n_1080)
);

AO21x1_ASAP7_75t_L g1081 ( 
.A1(n_1036),
.A2(n_922),
.B(n_888),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_996),
.Y(n_1082)
);

NOR4xp25_ASAP7_75t_L g1083 ( 
.A(n_1000),
.B(n_770),
.C(n_857),
.D(n_899),
.Y(n_1083)
);

AOI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_970),
.A2(n_856),
.B1(n_859),
.B2(n_839),
.C(n_895),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_1049),
.A2(n_886),
.B(n_926),
.Y(n_1085)
);

AO32x2_ASAP7_75t_L g1086 ( 
.A1(n_945),
.A2(n_869),
.A3(n_856),
.B1(n_859),
.B2(n_770),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1021),
.B(n_830),
.Y(n_1087)
);

CKINVDCx8_ASAP7_75t_R g1088 ( 
.A(n_1014),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_SL g1089 ( 
.A1(n_1047),
.A2(n_763),
.B(n_785),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1030),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_984),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1057),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_SL g1093 ( 
.A1(n_1028),
.A2(n_837),
.B(n_869),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_952),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_1029),
.A2(n_869),
.A3(n_926),
.B(n_923),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_1046),
.A2(n_926),
.B(n_763),
.Y(n_1096)
);

INVx8_ASAP7_75t_L g1097 ( 
.A(n_1004),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1037),
.B(n_785),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1039),
.B(n_973),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1055),
.A2(n_948),
.B(n_934),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_1048),
.B(n_938),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_959),
.A2(n_942),
.B(n_937),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1022),
.A2(n_1015),
.B(n_999),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_989),
.B(n_936),
.C(n_1053),
.Y(n_1104)
);

NAND3x1_ASAP7_75t_L g1105 ( 
.A(n_997),
.B(n_967),
.C(n_995),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_941),
.B(n_993),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1034),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1044),
.A2(n_943),
.B(n_1003),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_953),
.B(n_951),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_947),
.A2(n_1045),
.B(n_990),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1040),
.A2(n_1001),
.B(n_1011),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_987),
.A2(n_1002),
.B(n_1023),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_983),
.A2(n_962),
.B(n_961),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1017),
.A2(n_956),
.B(n_949),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1020),
.B(n_1032),
.Y(n_1115)
);

CKINVDCx11_ASAP7_75t_R g1116 ( 
.A(n_958),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_933),
.B(n_1018),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_944),
.Y(n_1118)
);

AND2x6_ASAP7_75t_L g1119 ( 
.A(n_951),
.B(n_1031),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_991),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_968),
.B(n_971),
.C(n_1038),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_946),
.A2(n_976),
.B(n_1024),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_991),
.B(n_1031),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_965),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1019),
.A2(n_1009),
.A3(n_1060),
.B(n_1016),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1035),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1052),
.A2(n_963),
.B(n_974),
.C(n_1059),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_938),
.B(n_1043),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1026),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_982),
.B(n_1058),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_978),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1043),
.B(n_1054),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1007),
.A2(n_1041),
.B(n_1008),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_953),
.B(n_1033),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_960),
.B(n_972),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_980),
.A2(n_988),
.B(n_994),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1042),
.B(n_1056),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_L g1138 ( 
.A1(n_1006),
.A2(n_1012),
.B(n_1013),
.C(n_940),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_944),
.A2(n_957),
.B(n_975),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1005),
.Y(n_1140)
);

AO21x1_ASAP7_75t_L g1141 ( 
.A1(n_1013),
.A2(n_1012),
.B(n_1010),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_975),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_SL g1143 ( 
.A1(n_986),
.A2(n_1028),
.B(n_1046),
.Y(n_1143)
);

NAND2x1_ASAP7_75t_L g1144 ( 
.A(n_1051),
.B(n_830),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_930),
.B(n_615),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1027),
.A2(n_761),
.B(n_898),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1049),
.A2(n_746),
.B(n_749),
.Y(n_1147)
);

AO21x1_ASAP7_75t_L g1148 ( 
.A1(n_1036),
.A2(n_935),
.B(n_1040),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_939),
.A2(n_842),
.B(n_979),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_964),
.A2(n_1027),
.A3(n_998),
.B(n_1029),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_SL g1151 ( 
.A1(n_998),
.A2(n_767),
.B(n_1036),
.Y(n_1151)
);

AOI31xp67_ASAP7_75t_L g1152 ( 
.A1(n_959),
.A2(n_892),
.A3(n_907),
.B(n_928),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_931),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_935),
.B(n_914),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_932),
.A2(n_588),
.B1(n_529),
.B2(n_560),
.C(n_914),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_930),
.B(n_615),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_979),
.A2(n_842),
.B(n_977),
.Y(n_1157)
);

OA22x2_ASAP7_75t_L g1158 ( 
.A1(n_933),
.A2(n_588),
.B1(n_623),
.B2(n_619),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_1049),
.A2(n_1044),
.B(n_939),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_932),
.A2(n_914),
.B(n_746),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_969),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_930),
.B(n_615),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_930),
.B(n_615),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_939),
.A2(n_842),
.B(n_979),
.Y(n_1164)
);

AOI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_935),
.A2(n_901),
.B(n_932),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_969),
.B(n_769),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_964),
.A2(n_1027),
.A3(n_998),
.B(n_1029),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_939),
.A2(n_842),
.B(n_979),
.Y(n_1168)
);

AOI31xp67_ASAP7_75t_L g1169 ( 
.A1(n_959),
.A2(n_892),
.A3(n_907),
.B(n_928),
.Y(n_1169)
);

NAND2x1_ASAP7_75t_L g1170 ( 
.A(n_1051),
.B(n_830),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_932),
.A2(n_914),
.B(n_428),
.C(n_433),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_SL g1172 ( 
.A1(n_932),
.A2(n_914),
.B(n_428),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_960),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_939),
.A2(n_842),
.B(n_979),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_935),
.B(n_914),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_939),
.A2(n_842),
.B(n_979),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_931),
.Y(n_1177)
);

NAND2x1_ASAP7_75t_L g1178 ( 
.A(n_1051),
.B(n_830),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_981),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_991),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_952),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1049),
.A2(n_746),
.B(n_749),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1027),
.A2(n_761),
.B(n_898),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1027),
.A2(n_761),
.B(n_898),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_932),
.A2(n_588),
.B1(n_529),
.B2(n_560),
.C(n_914),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_952),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_960),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1049),
.A2(n_746),
.B(n_749),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_939),
.A2(n_842),
.B(n_979),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1165),
.A2(n_1155),
.B(n_1185),
.C(n_1160),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1147),
.B(n_1182),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1072),
.A2(n_1100),
.B(n_1108),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1151),
.A2(n_1172),
.B(n_1121),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1172),
.A2(n_1121),
.B(n_1147),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1160),
.B(n_1162),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1166),
.B(n_1099),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_1085),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1164),
.A2(n_1174),
.B(n_1168),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1165),
.A2(n_1171),
.B(n_1113),
.C(n_1066),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1109),
.B(n_1098),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1182),
.A2(n_1188),
.B1(n_1105),
.B2(n_1154),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1188),
.B(n_1148),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1102),
.A2(n_1111),
.B(n_1113),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1175),
.A2(n_1158),
.B1(n_1063),
.B2(n_1163),
.Y(n_1205)
);

CKINVDCx11_ASAP7_75t_R g1206 ( 
.A(n_1116),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_1127),
.B(n_1075),
.C(n_1079),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1091),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1124),
.B(n_1088),
.Y(n_1209)
);

AOI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1143),
.A2(n_1180),
.B1(n_1173),
.B2(n_1135),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_R g1211 ( 
.A(n_1187),
.B(n_1173),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1126),
.B(n_1153),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1064),
.Y(n_1213)
);

OR3x4_ASAP7_75t_SL g1214 ( 
.A(n_1131),
.B(n_1097),
.C(n_1080),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1104),
.A2(n_1090),
.B1(n_1179),
.B2(n_1082),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1176),
.A2(n_1189),
.B(n_1146),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1183),
.A2(n_1068),
.B(n_1112),
.Y(n_1217)
);

AO21x1_ASAP7_75t_L g1218 ( 
.A1(n_1096),
.A2(n_1117),
.B(n_1101),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1062),
.A2(n_1114),
.B(n_1070),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_1073),
.B(n_1092),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1177),
.B(n_1071),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1084),
.A2(n_1130),
.B1(n_1074),
.B2(n_1137),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1083),
.A2(n_1141),
.A3(n_1086),
.B(n_1078),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1140),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1106),
.B(n_1107),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1159),
.A2(n_1085),
.B(n_1093),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1075),
.B(n_1061),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1086),
.A2(n_1152),
.A3(n_1169),
.B(n_1167),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1159),
.A2(n_1110),
.B(n_1136),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1094),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1122),
.A2(n_1110),
.B(n_1087),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1118),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1079),
.A2(n_1096),
.B(n_1067),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1077),
.A2(n_1101),
.B1(n_1115),
.B2(n_1119),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1128),
.A2(n_1138),
.B(n_1120),
.C(n_1123),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1077),
.A2(n_1119),
.B1(n_1122),
.B2(n_1132),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1181),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1097),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1092),
.A2(n_1065),
.B(n_1134),
.C(n_1139),
.Y(n_1239)
);

AOI221xp5_ASAP7_75t_L g1240 ( 
.A1(n_1097),
.A2(n_1186),
.B1(n_1133),
.B2(n_1089),
.C(n_1107),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1065),
.A2(n_1144),
.B1(n_1170),
.B2(n_1178),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1119),
.B(n_1142),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1119),
.B(n_1142),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_1118),
.A2(n_1061),
.B(n_1150),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1069),
.B(n_1129),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1167),
.B(n_1125),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1095),
.A2(n_1157),
.B(n_1072),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1125),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1146),
.A2(n_1184),
.B(n_1183),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1076),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1076),
.Y(n_1254)
);

O2A1O1Ixp5_ASAP7_75t_L g1255 ( 
.A1(n_1103),
.A2(n_1148),
.B(n_1111),
.C(n_1081),
.Y(n_1255)
);

AOI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1155),
.A2(n_1185),
.B1(n_932),
.B2(n_1172),
.C(n_1160),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1151),
.A2(n_1103),
.B(n_1040),
.Y(n_1257)
);

NOR2x1_ASAP7_75t_SL g1258 ( 
.A(n_1154),
.B(n_1036),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1117),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1172),
.A2(n_1171),
.B(n_1160),
.C(n_914),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1147),
.B(n_1182),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1180),
.B(n_1120),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1109),
.B(n_1098),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1158),
.A2(n_588),
.B1(n_872),
.B2(n_349),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1076),
.Y(n_1268)
);

CKINVDCx16_ASAP7_75t_R g1269 ( 
.A(n_1173),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1073),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1161),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1147),
.B(n_1182),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1151),
.A2(n_1103),
.B(n_1040),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1117),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1072),
.A2(n_1103),
.B(n_1100),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1160),
.B(n_1172),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1147),
.B(n_1182),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1161),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1076),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1165),
.A2(n_1185),
.B(n_1155),
.C(n_932),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1076),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1172),
.B(n_1185),
.C(n_1155),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1158),
.A2(n_588),
.B1(n_872),
.B2(n_349),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1117),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1155),
.A2(n_1185),
.B1(n_932),
.B2(n_914),
.Y(n_1291)
);

BUFx2_ASAP7_75t_R g1292 ( 
.A(n_1088),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1157),
.A2(n_1072),
.B(n_1149),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1160),
.B(n_1172),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1230),
.B(n_1237),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1257),
.B(n_1277),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1285),
.A2(n_1190),
.B(n_1260),
.C(n_1256),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1201),
.B(n_1250),
.Y(n_1298)
);

O2A1O1Ixp5_ASAP7_75t_L g1299 ( 
.A1(n_1257),
.A2(n_1277),
.B(n_1193),
.C(n_1194),
.Y(n_1299)
);

OA22x2_ASAP7_75t_L g1300 ( 
.A1(n_1205),
.A2(n_1291),
.B1(n_1193),
.B2(n_1194),
.Y(n_1300)
);

NOR2x1_ASAP7_75t_SL g1301 ( 
.A(n_1202),
.B(n_1207),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1288),
.A2(n_1256),
.B1(n_1294),
.B2(n_1281),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1255),
.A2(n_1204),
.B(n_1273),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1213),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1260),
.A2(n_1199),
.B(n_1233),
.C(n_1205),
.Y(n_1305)
);

AOI21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1203),
.A2(n_1262),
.B(n_1191),
.Y(n_1306)
);

O2A1O1Ixp5_ASAP7_75t_L g1307 ( 
.A1(n_1204),
.A2(n_1255),
.B(n_1202),
.C(n_1233),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1249),
.A2(n_1286),
.B(n_1274),
.Y(n_1308)
);

AOI21x1_ASAP7_75t_SL g1309 ( 
.A1(n_1191),
.A2(n_1282),
.B(n_1276),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1253),
.A2(n_1266),
.B(n_1261),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1262),
.A2(n_1276),
.B1(n_1282),
.B2(n_1267),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1264),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1212),
.B(n_1283),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1225),
.B(n_1200),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1267),
.A2(n_1289),
.B(n_1235),
.C(n_1227),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_SL g1316 ( 
.A1(n_1227),
.A2(n_1246),
.B(n_1214),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1258),
.A2(n_1239),
.B(n_1235),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1272),
.A2(n_1278),
.B(n_1275),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1240),
.A2(n_1242),
.B(n_1243),
.Y(n_1319)
);

AOI21x1_ASAP7_75t_SL g1320 ( 
.A1(n_1210),
.A2(n_1211),
.B(n_1206),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1290),
.B(n_1259),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1265),
.B(n_1279),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1269),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1289),
.A2(n_1222),
.B1(n_1234),
.B2(n_1236),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1232),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1292),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1208),
.A2(n_1252),
.B1(n_1268),
.B2(n_1287),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1238),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1224),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1254),
.B(n_1284),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1209),
.Y(n_1331)
);

O2A1O1Ixp5_ASAP7_75t_L g1332 ( 
.A1(n_1218),
.A2(n_1244),
.B(n_1231),
.C(n_1270),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1241),
.A2(n_1197),
.B(n_1263),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1223),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1220),
.A2(n_1244),
.B(n_1245),
.C(n_1251),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1215),
.A2(n_1248),
.B1(n_1280),
.B2(n_1219),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1293),
.A2(n_1247),
.B(n_1217),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1226),
.B(n_1228),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1192),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1198),
.B(n_1216),
.Y(n_1341)
);

INVx8_ASAP7_75t_L g1342 ( 
.A(n_1237),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1285),
.A2(n_1172),
.B(n_1190),
.C(n_1260),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1201),
.B(n_1250),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1257),
.A2(n_1277),
.B(n_1151),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1196),
.B(n_1195),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1190),
.A2(n_1285),
.B(n_1199),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1288),
.A2(n_1256),
.B1(n_1190),
.B2(n_1285),
.Y(n_1348)
);

OAI211xp5_ASAP7_75t_L g1349 ( 
.A1(n_1256),
.A2(n_1172),
.B(n_1193),
.C(n_1288),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1196),
.B(n_1221),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1285),
.A2(n_1172),
.B(n_1190),
.C(n_1260),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1288),
.A2(n_1256),
.B1(n_1190),
.B2(n_1285),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1191),
.B(n_1262),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1196),
.B(n_1221),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1191),
.B(n_1262),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1285),
.A2(n_1172),
.B(n_1190),
.C(n_1260),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1191),
.B(n_1262),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1201),
.B(n_1250),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1271),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1191),
.B(n_1262),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1257),
.A2(n_1277),
.B(n_1193),
.C(n_1148),
.Y(n_1361)
);

CKINVDCx6p67_ASAP7_75t_R g1362 ( 
.A(n_1206),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1191),
.B(n_1262),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1338),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1340),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1329),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1368)
);

OR2x6_ASAP7_75t_L g1369 ( 
.A(n_1345),
.B(n_1296),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1339),
.B(n_1303),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1308),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1357),
.B(n_1360),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1310),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1336),
.A2(n_1305),
.B(n_1334),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1360),
.B(n_1363),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1310),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1363),
.B(n_1299),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1318),
.A2(n_1337),
.B(n_1302),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1341),
.Y(n_1379)
);

AOI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1318),
.A2(n_1337),
.B(n_1302),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1300),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1330),
.B(n_1361),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1347),
.A2(n_1301),
.B(n_1311),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1325),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1307),
.B(n_1298),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1311),
.A2(n_1327),
.B(n_1348),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1332),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1348),
.A2(n_1352),
.B(n_1321),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1352),
.A2(n_1321),
.B(n_1315),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1335),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1344),
.B(n_1358),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1349),
.B(n_1297),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1359),
.B(n_1313),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1312),
.B(n_1300),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1333),
.A2(n_1324),
.B(n_1317),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1377),
.B(n_1346),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1370),
.B(n_1322),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1382),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1383),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1368),
.B(n_1350),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1369),
.B(n_1319),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1386),
.A2(n_1324),
.B1(n_1351),
.B2(n_1356),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1370),
.B(n_1354),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1365),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1370),
.B(n_1314),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1365),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1382),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1384),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1384),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1377),
.B(n_1343),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1392),
.A2(n_1326),
.B1(n_1331),
.B2(n_1323),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1371),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1377),
.B(n_1306),
.Y(n_1413)
);

NOR2x1_ASAP7_75t_SL g1414 ( 
.A(n_1383),
.B(n_1304),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1367),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1364),
.B(n_1316),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1375),
.B(n_1309),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1367),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_1413),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1406),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1406),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1402),
.B(n_1392),
.C(n_1377),
.Y(n_1422)
);

NAND2xp33_ASAP7_75t_R g1423 ( 
.A(n_1398),
.B(n_1394),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1415),
.Y(n_1424)
);

OAI222xp33_ASAP7_75t_L g1425 ( 
.A1(n_1402),
.A2(n_1381),
.B1(n_1410),
.B2(n_1398),
.C1(n_1407),
.C2(n_1394),
.Y(n_1425)
);

OAI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1410),
.A2(n_1381),
.B1(n_1387),
.B2(n_1394),
.C(n_1390),
.Y(n_1426)
);

NOR4xp25_ASAP7_75t_SL g1427 ( 
.A(n_1407),
.B(n_1390),
.C(n_1414),
.D(n_1379),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1415),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1405),
.B(n_1393),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1412),
.A2(n_1376),
.B(n_1373),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1414),
.B(n_1364),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1417),
.B(n_1396),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1400),
.Y(n_1433)
);

NAND2xp33_ASAP7_75t_SL g1434 ( 
.A(n_1417),
.B(n_1385),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1411),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1408),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1413),
.A2(n_1385),
.B1(n_1382),
.B2(n_1394),
.C(n_1366),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1412),
.A2(n_1380),
.B(n_1378),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1417),
.B(n_1385),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1401),
.A2(n_1383),
.B1(n_1386),
.B2(n_1381),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1412),
.A2(n_1376),
.B(n_1373),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_R g1442 ( 
.A(n_1408),
.B(n_1362),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1405),
.B(n_1393),
.Y(n_1443)
);

OAI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1399),
.A2(n_1381),
.B(n_1385),
.C(n_1382),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1396),
.A2(n_1386),
.B1(n_1389),
.B2(n_1388),
.C(n_1381),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1403),
.B(n_1375),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1404),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1409),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1399),
.A2(n_1395),
.B1(n_1383),
.B2(n_1381),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1418),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1409),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1430),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1447),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1447),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1438),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1420),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1422),
.B(n_1416),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1437),
.B(n_1405),
.Y(n_1458)
);

NOR2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1431),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1434),
.Y(n_1461)
);

NOR2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1399),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1438),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1424),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1431),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1411),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1420),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1429),
.B(n_1397),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1421),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1444),
.B(n_1399),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1429),
.B(n_1397),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1433),
.B(n_1386),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1441),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1445),
.B(n_1390),
.C(n_1387),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1431),
.B(n_1416),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1448),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1428),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1439),
.B(n_1386),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1432),
.B(n_1386),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1450),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1443),
.B(n_1397),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1443),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1474),
.B(n_1388),
.Y(n_1483)
);

NOR2x1_ASAP7_75t_L g1484 ( 
.A(n_1476),
.B(n_1383),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1461),
.B(n_1436),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1461),
.B(n_1436),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1476),
.B(n_1342),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1453),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1459),
.B(n_1431),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1474),
.B(n_1388),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1453),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1454),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1464),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1458),
.B(n_1436),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1458),
.B(n_1468),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1454),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1458),
.B(n_1451),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1452),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1478),
.B(n_1388),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1468),
.B(n_1451),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1478),
.B(n_1388),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1459),
.B(n_1440),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1476),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1464),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1478),
.B(n_1479),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1479),
.B(n_1446),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1456),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1468),
.B(n_1451),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_L g1509 ( 
.A(n_1476),
.B(n_1425),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1388),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1476),
.B(n_1342),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_SL g1512 ( 
.A(n_1457),
.B(n_1427),
.C(n_1440),
.Y(n_1512)
);

NAND5xp2_ASAP7_75t_L g1513 ( 
.A(n_1466),
.B(n_1449),
.C(n_1426),
.D(n_1380),
.E(n_1378),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1471),
.B(n_1450),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1457),
.A2(n_1423),
.B1(n_1387),
.B2(n_1366),
.C(n_1372),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1452),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1481),
.B(n_1442),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1456),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1467),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1467),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1469),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1469),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1466),
.A2(n_1395),
.B(n_1389),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1481),
.B(n_1403),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1493),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_L g1527 ( 
.A(n_1509),
.B(n_1455),
.C(n_1463),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1509),
.A2(n_1472),
.B(n_1470),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1504),
.B(n_1480),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1498),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1510),
.B(n_1477),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1503),
.B(n_1342),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1488),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1482),
.B(n_1471),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1491),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1491),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1492),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1516),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1485),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1494),
.B(n_1477),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1494),
.B(n_1471),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1482),
.B(n_1481),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1487),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1492),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1472),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1517),
.B(n_1460),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1513),
.A2(n_1395),
.B1(n_1389),
.B2(n_1374),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1511),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1496),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_L g1552 ( 
.A(n_1483),
.B(n_1455),
.C(n_1463),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1490),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1460),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1485),
.Y(n_1555)
);

AOI21xp33_ASAP7_75t_L g1556 ( 
.A1(n_1484),
.A2(n_1395),
.B(n_1389),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1497),
.B(n_1391),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1523),
.A2(n_1470),
.B(n_1475),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1484),
.B(n_1460),
.Y(n_1559)
);

OAI21xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1495),
.A2(n_1462),
.B(n_1475),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1536),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1540),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1548),
.A2(n_1512),
.B1(n_1553),
.B2(n_1502),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1515),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1526),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1540),
.B(n_1555),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1532),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1525),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1553),
.A2(n_1502),
.B1(n_1395),
.B2(n_1389),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1555),
.B(n_1495),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1486),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1514),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1549),
.B(n_1486),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1543),
.B(n_1500),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1514),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1529),
.B(n_1496),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1526),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1533),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1553),
.A2(n_1502),
.B1(n_1395),
.B2(n_1389),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1500),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1547),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1533),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1535),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1554),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1565),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1582),
.A2(n_1541),
.B(n_1554),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1568),
.A2(n_1527),
.B(n_1528),
.C(n_1556),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1581),
.B(n_1508),
.Y(n_1589)
);

OAI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1582),
.A2(n_1560),
.B(n_1558),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1565),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1581),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1563),
.A2(n_1560),
.B(n_1542),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1578),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1585),
.A2(n_1328),
.B1(n_1295),
.B2(n_1489),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1564),
.A2(n_1552),
.B(n_1538),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1585),
.A2(n_1559),
.B1(n_1552),
.B2(n_1546),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1569),
.A2(n_1499),
.B1(n_1501),
.B2(n_1537),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1508),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1578),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1573),
.B(n_1562),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1557),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1568),
.B(n_1489),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1579),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1589),
.B(n_1574),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1603),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1602),
.B(n_1567),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1592),
.B(n_1566),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1586),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1593),
.A2(n_1580),
.B1(n_1575),
.B2(n_1537),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_R g1612 ( 
.A1(n_1588),
.A2(n_1575),
.B1(n_1561),
.B2(n_1539),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1601),
.B(n_1587),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1596),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1591),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1608),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1614),
.A2(n_1596),
.B(n_1588),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1612),
.B(n_1597),
.C(n_1590),
.Y(n_1618)
);

NOR3xp33_ASAP7_75t_SL g1619 ( 
.A(n_1613),
.B(n_1609),
.C(n_1605),
.Y(n_1619)
);

NOR3xp33_ASAP7_75t_L g1620 ( 
.A(n_1613),
.B(n_1597),
.C(n_1595),
.Y(n_1620)
);

NAND4xp25_ASAP7_75t_L g1621 ( 
.A(n_1607),
.B(n_1603),
.C(n_1561),
.D(n_1570),
.Y(n_1621)
);

AOI322xp5_ASAP7_75t_L g1622 ( 
.A1(n_1611),
.A2(n_1598),
.A3(n_1604),
.B1(n_1594),
.B2(n_1600),
.C1(n_1530),
.C2(n_1551),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1611),
.A2(n_1577),
.B1(n_1531),
.B2(n_1579),
.C(n_1583),
.Y(n_1623)
);

OAI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1610),
.A2(n_1577),
.B1(n_1530),
.B2(n_1539),
.C(n_1551),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_SL g1625 ( 
.A(n_1606),
.B(n_1576),
.C(n_1572),
.Y(n_1625)
);

AOI222xp33_ASAP7_75t_L g1626 ( 
.A1(n_1618),
.A2(n_1615),
.B1(n_1584),
.B2(n_1583),
.C1(n_1559),
.C2(n_1473),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1617),
.A2(n_1584),
.B(n_1531),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1619),
.A2(n_1559),
.B(n_1538),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1616),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1620),
.B(n_1524),
.Y(n_1630)
);

AOI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1623),
.A2(n_1559),
.B(n_1550),
.C(n_1545),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1535),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1630),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1629),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1628),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1632),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1631),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_L g1638 ( 
.A(n_1626),
.B(n_1625),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1627),
.B(n_1622),
.C(n_1624),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_SL g1640 ( 
.A(n_1639),
.B(n_1427),
.C(n_1545),
.Y(n_1640)
);

OAI221xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1639),
.A2(n_1550),
.B1(n_1505),
.B2(n_1463),
.C(n_1455),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1634),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1638),
.A2(n_1463),
.B1(n_1455),
.B2(n_1505),
.C(n_1465),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1633),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1644),
.Y(n_1645)
);

NOR3xp33_ASAP7_75t_SL g1646 ( 
.A(n_1641),
.B(n_1635),
.C(n_1637),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1642),
.Y(n_1647)
);

OR2x6_ASAP7_75t_L g1648 ( 
.A(n_1647),
.B(n_1636),
.Y(n_1648)
);

OAI32xp33_ASAP7_75t_L g1649 ( 
.A1(n_1648),
.A2(n_1643),
.A3(n_1646),
.B1(n_1645),
.B2(n_1640),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1649),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1649),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1650),
.B(n_1507),
.Y(n_1652)
);

NAND2x1_ASAP7_75t_SL g1653 ( 
.A(n_1651),
.B(n_1489),
.Y(n_1653)
);

XNOR2xp5_ASAP7_75t_L g1654 ( 
.A(n_1652),
.B(n_1462),
.Y(n_1654)
);

AOI21xp33_ASAP7_75t_L g1655 ( 
.A1(n_1653),
.A2(n_1463),
.B(n_1455),
.Y(n_1655)
);

XNOR2x2_ASAP7_75t_L g1656 ( 
.A(n_1654),
.B(n_1507),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1655),
.B1(n_1518),
.B2(n_1522),
.Y(n_1657)
);

AOI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1520),
.B(n_1522),
.Y(n_1658)
);

AOI22x1_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1519),
.B1(n_1518),
.B2(n_1521),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1659),
.A2(n_1519),
.B1(n_1521),
.B2(n_1520),
.C(n_1506),
.Y(n_1660)
);

AOI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1660),
.A2(n_1320),
.B(n_1506),
.C(n_1465),
.Y(n_1661)
);


endmodule