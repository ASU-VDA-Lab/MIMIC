module fake_ariane_1662_n_176 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_176);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_176;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_128;
wire n_105;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVxp33_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_37),
.C(n_40),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_4),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_6),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_7),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_21),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

AOI21x1_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_52),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_48),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_52),
.B(n_49),
.C(n_43),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_50),
.B(n_43),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_42),
.B(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_42),
.B(n_41),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_65),
.B(n_58),
.C(n_71),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_10),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_11),
.B(n_12),
.C(n_17),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_31),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_24),
.B(n_26),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_64),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_63),
.B1(n_62),
.B2(n_70),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_75),
.Y(n_95)
);

OR2x6_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_74),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_70),
.B(n_73),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_70),
.B(n_74),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_63),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_91),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_80),
.B(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_103),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_94),
.C(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_96),
.B1(n_98),
.B2(n_104),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_93),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_96),
.C(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_96),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_96),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_79),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_86),
.C(n_74),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_73),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_122),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_108),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_72),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_72),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_127),
.B(n_132),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_128),
.C(n_130),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_133),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_134),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_88),
.C(n_81),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_87),
.C(n_131),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_141),
.B1(n_66),
.B2(n_100),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_145),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_143),
.C(n_148),
.Y(n_162)
);

AOI211x1_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_83),
.B(n_100),
.C(n_110),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_159),
.Y(n_164)
);

NAND2x1p5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_112),
.Y(n_167)
);

OAI221xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.C(n_157),
.Y(n_168)
);

OAI222xp33_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_157),
.B1(n_108),
.B2(n_107),
.C1(n_105),
.C2(n_70),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_112),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_107),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_105),
.B1(n_101),
.B2(n_112),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_166),
.B(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_105),
.B1(n_101),
.B2(n_70),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_173),
.B(n_170),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_174),
.B1(n_172),
.B2(n_169),
.C(n_105),
.Y(n_176)
);


endmodule