module real_aes_7451_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_755;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_1), .A2(n_146), .B(n_149), .C(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_2), .A2(n_174), .B(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g502 ( .A(n_3), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_4), .B(n_185), .Y(n_184) );
AOI21xp33_ASAP7_75t_L g479 ( .A1(n_5), .A2(n_174), .B(n_480), .Y(n_479) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g249 ( .A(n_7), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_41), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_9), .A2(n_273), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_10), .B(n_158), .Y(n_226) );
INVx1_ASAP7_75t_L g484 ( .A(n_11), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_12), .B(n_179), .Y(n_535) );
INVx1_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
INVx1_ASAP7_75t_L g547 ( .A(n_14), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_15), .A2(n_193), .B(n_234), .C(n_236), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_16), .B(n_185), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_17), .B(n_473), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_18), .B(n_174), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_19), .B(n_281), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_20), .A2(n_179), .B(n_210), .C(n_213), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_21), .B(n_185), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_22), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_23), .A2(n_212), .B(n_236), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_24), .B(n_158), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_25), .Y(n_140) );
INVx1_ASAP7_75t_L g191 ( .A(n_26), .Y(n_191) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_28), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_29), .B(n_158), .Y(n_503) );
INVx1_ASAP7_75t_L g278 ( .A(n_30), .Y(n_278) );
INVx1_ASAP7_75t_L g492 ( .A(n_31), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_32), .A2(n_122), .B1(n_123), .B2(n_448), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_32), .Y(n_448) );
INVx2_ASAP7_75t_L g144 ( .A(n_33), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_34), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_35), .B(n_453), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_36), .A2(n_179), .B(n_180), .C(n_182), .Y(n_178) );
INVxp67_ASAP7_75t_L g279 ( .A(n_37), .Y(n_279) );
CKINVDCx14_ASAP7_75t_R g176 ( .A(n_38), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_39), .A2(n_149), .B(n_190), .C(n_197), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_40), .A2(n_146), .B(n_149), .C(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_42), .A2(n_104), .B1(n_115), .B2(n_756), .Y(n_103) );
INVx1_ASAP7_75t_L g491 ( .A(n_43), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_44), .A2(n_52), .B1(n_446), .B2(n_447), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_44), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_45), .A2(n_65), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_45), .Y(n_749) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_46), .A2(n_746), .B1(n_747), .B2(n_750), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_46), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_47), .A2(n_160), .B(n_247), .C(n_248), .Y(n_246) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_48), .A2(n_456), .B1(n_744), .B2(n_745), .C1(n_751), .C2(n_752), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_49), .B(n_158), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_50), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_51), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_52), .Y(n_446) );
INVx1_ASAP7_75t_L g208 ( .A(n_53), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_54), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_55), .B(n_174), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_56), .A2(n_149), .B1(n_213), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_57), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_58), .Y(n_499) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_59), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_60), .A2(n_182), .B(n_247), .C(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_61), .Y(n_527) );
INVx1_ASAP7_75t_L g481 ( .A(n_62), .Y(n_481) );
INVx1_ASAP7_75t_L g147 ( .A(n_63), .Y(n_147) );
INVx1_ASAP7_75t_L g137 ( .A(n_64), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_65), .Y(n_748) );
INVx1_ASAP7_75t_SL g181 ( .A(n_66), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_68), .B(n_185), .Y(n_215) );
INVx1_ASAP7_75t_L g153 ( .A(n_69), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_SL g472 ( .A1(n_70), .A2(n_182), .B(n_473), .C(n_474), .Y(n_472) );
INVxp67_ASAP7_75t_L g475 ( .A(n_71), .Y(n_475) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_73), .A2(n_174), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_74), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_75), .A2(n_174), .B(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_76), .Y(n_495) );
INVx1_ASAP7_75t_L g521 ( .A(n_77), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_78), .A2(n_273), .B(n_274), .Y(n_272) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_79), .Y(n_188) );
INVx1_ASAP7_75t_L g232 ( .A(n_80), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_81), .A2(n_146), .B(n_149), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_82), .A2(n_174), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g235 ( .A(n_83), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_84), .B(n_192), .Y(n_515) );
INVx2_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx1_ASAP7_75t_L g225 ( .A(n_86), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_87), .B(n_473), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_88), .A2(n_146), .B(n_149), .C(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
OR2x2_ASAP7_75t_L g451 ( .A(n_89), .B(n_111), .Y(n_451) );
OR2x2_ASAP7_75t_L g742 ( .A(n_89), .B(n_112), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_90), .A2(n_149), .B(n_152), .C(n_162), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_91), .B(n_167), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_92), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_93), .A2(n_146), .B(n_149), .C(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_94), .Y(n_539) );
INVx1_ASAP7_75t_L g471 ( .A(n_95), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_96), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_97), .B(n_192), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_98), .B(n_133), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_99), .B(n_133), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_100), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g211 ( .A(n_101), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_102), .A2(n_174), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g756 ( .A(n_105), .Y(n_756) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g751 ( .A(n_108), .Y(n_751) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g459 ( .A(n_110), .B(n_112), .Y(n_459) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_454), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g755 ( .A(n_117), .Y(n_755) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_449), .B(n_452), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_445), .Y(n_123) );
INVx3_ASAP7_75t_L g743 ( .A(n_124), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_124), .A2(n_458), .B1(n_741), .B2(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_400), .Y(n_124) );
NOR4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_337), .C(n_371), .D(n_387), .Y(n_125) );
NAND4xp25_ASAP7_75t_SL g126 ( .A(n_127), .B(n_263), .C(n_301), .D(n_317), .Y(n_126) );
AOI222xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_200), .B1(n_238), .B2(n_251), .C1(n_256), .C2(n_262), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI31xp33_ASAP7_75t_L g433 ( .A1(n_129), .A2(n_434), .A3(n_435), .B(n_437), .Y(n_433) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_168), .Y(n_129) );
AND2x2_ASAP7_75t_L g408 ( .A(n_130), .B(n_170), .Y(n_408) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g255 ( .A(n_131), .Y(n_255) );
AND2x2_ASAP7_75t_L g262 ( .A(n_131), .B(n_186), .Y(n_262) );
AND2x2_ASAP7_75t_L g322 ( .A(n_131), .B(n_171), .Y(n_322) );
AO21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_164), .Y(n_131) );
INVx3_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_132), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_132), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_SL g517 ( .A(n_132), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_133), .A2(n_469), .B(n_476), .Y(n_468) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g271 ( .A(n_134), .Y(n_271) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_135), .B(n_136), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_148), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_141), .A2(n_167), .B(n_188), .C(n_189), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_141), .A2(n_222), .B(n_223), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_141), .A2(n_163), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_141), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_141), .A2(n_521), .B(n_522), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
AND2x4_ASAP7_75t_L g174 ( .A(n_142), .B(n_146), .Y(n_174) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g196 ( .A(n_143), .Y(n_196) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx1_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
INVx1_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
INVx3_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
INVx1_ASAP7_75t_L g473 ( .A(n_145), .Y(n_473) );
INVx4_ASAP7_75t_SL g163 ( .A(n_146), .Y(n_163) );
BUFx3_ASAP7_75t_L g197 ( .A(n_146), .Y(n_197) );
INVx5_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx3_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_150), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .C(n_159), .Y(n_152) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_159), .B(n_225), .C(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_155), .A2(n_156), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
INVx4_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
INVx2_ASAP7_75t_L g247 ( .A(n_158), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_159), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_159), .A2(n_524), .B(n_525), .Y(n_523) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_163), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g207 ( .A1(n_163), .A2(n_177), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_163), .A2(n_177), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_163), .A2(n_177), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g274 ( .A1(n_163), .A2(n_177), .B(n_275), .C(n_276), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_163), .A2(n_177), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_163), .A2(n_177), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_163), .A2(n_177), .B(n_544), .C(n_545), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g281 ( .A(n_166), .Y(n_281) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_166), .A2(n_531), .B(n_538), .Y(n_530) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_167), .A2(n_243), .B(n_250), .Y(n_242) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_167), .A2(n_542), .B(n_548), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_168), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_169), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_169), .B(n_266), .Y(n_312) );
AND2x2_ASAP7_75t_L g405 ( .A(n_169), .B(n_345), .Y(n_405) );
OAI321xp33_ASAP7_75t_L g439 ( .A1(n_169), .A2(n_255), .A3(n_412), .B1(n_440), .B2(n_442), .C(n_443), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_169), .B(n_241), .C(n_352), .D(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_186), .Y(n_169) );
AND2x2_ASAP7_75t_L g307 ( .A(n_170), .B(n_253), .Y(n_307) );
AND2x2_ASAP7_75t_L g326 ( .A(n_170), .B(n_255), .Y(n_326) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g254 ( .A(n_171), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g282 ( .A(n_171), .B(n_186), .Y(n_282) );
AND2x2_ASAP7_75t_L g368 ( .A(n_171), .B(n_253), .Y(n_368) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_184), .Y(n_171) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_172), .A2(n_206), .B(n_215), .Y(n_205) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_172), .A2(n_230), .B(n_237), .Y(n_229) );
BUFx2_ASAP7_75t_L g273 ( .A(n_174), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_179), .B(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_183), .Y(n_536) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_185), .A2(n_479), .B(n_485), .Y(n_478) );
INVx3_ASAP7_75t_SL g253 ( .A(n_186), .Y(n_253) );
AND2x2_ASAP7_75t_L g300 ( .A(n_186), .B(n_287), .Y(n_300) );
OR2x2_ASAP7_75t_L g333 ( .A(n_186), .B(n_255), .Y(n_333) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_186), .Y(n_340) );
AND2x2_ASAP7_75t_L g369 ( .A(n_186), .B(n_254), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_186), .B(n_342), .Y(n_384) );
AND2x2_ASAP7_75t_L g416 ( .A(n_186), .B(n_408), .Y(n_416) );
AND2x2_ASAP7_75t_L g425 ( .A(n_186), .B(n_267), .Y(n_425) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_198), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_194), .C(n_195), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_192), .A2(n_212), .B1(n_278), .B2(n_279), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_192), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
INVx5_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_193), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_193), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_193), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_196), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_216), .Y(n_201) );
INVx1_ASAP7_75t_SL g393 ( .A(n_202), .Y(n_393) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g258 ( .A(n_203), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g240 ( .A(n_204), .B(n_218), .Y(n_240) );
AND2x2_ASAP7_75t_L g329 ( .A(n_204), .B(n_242), .Y(n_329) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g299 ( .A(n_205), .B(n_229), .Y(n_299) );
OR2x2_ASAP7_75t_L g310 ( .A(n_205), .B(n_242), .Y(n_310) );
AND2x2_ASAP7_75t_L g336 ( .A(n_205), .B(n_242), .Y(n_336) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_205), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_212), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_212), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g504 ( .A(n_213), .Y(n_504) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_216), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_216), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g309 ( .A(n_217), .B(n_310), .Y(n_309) );
AOI322xp5_ASAP7_75t_L g395 ( .A1(n_217), .A2(n_299), .A3(n_305), .B1(n_336), .B2(n_386), .C1(n_396), .C2(n_398), .Y(n_395) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_229), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_218), .B(n_241), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_218), .B(n_242), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_218), .B(n_259), .Y(n_316) );
AND2x2_ASAP7_75t_L g370 ( .A(n_218), .B(n_336), .Y(n_370) );
INVx1_ASAP7_75t_L g374 ( .A(n_218), .Y(n_374) );
AND2x2_ASAP7_75t_L g386 ( .A(n_218), .B(n_229), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_218), .B(n_258), .Y(n_418) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g283 ( .A(n_219), .B(n_229), .Y(n_283) );
BUFx3_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
AND3x2_ASAP7_75t_L g379 ( .A(n_219), .B(n_359), .C(n_380), .Y(n_379) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_227), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_220), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_220), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_220), .B(n_539), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g239 ( .A(n_229), .B(n_240), .C(n_241), .Y(n_239) );
INVx1_ASAP7_75t_SL g259 ( .A(n_229), .Y(n_259) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_229), .Y(n_364) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g358 ( .A(n_240), .B(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g365 ( .A(n_240), .Y(n_365) );
AND2x2_ASAP7_75t_L g403 ( .A(n_241), .B(n_381), .Y(n_403) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx3_ASAP7_75t_L g284 ( .A(n_242), .Y(n_284) );
AND2x2_ASAP7_75t_L g359 ( .A(n_242), .B(n_259), .Y(n_359) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OR2x2_ASAP7_75t_L g303 ( .A(n_253), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g422 ( .A(n_253), .B(n_322), .Y(n_422) );
AND2x2_ASAP7_75t_L g436 ( .A(n_253), .B(n_255), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_254), .B(n_267), .Y(n_377) );
AND2x2_ASAP7_75t_L g424 ( .A(n_254), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g287 ( .A(n_255), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g304 ( .A(n_255), .B(n_267), .Y(n_304) );
INVx1_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
AND2x2_ASAP7_75t_L g345 ( .A(n_255), .B(n_267), .Y(n_345) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_257), .A2(n_388), .B1(n_392), .B2(n_394), .C(n_395), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x2_ASAP7_75t_L g291 ( .A(n_258), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_261), .B(n_298), .Y(n_441) );
AOI322xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_283), .A3(n_284), .B1(n_285), .B2(n_291), .C1(n_293), .C2(n_300), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_282), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_266), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_266), .B(n_332), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_266), .A2(n_282), .B(n_356), .C(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_266), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_266), .B(n_326), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_266), .B(n_408), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_266), .B(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_267), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_267), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g397 ( .A(n_267), .B(n_284), .Y(n_397) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B(n_280), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_269), .A2(n_289), .B(n_290), .Y(n_288) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_269), .A2(n_520), .B(n_526), .Y(n_519) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AOI21xp5_ASAP7_75t_SL g511 ( .A1(n_270), .A2(n_512), .B(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_271), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_271), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_271), .A2(n_498), .B(n_505), .Y(n_497) );
INVx1_ASAP7_75t_L g289 ( .A(n_272), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_280), .Y(n_290) );
INVx1_ASAP7_75t_L g372 ( .A(n_282), .Y(n_372) );
OAI31xp33_ASAP7_75t_L g382 ( .A1(n_282), .A2(n_307), .A3(n_383), .B(n_385), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_282), .B(n_288), .Y(n_434) );
INVx1_ASAP7_75t_SL g295 ( .A(n_283), .Y(n_295) );
AND2x2_ASAP7_75t_L g328 ( .A(n_283), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g409 ( .A(n_283), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g294 ( .A(n_284), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
AND2x2_ASAP7_75t_L g346 ( .A(n_284), .B(n_299), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_284), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g438 ( .A(n_284), .B(n_386), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_286), .B(n_356), .Y(n_429) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g343 ( .A(n_288), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
OAI211xp5_ASAP7_75t_SL g337 ( .A1(n_295), .A2(n_338), .B(n_344), .C(n_360), .Y(n_337) );
OR2x2_ASAP7_75t_L g412 ( .A(n_295), .B(n_393), .Y(n_412) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g349 ( .A(n_297), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_297), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g318 ( .A(n_299), .B(n_319), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B(n_308), .C(n_311), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g352 ( .A(n_304), .Y(n_352) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_307), .B(n_345), .Y(n_350) );
INVx1_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g315 ( .A(n_310), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g348 ( .A(n_310), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g410 ( .A(n_310), .Y(n_410) );
AOI21xp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_313), .B(n_315), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_313), .A2(n_324), .B(n_327), .Y(n_323) );
AOI211xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B(n_323), .C(n_330), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_318), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_321), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g334 ( .A(n_322), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_324), .A2(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_329), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g354 ( .A(n_329), .Y(n_354) );
AOI21xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_334), .B(n_335), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g385 ( .A(n_336), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_342), .B(n_368), .Y(n_394) );
AND2x2_ASAP7_75t_L g407 ( .A(n_342), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g421 ( .A(n_342), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g431 ( .A(n_342), .B(n_369), .Y(n_431) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B(n_347), .C(n_355), .Y(n_344) );
INVx1_ASAP7_75t_L g391 ( .A(n_345), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B1(n_351), .B2(n_353), .Y(n_347) );
OR2x2_ASAP7_75t_L g353 ( .A(n_349), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_349), .B(n_410), .Y(n_432) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g426 ( .A(n_359), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_366), .B1(n_369), .B2(n_370), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g444 ( .A(n_364), .Y(n_444) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g390 ( .A(n_368), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_373), .B(n_375), .C(n_382), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_390), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR5xp2_ASAP7_75t_L g400 ( .A(n_401), .B(n_419), .C(n_427), .D(n_433), .E(n_439), .Y(n_400) );
OAI211xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_404), .B(n_406), .C(n_413), .Y(n_401) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B(n_411), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_416), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B(n_426), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g442 ( .A(n_422), .Y(n_442) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B(n_432), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_451), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g454 ( .A1(n_452), .A2(n_455), .B(n_755), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B1(n_741), .B2(n_743), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g754 ( .A(n_460), .Y(n_754) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND4x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_659), .C(n_706), .D(n_726), .Y(n_461) );
NOR3xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_589), .C(n_614), .Y(n_462) );
OAI211xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_507), .B(n_549), .C(n_579), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_486), .Y(n_465) );
INVx3_ASAP7_75t_SL g631 ( .A(n_466), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_466), .B(n_562), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_466), .B(n_496), .Y(n_712) );
AND2x2_ASAP7_75t_L g735 ( .A(n_466), .B(n_601), .Y(n_735) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g553 ( .A(n_468), .B(n_478), .Y(n_553) );
INVx3_ASAP7_75t_L g566 ( .A(n_468), .Y(n_566) );
AND2x2_ASAP7_75t_L g571 ( .A(n_468), .B(n_477), .Y(n_571) );
OR2x2_ASAP7_75t_L g622 ( .A(n_468), .B(n_563), .Y(n_622) );
BUFx2_ASAP7_75t_L g642 ( .A(n_468), .Y(n_642) );
AND2x2_ASAP7_75t_L g652 ( .A(n_468), .B(n_563), .Y(n_652) );
AND2x2_ASAP7_75t_L g658 ( .A(n_468), .B(n_487), .Y(n_658) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_478), .B(n_563), .Y(n_577) );
INVx2_ASAP7_75t_L g587 ( .A(n_478), .Y(n_587) );
AND2x2_ASAP7_75t_L g600 ( .A(n_478), .B(n_566), .Y(n_600) );
OR2x2_ASAP7_75t_L g611 ( .A(n_478), .B(n_563), .Y(n_611) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_478), .B(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g669 ( .A(n_478), .Y(n_669) );
AND2x2_ASAP7_75t_L g715 ( .A(n_478), .B(n_487), .Y(n_715) );
INVx3_ASAP7_75t_SL g588 ( .A(n_486), .Y(n_588) );
OR2x2_ASAP7_75t_L g641 ( .A(n_486), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
INVx3_ASAP7_75t_L g563 ( .A(n_487), .Y(n_563) );
AND2x2_ASAP7_75t_L g630 ( .A(n_487), .B(n_497), .Y(n_630) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_487), .Y(n_698) );
AOI33xp33_ASAP7_75t_L g702 ( .A1(n_487), .A2(n_631), .A3(n_638), .B1(n_647), .B2(n_703), .B3(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_496), .B(n_566), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_496), .B(n_626), .C(n_628), .Y(n_625) );
AND2x2_ASAP7_75t_L g651 ( .A(n_496), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_496), .B(n_658), .Y(n_661) );
AND2x2_ASAP7_75t_L g714 ( .A(n_496), .B(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
OR2x2_ASAP7_75t_L g664 ( .A(n_497), .B(n_563), .Y(n_664) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_528), .Y(n_507) );
AOI32xp33_ASAP7_75t_L g615 ( .A1(n_508), .A2(n_616), .A3(n_618), .B1(n_620), .B2(n_623), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_508), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g718 ( .A(n_508), .Y(n_718) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g650 ( .A(n_509), .B(n_634), .Y(n_650) );
AND2x2_ASAP7_75t_L g670 ( .A(n_509), .B(n_596), .Y(n_670) );
AND2x2_ASAP7_75t_L g738 ( .A(n_509), .B(n_656), .Y(n_738) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
INVx3_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
AND2x2_ASAP7_75t_L g573 ( .A(n_510), .B(n_557), .Y(n_573) );
OR2x2_ASAP7_75t_L g578 ( .A(n_510), .B(n_556), .Y(n_578) );
INVx1_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
AND2x2_ASAP7_75t_L g593 ( .A(n_510), .B(n_567), .Y(n_593) );
AND2x2_ASAP7_75t_L g595 ( .A(n_510), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_510), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g648 ( .A(n_510), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_510), .B(n_733), .Y(n_732) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_517), .Y(n_510) );
INVx2_ASAP7_75t_L g557 ( .A(n_519), .Y(n_557) );
AND2x2_ASAP7_75t_L g603 ( .A(n_519), .B(n_529), .Y(n_603) );
AND2x2_ASAP7_75t_L g613 ( .A(n_519), .B(n_541), .Y(n_613) );
INVx2_ASAP7_75t_L g733 ( .A(n_528), .Y(n_733) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_529), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g574 ( .A(n_529), .Y(n_574) );
AND2x2_ASAP7_75t_L g618 ( .A(n_529), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g634 ( .A(n_529), .B(n_597), .Y(n_634) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
AND2x2_ASAP7_75t_L g596 ( .A(n_530), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g647 ( .A(n_530), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_530), .B(n_557), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
AND2x2_ASAP7_75t_L g558 ( .A(n_540), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g619 ( .A(n_540), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_540), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g656 ( .A(n_540), .Y(n_656) );
INVx1_ASAP7_75t_L g689 ( .A(n_540), .Y(n_689) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g567 ( .A(n_541), .B(n_557), .Y(n_567) );
INVx1_ASAP7_75t_L g597 ( .A(n_541), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B1(n_560), .B2(n_567), .C(n_568), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_551), .B(n_571), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_551), .B(n_634), .Y(n_711) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_553), .B(n_601), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_553), .B(n_562), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_553), .B(n_576), .Y(n_705) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
AND2x2_ASAP7_75t_L g602 ( .A(n_558), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g680 ( .A(n_558), .Y(n_680) );
AND2x2_ASAP7_75t_L g612 ( .A(n_559), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_559), .B(n_582), .Y(n_628) );
AND2x2_ASAP7_75t_L g692 ( .A(n_559), .B(n_618), .Y(n_692) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g601 ( .A(n_563), .B(n_570), .Y(n_601) );
AND2x2_ASAP7_75t_L g697 ( .A(n_564), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_566), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_567), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_567), .B(n_574), .Y(n_662) );
AND2x2_ASAP7_75t_L g682 ( .A(n_567), .B(n_582), .Y(n_682) );
AND2x2_ASAP7_75t_L g703 ( .A(n_567), .B(n_647), .Y(n_703) );
OAI32xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .A3(n_574), .B1(n_575), .B2(n_578), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_SL g576 ( .A(n_570), .Y(n_576) );
NAND2x1_ASAP7_75t_L g617 ( .A(n_570), .B(n_600), .Y(n_617) );
OR2x2_ASAP7_75t_L g621 ( .A(n_570), .B(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_570), .B(n_669), .Y(n_722) );
INVx1_ASAP7_75t_L g590 ( .A(n_571), .Y(n_590) );
OAI221xp5_ASAP7_75t_SL g708 ( .A1(n_572), .A2(n_663), .B1(n_709), .B2(n_712), .C(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g580 ( .A(n_573), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g623 ( .A(n_573), .B(n_596), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_573), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g701 ( .A(n_573), .B(n_634), .Y(n_701) );
INVxp67_ASAP7_75t_L g637 ( .A(n_574), .Y(n_637) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g707 ( .A(n_576), .B(n_694), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_576), .B(n_657), .Y(n_730) );
INVx1_ASAP7_75t_L g605 ( .A(n_578), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_578), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g723 ( .A(n_578), .B(n_724), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_583), .B(n_586), .Y(n_579) );
AND2x2_ASAP7_75t_L g592 ( .A(n_581), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g676 ( .A(n_585), .B(n_596), .Y(n_676) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AND2x2_ASAP7_75t_L g694 ( .A(n_587), .B(n_652), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_587), .B(n_651), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_588), .B(n_600), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_594), .C(n_604), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_590), .A2(n_625), .B1(n_629), .B2(n_632), .C(n_635), .Y(n_624) );
AOI31xp33_ASAP7_75t_L g719 ( .A1(n_590), .A2(n_720), .A3(n_721), .B(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_598), .B1(n_600), .B2(n_602), .Y(n_594) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g720 ( .A(n_600), .Y(n_720) );
INVx1_ASAP7_75t_L g683 ( .A(n_601), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_603), .A2(n_727), .B(n_729), .C(n_731), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_608), .B2(n_612), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_609), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g699 ( .A1(n_611), .A2(n_645), .B1(n_664), .B2(n_700), .C(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g695 ( .A(n_612), .Y(n_695) );
INVx1_ASAP7_75t_L g649 ( .A(n_613), .Y(n_649) );
NAND3xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_624), .C(n_639), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_616), .A2(n_666), .B(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_618), .B(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g725 ( .A(n_619), .Y(n_725) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g663 ( .A(n_626), .B(n_646), .Y(n_663) );
INVx1_ASAP7_75t_L g638 ( .A(n_627), .Y(n_638) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g636 ( .A(n_630), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_630), .B(n_668), .Y(n_667) );
NOR4xp25_ASAP7_75t_L g635 ( .A(n_631), .B(n_636), .C(n_637), .D(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_644), .B1(n_650), .B2(n_651), .C1(n_653), .C2(n_657), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g737 ( .A(n_641), .Y(n_737) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_653), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g713 ( .A1(n_658), .A2(n_714), .B(n_716), .Y(n_713) );
NOR4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_671), .C(n_684), .D(n_699), .Y(n_659) );
OAI221xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B1(n_663), .B2(n_664), .C(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g740 ( .A(n_661), .Y(n_740) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_668), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
OAI222xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .B1(n_677), .B2(n_678), .C1(n_681), .C2(n_683), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_676), .A2(n_707), .B(n_708), .C(n_719), .Y(n_706) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
OAI222xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_690), .B1(n_691), .B2(n_693), .C1(n_695), .C2(n_696), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_701), .A2(n_704), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI211xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_734), .B(n_736), .C(n_739), .Y(n_731) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule