module fake_jpeg_30859_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_73),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_1),
.B(n_2),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_75),
.B(n_60),
.C(n_64),
.Y(n_91)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_53),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_66),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_87),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_66),
.B1(n_65),
.B2(n_59),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_79),
.B1(n_68),
.B2(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_96),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_58),
.B1(n_65),
.B2(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_69),
.B1(n_63),
.B2(n_55),
.Y(n_102)
);

NAND2x1_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_63),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_105),
.B1(n_115),
.B2(n_11),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_110),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_113),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_63),
.B1(n_69),
.B2(n_72),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_114),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_71),
.B(n_51),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_42),
.B(n_22),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_57),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_62),
.B1(n_61),
.B2(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_86),
.Y(n_117)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_8),
.C(n_9),
.Y(n_124)
);

AO32x1_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_20),
.A3(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_28),
.C(n_48),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_131),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_108),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_31),
.B1(n_45),
.B2(n_44),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_27),
.C(n_43),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_13),
.B(n_17),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_49),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_131),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_144),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_151),
.B(n_125),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_39),
.A3(n_41),
.B1(n_122),
.B2(n_135),
.C1(n_130),
.C2(n_128),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_125),
.C(n_133),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_129),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_126),
.C(n_127),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_142),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_151),
.B(n_145),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_161),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_158),
.B(n_153),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_160),
.CI(n_140),
.CON(n_164),
.SN(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_153),
.B(n_146),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_146),
.B(n_164),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_164),
.C(n_143),
.Y(n_167)
);


endmodule