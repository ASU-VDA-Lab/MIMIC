module fake_jpeg_14856_n_352 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_49),
.B(n_54),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_11),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_58),
.Y(n_82)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_29),
.Y(n_94)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_69),
.Y(n_92)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_27),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_39),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_35),
.B1(n_19),
.B2(n_34),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_78),
.A2(n_106),
.B1(n_115),
.B2(n_1),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_19),
.B1(n_35),
.B2(n_33),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_81),
.A2(n_86),
.B1(n_90),
.B2(n_4),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_19),
.B1(n_35),
.B2(n_33),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_32),
.B(n_33),
.C(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_94),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_16),
.B1(n_39),
.B2(n_31),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_34),
.B1(n_16),
.B2(n_32),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_117),
.B1(n_120),
.B2(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_39),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_107),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_105),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_37),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_20),
.B1(n_37),
.B2(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_30),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_48),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_41),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_114),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_20),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_0),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_61),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_50),
.B(n_30),
.C(n_2),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_118),
.C(n_119),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_131),
.B1(n_139),
.B2(n_142),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_90),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_SL g207 ( 
.A(n_126),
.B(n_134),
.C(n_152),
.Y(n_207)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_74),
.B(n_65),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_140),
.C(n_166),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_79),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_150),
.B1(n_157),
.B2(n_169),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_9),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_76),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_153),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_6),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_156),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_81),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_7),
.B(n_9),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_76),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_158),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_7),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_72),
.B(n_7),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_94),
.A2(n_121),
.B1(n_86),
.B2(n_117),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_113),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_79),
.B1(n_85),
.B2(n_98),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_163),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_92),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_170),
.Y(n_182)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_108),
.A2(n_118),
.B1(n_122),
.B2(n_101),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_116),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_89),
.B(n_102),
.C(n_119),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_170),
.C(n_140),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_82),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_191),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_108),
.B(n_101),
.C(n_116),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_73),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_133),
.A2(n_95),
.B(n_89),
.C(n_87),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_73),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_142),
.A3(n_169),
.B1(n_136),
.B2(n_163),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_135),
.A3(n_124),
.B1(n_141),
.B2(n_153),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_87),
.B1(n_93),
.B2(n_110),
.Y(n_193)
);

AO21x2_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_138),
.B(n_164),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_87),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_128),
.B(n_93),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_137),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_93),
.B1(n_110),
.B2(n_119),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_199),
.B1(n_204),
.B2(n_205),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_110),
.CI(n_156),
.CON(n_198),
.SN(n_198)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_155),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_159),
.B1(n_146),
.B2(n_130),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_130),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_188),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_146),
.A2(n_130),
.B1(n_163),
.B2(n_161),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_150),
.B1(n_155),
.B2(n_140),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.C(n_148),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_167),
.C(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_226),
.C(n_233),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_174),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_207),
.B(n_202),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_219),
.A2(n_220),
.B(n_240),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_193),
.B(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_193),
.B1(n_228),
.B2(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_185),
.A2(n_152),
.B1(n_154),
.B2(n_149),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_232),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_129),
.C(n_144),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_236),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_176),
.A2(n_125),
.B(n_168),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_132),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_132),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_125),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_185),
.A2(n_145),
.B1(n_168),
.B2(n_180),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_192),
.B(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_190),
.C(n_182),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_243),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_254),
.B1(n_267),
.B2(n_268),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_207),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_260),
.B(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_179),
.B1(n_172),
.B2(n_193),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_193),
.B(n_176),
.C(n_180),
.D(n_181),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_214),
.B(n_173),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_265),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_199),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_221),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_224),
.A2(n_172),
.B1(n_184),
.B2(n_209),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_190),
.B1(n_205),
.B2(n_211),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_227),
.C(n_212),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_173),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

AO22x1_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_224),
.B1(n_228),
.B2(n_213),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_280),
.B1(n_293),
.B2(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_238),
.B1(n_236),
.B2(n_213),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_279),
.A2(n_283),
.B1(n_258),
.B2(n_253),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_217),
.B1(n_225),
.B2(n_197),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_241),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_290),
.C(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_243),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_217),
.B1(n_230),
.B2(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_265),
.B(n_225),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_287),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_235),
.B(n_244),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_226),
.B(n_216),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_295),
.Y(n_297)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_232),
.C(n_218),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_215),
.B1(n_237),
.B2(n_187),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_186),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_258),
.C(n_253),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_186),
.B(n_191),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_301),
.A2(n_309),
.B1(n_312),
.B2(n_287),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_306),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_307),
.C(n_311),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_288),
.B(n_279),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_272),
.C(n_260),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_275),
.A2(n_250),
.B1(n_254),
.B2(n_266),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_269),
.C(n_259),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_264),
.B1(n_257),
.B2(n_262),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_285),
.B1(n_293),
.B2(n_273),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_314),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_294),
.C(n_290),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_319),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_278),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_316),
.A2(n_270),
.B(n_299),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_275),
.B(n_274),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_321),
.B(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_284),
.B1(n_292),
.B2(n_289),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_283),
.C(n_277),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_270),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_277),
.C(n_295),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_287),
.C(n_256),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_298),
.A2(n_257),
.B1(n_274),
.B2(n_259),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_297),
.B1(n_304),
.B2(n_306),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_328),
.A2(n_330),
.B(n_324),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_301),
.B(n_300),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_336),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_333),
.A2(n_313),
.B1(n_315),
.B2(n_334),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_317),
.A2(n_305),
.B1(n_308),
.B2(n_297),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_335),
.B1(n_331),
.B2(n_336),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_323),
.A2(n_308),
.B1(n_255),
.B2(n_256),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_255),
.B(n_203),
.C(n_229),
.D(n_222),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_338),
.A2(n_339),
.B(n_340),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_330),
.A2(n_320),
.B(n_322),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_319),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_327),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_327),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_345),
.C(n_346),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_338),
.A2(n_329),
.B(n_335),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

OAI21x1_ASAP7_75t_L g349 ( 
.A1(n_347),
.A2(n_337),
.B(n_340),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_348),
.B(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_350),
.B(n_329),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_313),
.Y(n_352)
);


endmodule