module fake_netlist_1_539_n_688 (n_52, n_50, n_7, n_3, n_34, n_25, n_9, n_72, n_43, n_73, n_62, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_66, n_46, n_37, n_18, n_65, n_5, n_47, n_1, n_16, n_40, n_68, n_36, n_11, n_15, n_71, n_70, n_2, n_17, n_58, n_20, n_12, n_56, n_67, n_22, n_19, n_26, n_39, n_38, n_24, n_35, n_32, n_48, n_63, n_54, n_41, n_55, n_29, n_60, n_10, n_30, n_13, n_75, n_53, n_64, n_69, n_23, n_0, n_57, n_51, n_45, n_42, n_21, n_27, n_28, n_49, n_14, n_31, n_688, n_656);
input n_52;
input n_50;
input n_7;
input n_3;
input n_34;
input n_25;
input n_9;
input n_72;
input n_43;
input n_73;
input n_62;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_66;
input n_46;
input n_37;
input n_18;
input n_65;
input n_5;
input n_47;
input n_1;
input n_16;
input n_40;
input n_68;
input n_36;
input n_11;
input n_15;
input n_71;
input n_70;
input n_2;
input n_17;
input n_58;
input n_20;
input n_12;
input n_56;
input n_67;
input n_22;
input n_19;
input n_26;
input n_39;
input n_38;
input n_24;
input n_35;
input n_32;
input n_48;
input n_63;
input n_54;
input n_41;
input n_55;
input n_29;
input n_60;
input n_10;
input n_30;
input n_13;
input n_75;
input n_53;
input n_64;
input n_69;
input n_23;
input n_0;
input n_57;
input n_51;
input n_45;
input n_42;
input n_21;
input n_27;
input n_28;
input n_49;
input n_14;
input n_31;
output n_688;
output n_656;
wire n_107;
wire n_646;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_169;
wire n_370;
wire n_384;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_357;
wire n_74;
wire n_308;
wire n_518;
wire n_394;
wire n_44;
wire n_189;
wire n_681;
wire n_352;
wire n_226;
wire n_447;
wire n_66;
wire n_379;
wire n_535;
wire n_595;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_475;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_436;
wire n_438;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_223;
wire n_405;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_534;
wire n_569;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_303;
wire n_502;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_246;
wire n_676;
wire n_191;
wire n_143;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_555;
wire n_553;
wire n_135;
wire n_481;
wire n_621;
wire n_315;
wire n_397;
wire n_53;
wire n_213;
wire n_196;
wire n_293;
wire n_127;
wire n_312;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_155;
wire n_162;
wire n_114;
wire n_50;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_636;
wire n_330;
wire n_231;
wire n_9;
wire n_428;
wire n_178;
wire n_478;
wire n_652;
wire n_678;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_441;
wire n_628;
wire n_425;
wire n_314;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_172;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_228;
wire n_671;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_599;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_362;
wire n_617;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_152;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_491;
wire n_388;
wire n_266;
wire n_80;
wire n_632;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_326;
wire n_532;
wire n_635;
wire n_544;
wire n_576;
wire n_275;
wire n_622;
wire n_661;
wire n_493;
wire n_274;
wire n_150;
wire n_235;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_100;
wire n_299;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_193;
wire n_232;
wire n_344;
wire n_147;
wire n_185;
wire n_367;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_212;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_435;
wire n_583;
wire n_64;
wire n_69;
wire n_248;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_119;
wire n_667;
wire n_503;
wire n_339;
wire n_347;
wire n_124;
wire n_79;
wire n_129;
wire n_611;
wire n_521;
wire n_157;
wire n_103;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_325;
wire n_273;
wire n_571;
wire n_524;
wire n_530;
wire n_163;
wire n_348;
wire n_96;
wire n_685;
wire n_669;
wire n_72;
wire n_77;
wire n_90;
wire n_594;
wire n_214;
wire n_167;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_413;
wire n_65;
wire n_537;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_290;
wire n_217;
wire n_201;
wire n_277;
wire n_259;
wire n_612;
wire n_244;
wire n_666;
wire n_297;
wire n_276;
wire n_225;
wire n_631;
wire n_350;
wire n_208;
wire n_616;
wire n_523;
wire n_528;
wire n_419;
wire n_252;
wire n_519;
wire n_168;
wire n_271;
wire n_94;
wire n_194;
wire n_282;
wire n_58;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_116;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_597;
wire n_554;
wire n_257;
wire n_203;
wire n_26;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_146;
wire n_337;
wire n_32;
wire n_637;
wire n_641;
wire n_531;
wire n_93;
wire n_539;
wire n_406;
wire n_372;
wire n_467;
wire n_41;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_647;
wire n_445;
wire n_500;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_75;
wire n_82;
wire n_183;
wire n_550;
wire n_132;
wire n_643;
wire n_582;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_510;
wire n_360;
wire n_363;
wire n_427;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_437;
wire n_620;
wire n_89;
wire n_480;
wire n_130;
wire n_310;
wire n_341;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_136;
wire n_260;
wire n_580;
wire n_610;
wire n_222;
wire n_657;
wire n_381;
wire n_34;
wire n_142;
wire n_385;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_376;
wire n_240;
wire n_459;
wire n_88;
wire n_568;
wire n_46;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_672;
wire n_87;
wire n_466;
wire n_349;
wire n_207;
wire n_197;
wire n_81;
wire n_541;
wire n_572;
wire n_298;
wire n_112;
wire n_630;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_36;
wire n_416;
wire n_432;
wire n_465;
wire n_414;
wire n_680;
wire n_369;
wire n_469;
wire n_361;
wire n_237;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_591;
wire n_391;
wire n_241;
wire n_209;
wire n_20;
wire n_84;
wire n_449;
wire n_56;
wire n_12;
wire n_412;
wire n_455;
wire n_504;
wire n_67;
wire n_618;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_383;
wire n_202;
wire n_319;
wire n_542;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_508;
wire n_486;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_400;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_60;
wire n_138;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_505;
wire n_92;
wire n_313;
wire n_358;
wire n_333;
wire n_627;
wire n_589;
wire n_175;
wire n_128;
wire n_306;
wire n_415;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_234;
wire n_607;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_31;
INVx2_ASAP7_75t_L g77 ( .A(n_60), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_7), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_71), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_72), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_34), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_75), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_39), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_30), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_37), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_27), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_57), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_73), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_52), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_47), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_32), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_76), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_56), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_43), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_66), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_4), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_10), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_63), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_42), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_20), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_11), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_31), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_35), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_7), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_3), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_41), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_45), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_18), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_38), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_18), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_36), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_33), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_15), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_8), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_2), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_5), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_107), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_99), .B(n_0), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_99), .B(n_3), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_80), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_114), .B(n_4), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_77), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_101), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_119), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_119), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_87), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g144 ( .A1(n_78), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_85), .B(n_6), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_122), .B(n_9), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_123), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_77), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_88), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_89), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_91), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_91), .B(n_9), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_94), .B(n_10), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_85), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_113), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_92), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_110), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_93), .B(n_11), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_95), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_103), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_153), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_134), .B(n_112), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_131), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_134), .B(n_112), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_129), .B(n_105), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_142), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_132), .B(n_105), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_126), .B(n_136), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_159), .B(n_115), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_126), .B(n_104), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_128), .A2(n_108), .B1(n_118), .B2(n_93), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_160), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_128), .B(n_115), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
AO22x2_ASAP7_75t_L g191 ( .A1(n_128), .A2(n_103), .B1(n_104), .B2(n_120), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_165), .B(n_116), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_141), .B(n_116), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_139), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_128), .B(n_102), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_145), .B(n_117), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_144), .B(n_102), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_161), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_136), .B(n_120), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_145), .A2(n_121), .B1(n_111), .B2(n_106), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_140), .B(n_106), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_151), .B(n_140), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_150), .B(n_117), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_166), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_133), .B(n_111), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_150), .B(n_121), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_143), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_143), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_143), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_143), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_127), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_127), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_151), .B(n_100), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_151), .B(n_109), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_156), .B(n_97), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_207), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_191), .A2(n_152), .B1(n_158), .B2(n_156), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_207), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_207), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_224), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_202), .Y(n_234) );
BUFx12f_ASAP7_75t_L g235 ( .A(n_199), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_202), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_169), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_172), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_197), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_226), .B(n_158), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_226), .B(n_152), .Y(n_241) );
INVxp67_ASAP7_75t_L g242 ( .A(n_180), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_173), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_176), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_196), .B(n_163), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_197), .B(n_130), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_224), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_226), .B(n_151), .Y(n_250) );
BUFx4f_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_173), .Y(n_252) );
NOR3xp33_ASAP7_75t_SL g253 ( .A(n_192), .B(n_144), .C(n_146), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_196), .B(n_164), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_226), .B(n_157), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_225), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g258 ( .A(n_187), .B(n_124), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_227), .B(n_162), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_182), .Y(n_260) );
AND2x6_ASAP7_75t_SL g261 ( .A(n_198), .B(n_168), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_227), .B(n_162), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_183), .B(n_164), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_175), .B(n_155), .C(n_79), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_206), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_196), .B(n_214), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_216), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_173), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_227), .B(n_162), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_210), .Y(n_271) );
NOR3xp33_ASAP7_75t_SL g272 ( .A(n_177), .B(n_81), .C(n_84), .Y(n_272) );
OR2x4_ASAP7_75t_L g273 ( .A(n_194), .B(n_143), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_189), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_214), .B(n_154), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_210), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_227), .B(n_154), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_191), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_198), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_189), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_184), .Y(n_281) );
AND3x1_ASAP7_75t_SL g282 ( .A(n_198), .B(n_125), .C(n_13), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_210), .Y(n_283) );
AND3x2_ASAP7_75t_SL g284 ( .A(n_191), .B(n_154), .C(n_149), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_183), .B(n_149), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
AOI22xp33_ASAP7_75t_SL g287 ( .A1(n_198), .A2(n_149), .B1(n_125), .B2(n_86), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_191), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_185), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_184), .Y(n_290) );
INVx5_ASAP7_75t_L g291 ( .A(n_205), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_168), .B(n_148), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_174), .Y(n_293) );
INVx6_ASAP7_75t_L g294 ( .A(n_205), .Y(n_294) );
CKINVDCx8_ASAP7_75t_R g295 ( .A(n_238), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_229), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_233), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_278), .Y(n_298) );
BUFx4f_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_231), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_263), .B(n_260), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_237), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_278), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_232), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_233), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_288), .A2(n_198), .B1(n_186), .B2(n_204), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_232), .Y(n_312) );
NOR4xp25_ASAP7_75t_L g313 ( .A(n_230), .B(n_127), .C(n_135), .D(n_148), .Y(n_313) );
OAI21x1_ASAP7_75t_SL g314 ( .A1(n_239), .A2(n_186), .B(n_204), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_289), .A2(n_203), .B(n_208), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_288), .A2(n_174), .B1(n_228), .B2(n_135), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_257), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_257), .Y(n_318) );
AOI21xp33_ASAP7_75t_SL g319 ( .A1(n_279), .A2(n_12), .B(n_13), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_244), .B(n_135), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_SL g321 ( .A1(n_275), .A2(n_217), .B(n_222), .C(n_195), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_248), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
AND2x2_ASAP7_75t_SL g324 ( .A(n_251), .B(n_148), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_263), .B(n_12), .Y(n_326) );
BUFx2_ASAP7_75t_R g327 ( .A(n_279), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_254), .A2(n_205), .B1(n_143), .B2(n_223), .Y(n_329) );
INVx5_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_251), .B(n_205), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_254), .A2(n_98), .B1(n_200), .B2(n_221), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_254), .A2(n_223), .B1(n_220), .B2(n_221), .Y(n_333) );
CKINVDCx11_ASAP7_75t_R g334 ( .A(n_235), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_246), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_260), .B(n_14), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_249), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_258), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_293), .A2(n_220), .B(n_167), .C(n_218), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_249), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_242), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_235), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_289), .A2(n_200), .B1(n_178), .B2(n_179), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_243), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_301), .B(n_247), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_301), .A2(n_256), .B1(n_267), .B2(n_265), .C(n_268), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_319), .B(n_272), .C(n_253), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_314), .A2(n_284), .B1(n_247), .B2(n_282), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_334), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_326), .A2(n_284), .B1(n_277), .B2(n_259), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_296), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_295), .A2(n_293), .B1(n_285), .B2(n_255), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_315), .B(n_299), .Y(n_356) );
NAND2xp33_ASAP7_75t_SL g357 ( .A(n_298), .B(n_284), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_321), .A2(n_250), .B(n_262), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_295), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_341), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_326), .B(n_266), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_299), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_312), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_314), .A2(n_287), .B1(n_274), .B2(n_280), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_325), .A2(n_201), .B(n_222), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_336), .B(n_268), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_304), .B(n_292), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_312), .B(n_234), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
O2A1O1Ixp5_ASAP7_75t_L g373 ( .A1(n_338), .A2(n_195), .B(n_188), .C(n_201), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_217), .B(n_201), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_297), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_306), .A2(n_236), .B1(n_245), .B2(n_240), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_306), .A2(n_241), .B1(n_270), .B2(n_294), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_350), .A2(n_336), .B1(n_339), .B2(n_324), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_366), .B1(n_355), .B2(n_348), .C(n_346), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_346), .B(n_310), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_364), .B(n_330), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_350), .A2(n_310), .B1(n_342), .B2(n_320), .C(n_305), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_347), .A2(n_320), .B1(n_264), .B2(n_316), .C(n_335), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_352), .A2(n_298), .B1(n_324), .B2(n_296), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_298), .B1(n_324), .B2(n_296), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_370), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_370), .Y(n_387) );
AND2x4_ASAP7_75t_SL g388 ( .A(n_364), .B(n_307), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_374), .A2(n_344), .B(n_345), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_298), .B1(n_300), .B2(n_302), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_361), .A2(n_335), .B1(n_343), .B2(n_307), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_348), .A2(n_316), .B1(n_343), .B2(n_313), .C(n_332), .Y(n_392) );
AND2x4_ASAP7_75t_SL g393 ( .A(n_356), .B(n_307), .Y(n_393) );
CKINVDCx8_ASAP7_75t_R g394 ( .A(n_360), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_368), .B(n_296), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_363), .A2(n_296), .B1(n_308), .B2(n_302), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_365), .A2(n_302), .B1(n_308), .B2(n_300), .Y(n_397) );
AND2x4_ASAP7_75t_SL g398 ( .A(n_356), .B(n_307), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_360), .B(n_330), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_372), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_357), .A2(n_309), .B1(n_311), .B2(n_303), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_368), .B(n_261), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_358), .B(n_319), .C(n_313), .Y(n_405) );
NOR4xp25_ASAP7_75t_SL g406 ( .A(n_382), .B(n_365), .C(n_353), .D(n_362), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_379), .A2(n_376), .B1(n_369), .B2(n_377), .C(n_332), .Y(n_407) );
OR2x6_ASAP7_75t_SL g408 ( .A(n_384), .B(n_327), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_387), .B(n_369), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_405), .A2(n_374), .B(n_358), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_395), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_380), .B(n_349), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_405), .B(n_378), .C(n_392), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_387), .B(n_349), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_353), .B(n_362), .C(n_359), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_400), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_400), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_404), .B(n_359), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_404), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_385), .A2(n_367), .B(n_374), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
BUFx10_ASAP7_75t_L g422 ( .A(n_399), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_383), .A2(n_329), .B1(n_333), .B2(n_317), .C(n_311), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_394), .A2(n_351), .B(n_330), .C(n_331), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_393), .A2(n_371), .B1(n_330), .B2(n_308), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_393), .B(n_375), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g429 ( .A1(n_402), .A2(n_211), .A3(n_178), .B1(n_179), .B2(n_181), .B3(n_193), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_403), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_398), .B(n_375), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_398), .A2(n_371), .B1(n_308), .B2(n_302), .Y(n_432) );
NOR4xp25_ASAP7_75t_L g433 ( .A(n_401), .B(n_375), .C(n_354), .D(n_317), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_390), .A2(n_371), .B1(n_303), .B2(n_309), .C(n_323), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g438 ( .A1(n_388), .A2(n_371), .A3(n_309), .B(n_297), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
NAND4xp75_ASAP7_75t_L g440 ( .A(n_381), .B(n_367), .C(n_373), .D(n_273), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_409), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_421), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_416), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_416), .B(n_403), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_419), .B(n_403), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_354), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_421), .Y(n_448) );
NAND4xp25_ASAP7_75t_SL g449 ( .A(n_426), .B(n_14), .C(n_16), .D(n_17), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_408), .Y(n_450) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_438), .B(n_397), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_421), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_419), .B(n_354), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_423), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_409), .B(n_381), .Y(n_456) );
AND4x1_ASAP7_75t_L g457 ( .A(n_438), .B(n_16), .C(n_17), .D(n_19), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_422), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_417), .B(n_396), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_411), .B(n_388), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_417), .B(n_367), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_436), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_407), .B(n_330), .Y(n_463) );
NOR2x1p5_ASAP7_75t_L g464 ( .A(n_441), .B(n_300), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_426), .B(n_373), .C(n_218), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_415), .B(n_330), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_420), .A2(n_367), .B(n_300), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_415), .B(n_302), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_407), .A2(n_308), .B1(n_300), .B2(n_328), .Y(n_474) );
OAI321xp33_ASAP7_75t_L g475 ( .A1(n_413), .A2(n_211), .A3(n_181), .B1(n_193), .B2(n_167), .C(n_212), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_412), .B(n_19), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_418), .B(n_345), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_418), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_430), .B(n_431), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_413), .A2(n_429), .B1(n_437), .B2(n_435), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_430), .B(n_188), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_412), .B(n_273), .Y(n_482) );
AOI33xp33_ASAP7_75t_L g483 ( .A1(n_406), .A2(n_212), .A3(n_213), .B1(n_222), .B2(n_171), .B3(n_195), .Y(n_483) );
INVx4_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_428), .B(n_337), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_337), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_427), .A2(n_328), .B1(n_323), .B2(n_337), .C(n_318), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_435), .B(n_337), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_439), .Y(n_491) );
OAI31xp33_ASAP7_75t_SL g492 ( .A1(n_408), .A2(n_273), .A3(n_318), .B(n_24), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_450), .B(n_441), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_454), .B(n_410), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_442), .B(n_435), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_478), .B(n_441), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_479), .B(n_422), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_450), .B(n_441), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_472), .B(n_428), .Y(n_499) );
HB1xp67_ASAP7_75t_SL g500 ( .A(n_484), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_467), .B(n_434), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_455), .B(n_410), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_467), .B(n_433), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_455), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_443), .B(n_410), .Y(n_505) );
NAND4xp25_ASAP7_75t_L g506 ( .A(n_463), .B(n_437), .C(n_432), .D(n_420), .Y(n_506) );
NOR4xp25_ASAP7_75t_SL g507 ( .A(n_466), .B(n_406), .C(n_425), .D(n_433), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_443), .B(n_410), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_470), .B(n_440), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_448), .B(n_422), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_470), .B(n_477), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_449), .B(n_425), .C(n_440), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_477), .B(n_337), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_476), .B(n_171), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_448), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_444), .B(n_171), .Y(n_517) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_484), .B(n_217), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_476), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_452), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_479), .B(n_188), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_456), .B(n_485), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_461), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_461), .B(n_219), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_459), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_445), .B(n_215), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_458), .Y(n_528) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_484), .B(n_170), .Y(n_529) );
NOR2xp33_ASAP7_75t_R g530 ( .A(n_484), .B(n_451), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_462), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_482), .B(n_219), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g533 ( .A1(n_460), .A2(n_213), .A3(n_215), .B1(n_190), .B2(n_170), .B3(n_29), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_485), .B(n_190), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_445), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_462), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_462), .Y(n_537) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_464), .B(n_323), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_446), .B(n_219), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_447), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_446), .B(n_219), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_446), .B(n_219), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_483), .B(n_184), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_447), .Y(n_545) );
OAI211xp5_ASAP7_75t_SL g546 ( .A1(n_492), .A2(n_220), .B(n_328), .C(n_276), .Y(n_546) );
NOR4xp25_ASAP7_75t_SL g547 ( .A(n_471), .B(n_21), .C(n_22), .D(n_26), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_446), .B(n_28), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_453), .B(n_219), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_535), .B(n_497), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_519), .A2(n_480), .B1(n_474), .B2(n_451), .C(n_487), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_525), .B(n_453), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_500), .A2(n_464), .B1(n_488), .B2(n_490), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_522), .B(n_487), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_512), .A2(n_488), .B1(n_490), .B2(n_481), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_493), .A2(n_481), .B1(n_489), .B2(n_457), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_504), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_515), .Y(n_559) );
AOI21xp33_ASAP7_75t_L g560 ( .A1(n_503), .A2(n_481), .B(n_486), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_528), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_526), .B(n_486), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_523), .B(n_457), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_540), .B(n_468), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_507), .B(n_481), .C(n_465), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_516), .Y(n_566) );
AND2x4_ASAP7_75t_SL g567 ( .A(n_510), .B(n_468), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_506), .A2(n_469), .B1(n_468), .B2(n_473), .Y(n_568) );
O2A1O1Ixp5_ASAP7_75t_L g569 ( .A1(n_538), .A2(n_468), .B(n_491), .C(n_220), .Y(n_569) );
NAND2xp33_ASAP7_75t_L g570 ( .A(n_530), .B(n_491), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_545), .B(n_491), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_511), .B(n_209), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_493), .A2(n_475), .B1(n_291), .B2(n_209), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_498), .A2(n_184), .B1(n_209), .B2(n_276), .C(n_269), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_510), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_520), .Y(n_577) );
OAI31xp33_ASAP7_75t_SL g578 ( .A1(n_498), .A2(n_40), .A3(n_44), .B(n_46), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_48), .Y(n_579) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_531), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_529), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_501), .Y(n_582) );
AOI22xp5_ASAP7_75t_SL g583 ( .A1(n_530), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_494), .B(n_184), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_518), .A2(n_291), .B(n_271), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g586 ( .A1(n_496), .A2(n_184), .A3(n_209), .B1(n_59), .B2(n_61), .C1(n_62), .C2(n_64), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_509), .A2(n_291), .B1(n_209), .B2(n_294), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_495), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_209), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_538), .A2(n_53), .B(n_55), .C(n_65), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_544), .A2(n_291), .B(n_269), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_494), .B(n_67), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_527), .B(n_68), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_502), .B(n_69), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_549), .A2(n_281), .B1(n_290), .B2(n_70), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_502), .B(n_281), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_505), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_524), .B(n_243), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_508), .B(n_271), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_549), .A2(n_281), .B1(n_290), .B2(n_283), .Y(n_601) );
XNOR2xp5_ASAP7_75t_L g602 ( .A(n_561), .B(n_521), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_556), .B(n_578), .C(n_565), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_597), .B(n_508), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_558), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_570), .A2(n_546), .B(n_544), .C(n_549), .Y(n_606) );
INVxp33_ASAP7_75t_L g607 ( .A(n_583), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_582), .B(n_531), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_574), .B(n_536), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_588), .B(n_548), .Y(n_610) );
NOR4xp25_ASAP7_75t_SL g611 ( .A(n_552), .B(n_533), .C(n_547), .D(n_517), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_559), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_598), .B(n_536), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_570), .A2(n_532), .B(n_514), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_566), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_576), .A2(n_542), .B(n_541), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_577), .Y(n_617) );
NAND2xp33_ASAP7_75t_SL g618 ( .A(n_554), .B(n_537), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_581), .B(n_542), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_563), .A2(n_541), .B1(n_550), .B2(n_537), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_553), .B(n_548), .Y(n_622) );
AOI211xp5_ASAP7_75t_SL g623 ( .A1(n_568), .A2(n_534), .B(n_539), .C(n_550), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_562), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_551), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_571), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_580), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_580), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_560), .A2(n_543), .B(n_281), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_564), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_557), .B(n_281), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_572), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_567), .B(n_283), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_552), .B(n_290), .Y(n_635) );
AOI221x1_ASAP7_75t_L g636 ( .A1(n_618), .A2(n_591), .B1(n_592), .B2(n_594), .C(n_590), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_607), .B(n_568), .Y(n_637) );
XNOR2x1_ASAP7_75t_L g638 ( .A(n_602), .B(n_579), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_608), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_603), .B(n_575), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_624), .A2(n_587), .B1(n_573), .B2(n_595), .C(n_600), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_630), .B(n_596), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_621), .B(n_589), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_625), .B(n_593), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g645 ( .A(n_631), .B(n_569), .C(n_585), .D(n_587), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_627), .Y(n_646) );
XNOR2xp5_ASAP7_75t_L g647 ( .A(n_620), .B(n_599), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_616), .A2(n_590), .B(n_601), .C(n_569), .Y(n_648) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_628), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_605), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_623), .A2(n_586), .B(n_290), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_626), .B(n_290), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_632), .B(n_252), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_619), .A2(n_252), .B1(n_286), .B2(n_606), .Y(n_654) );
O2A1O1Ixp5_ASAP7_75t_L g655 ( .A1(n_623), .A2(n_286), .B(n_610), .C(n_615), .Y(n_655) );
UNKNOWN g656 ( );
INVx1_ASAP7_75t_L g657 ( .A(n_612), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_638), .B(n_617), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_646), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_637), .B(n_604), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_639), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_649), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_649), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_637), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_647), .Y(n_665) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_645), .B(n_633), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_650), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_640), .B(n_629), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_640), .A2(n_634), .B1(n_635), .B2(n_619), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_643), .A2(n_644), .B1(n_656), .B2(n_642), .Y(n_670) );
AND4x1_ASAP7_75t_L g671 ( .A(n_655), .B(n_611), .C(n_604), .D(n_613), .Y(n_671) );
NAND2x1_ASAP7_75t_SL g672 ( .A(n_643), .B(n_613), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_657), .Y(n_673) );
AND4x1_ASAP7_75t_L g674 ( .A(n_636), .B(n_609), .C(n_622), .D(n_648), .Y(n_674) );
NAND4xp25_ASAP7_75t_SL g675 ( .A(n_651), .B(n_641), .C(n_653), .D(n_652), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_654), .A2(n_637), .B1(n_640), .B2(n_603), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_664), .B(n_676), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_659), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_675), .B(n_666), .C(n_668), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_662), .Y(n_680) );
NOR3xp33_ASAP7_75t_SL g681 ( .A(n_677), .B(n_658), .C(n_660), .Y(n_681) );
NOR4xp75_ASAP7_75t_L g682 ( .A(n_679), .B(n_672), .C(n_674), .D(n_671), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_678), .B(n_665), .Y(n_683) );
OAI21x1_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_680), .B(n_663), .Y(n_684) );
XNOR2xp5_ASAP7_75t_L g685 ( .A(n_682), .B(n_665), .Y(n_685) );
AOI22x1_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_662), .B1(n_681), .B2(n_673), .Y(n_686) );
AOI322xp5_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_684), .A3(n_663), .B1(n_669), .B2(n_670), .C1(n_661), .C2(n_667), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_687), .Y(n_688) );
endmodule