module fake_netlist_6_4391_n_488 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_488);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_488;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_466;
wire n_360;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_153;
wire n_156;
wire n_145;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_6),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_46),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_53),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_62),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_122),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVxp33_ASAP7_75t_SL g158 ( 
.A(n_109),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_33),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVxp33_ASAP7_75t_SL g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_48),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_3),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_25),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_0),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_30),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_24),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_64),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_37),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_50),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_3),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_137),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_28),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_92),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_76),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_102),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_82),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_69),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_18),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_16),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_85),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_26),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_52),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_84),
.Y(n_218)
);

INVxp33_ASAP7_75t_SL g219 ( 
.A(n_36),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_21),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_63),
.Y(n_223)
);

INVxp33_ASAP7_75t_SL g224 ( 
.A(n_19),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_51),
.Y(n_225)
);

INVxp33_ASAP7_75t_SL g226 ( 
.A(n_86),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_1),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_190),
.B(n_2),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_2),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_155),
.B(n_4),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_203),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_155),
.B(n_5),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_153),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_175),
.B(n_6),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_151),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_160),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_145),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_7),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_152),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_165),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_216),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_193),
.B(n_7),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_175),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_157),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_145),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_143),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_238),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_143),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_161),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_161),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_206),
.Y(n_286)
);

OAI22x1_ASAP7_75t_L g287 ( 
.A1(n_231),
.A2(n_206),
.B1(n_169),
.B2(n_225),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_188),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_8),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_251),
.B(n_188),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_262),
.A2(n_214),
.B1(n_146),
.B2(n_226),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_228),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_214),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_218),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_231),
.A2(n_158),
.B1(n_163),
.B2(n_185),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_221),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_251),
.B(n_202),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_253),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

OR2x6_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_236),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_261),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_149),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_283),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_154),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_156),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_303),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

NAND2xp33_ASAP7_75t_SL g323 ( 
.A(n_287),
.B(n_159),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_SL g324 ( 
.A(n_295),
.B(n_234),
.C(n_201),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_291),
.Y(n_326)
);

O2A1O1Ixp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_232),
.B(n_229),
.C(n_174),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_303),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_219),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_300),
.B(n_194),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_SL g332 ( 
.A(n_295),
.B(n_200),
.C(n_173),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_284),
.Y(n_336)
);

OR2x2_ASAP7_75t_SL g337 ( 
.A(n_292),
.B(n_196),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_170),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_178),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_278),
.B(n_232),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_179),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_314),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_331),
.A2(n_304),
.B1(n_286),
.B2(n_276),
.Y(n_351)
);

BUFx4f_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_276),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_347),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_347),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_310),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_334),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_313),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_328),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_233),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_346),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_329),
.A2(n_286),
.B1(n_224),
.B2(n_181),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_338),
.A2(n_301),
.B(n_299),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_271),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_274),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_326),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_301),
.Y(n_373)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_330),
.B(n_223),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_280),
.B(n_222),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

BUFx12f_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_337),
.A2(n_220),
.B1(n_215),
.B2(n_213),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_182),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_183),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_331),
.A2(n_211),
.B1(n_210),
.B2(n_209),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_320),
.B(n_184),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_341),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_311),
.A2(n_208),
.B(n_207),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_324),
.Y(n_389)
);

AOI222xp33_ASAP7_75t_L g390 ( 
.A1(n_364),
.A2(n_366),
.B1(n_381),
.B2(n_363),
.C1(n_358),
.C2(n_389),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_349),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_387),
.Y(n_393)
);

OR2x6_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_345),
.Y(n_394)
);

AOI221xp5_ASAP7_75t_SL g395 ( 
.A1(n_384),
.A2(n_366),
.B1(n_351),
.B2(n_373),
.C(n_367),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_373),
.A2(n_324),
.B1(n_332),
.B2(n_349),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_353),
.A2(n_323),
.B1(n_309),
.B2(n_308),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_323),
.B1(n_309),
.B2(n_308),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_322),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_332),
.B1(n_186),
.B2(n_205),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_356),
.A2(n_322),
.B1(n_325),
.B2(n_187),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_357),
.A2(n_327),
.B(n_319),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_325),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_382),
.A2(n_189),
.B1(n_192),
.B2(n_199),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_372),
.A2(n_204),
.B1(n_319),
.B2(n_317),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_327),
.B(n_315),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_318),
.Y(n_408)
);

OAI211xp5_ASAP7_75t_SL g409 ( 
.A1(n_361),
.A2(n_318),
.B(n_9),
.C(n_8),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_359),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_312),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_312),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_374),
.A2(n_317),
.B1(n_315),
.B2(n_12),
.Y(n_415)
);

NOR3xp33_ASAP7_75t_SL g416 ( 
.A(n_381),
.B(n_9),
.C(n_10),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_350),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_315),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_395),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

OAI21xp33_ASAP7_75t_SL g421 ( 
.A1(n_397),
.A2(n_368),
.B(n_386),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_396),
.B(n_407),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_412),
.Y(n_423)
);

OAI211xp5_ASAP7_75t_L g424 ( 
.A1(n_390),
.A2(n_375),
.B(n_376),
.C(n_352),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_399),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_354),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_414),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_405),
.A2(n_371),
.B1(n_369),
.B2(n_352),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_355),
.B1(n_354),
.B2(n_371),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_392),
.A2(n_355),
.B1(n_354),
.B2(n_388),
.Y(n_430)
);

OAI221xp5_ASAP7_75t_L g431 ( 
.A1(n_404),
.A2(n_400),
.B1(n_401),
.B2(n_406),
.C(n_416),
.Y(n_431)
);

BUFx12f_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

OAI22xp33_ASAP7_75t_L g434 ( 
.A1(n_415),
.A2(n_142),
.B1(n_14),
.B2(n_17),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_393),
.A2(n_13),
.B1(n_20),
.B2(n_23),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_408),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_392),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_431),
.A2(n_398),
.B(n_409),
.C(n_411),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_418),
.C(n_412),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_141),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_38),
.B(n_39),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_433),
.Y(n_442)
);

BUFx12f_ASAP7_75t_L g443 ( 
.A(n_432),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_41),
.Y(n_444)
);

OAI211xp5_ASAP7_75t_SL g445 ( 
.A1(n_427),
.A2(n_140),
.B(n_43),
.C(n_44),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_42),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g448 ( 
.A1(n_421),
.A2(n_45),
.B(n_47),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_434),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_57),
.Y(n_450)
);

OAI221xp5_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.C(n_65),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_437),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_446),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_426),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_435),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_439),
.B(n_429),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_430),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_444),
.Y(n_459)
);

AOI33xp33_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_66),
.A3(n_67),
.B1(n_70),
.B2(n_71),
.B3(n_72),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_74),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_444),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_133),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_88),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_90),
.C(n_91),
.Y(n_465)
);

OAI31xp33_ASAP7_75t_SL g466 ( 
.A1(n_463),
.A2(n_445),
.A3(n_451),
.B(n_448),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_455),
.A2(n_443),
.B(n_94),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_93),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_97),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_458),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_98),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_460),
.B(n_100),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_462),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_456),
.Y(n_476)
);

AOI221x1_ASAP7_75t_L g477 ( 
.A1(n_473),
.A2(n_465),
.B1(n_464),
.B2(n_460),
.C(n_461),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_474),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_SL g479 ( 
.A1(n_478),
.A2(n_466),
.B(n_476),
.Y(n_479)
);

OAI211xp5_ASAP7_75t_L g480 ( 
.A1(n_479),
.A2(n_477),
.B(n_467),
.C(n_472),
.Y(n_480)
);

AOI211xp5_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_472),
.B(n_470),
.C(n_468),
.Y(n_481)
);

NAND4xp25_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_105),
.C(n_107),
.D(n_108),
.Y(n_482)
);

NAND4xp25_ASAP7_75t_L g483 ( 
.A(n_482),
.B(n_111),
.C(n_114),
.D(n_115),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_483),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_483),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_484),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_485),
.B1(n_119),
.B2(n_121),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_130),
.B(n_132),
.Y(n_488)
);


endmodule