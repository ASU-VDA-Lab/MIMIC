module fake_jpeg_2741_n_251 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_1),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_54),
.B(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_62),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_20),
.B(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_26),
.B1(n_28),
.B2(n_19),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_81),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_32),
.B1(n_21),
.B2(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_80),
.B1(n_83),
.B2(n_2),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_21),
.B1(n_29),
.B2(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_34),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_21),
.B1(n_29),
.B2(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_18),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_98),
.C(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_97),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_27),
.B1(n_35),
.B2(n_30),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_85),
.B1(n_101),
.B2(n_84),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_27),
.Y(n_98)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_67),
.A3(n_41),
.B1(n_30),
.B2(n_36),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_40),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_110),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_26),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_120),
.C(n_121),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_123),
.B1(n_130),
.B2(n_132),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_122),
.B1(n_84),
.B2(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_2),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_28),
.C(n_19),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_70),
.A2(n_28),
.B1(n_3),
.B2(n_6),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_126),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_7),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_131),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_89),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_11),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_74),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_148),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_82),
.B1(n_75),
.B2(n_101),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_144),
.B1(n_145),
.B2(n_108),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_89),
.B(n_100),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_150),
.B(n_13),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_82),
.B1(n_74),
.B2(n_96),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_96),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_112),
.B(n_120),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_113),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_11),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_99),
.B1(n_8),
.B2(n_13),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_125),
.B1(n_112),
.B2(n_111),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_99),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_135),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_107),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_124),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_180),
.B1(n_155),
.B2(n_139),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_108),
.B1(n_102),
.B2(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_129),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_172),
.B(n_176),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_132),
.Y(n_173)
);

BUFx4f_ASAP7_75t_SL g193 ( 
.A(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_122),
.B1(n_8),
.B2(n_99),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_15),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_15),
.B1(n_144),
.B2(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_197),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_134),
.C(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_160),
.C(n_161),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_136),
.B(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_189),
.A2(n_173),
.B(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_196),
.B1(n_157),
.B2(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_135),
.B1(n_151),
.B2(n_157),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_161),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_199),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_181),
.B(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_165),
.C(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_209),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_180),
.B(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_212),
.A2(n_213),
.B1(n_185),
.B2(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_187),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_218),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_183),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_204),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_186),
.B(n_206),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_230),
.B(n_192),
.C(n_217),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_186),
.B(n_202),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_207),
.Y(n_231)
);

XOR2x1_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_221),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_228),
.B(n_182),
.C(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_231),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_226),
.B(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_226),
.C(n_227),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_235),
.A2(n_207),
.B1(n_211),
.B2(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_190),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_235),
.B(n_234),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_197),
.C(n_193),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_238),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_247),
.B(n_244),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_193),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_193),
.Y(n_251)
);


endmodule