module real_jpeg_22118_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_331, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_331;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_33),
.B1(n_43),
.B2(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_0),
.A2(n_33),
.B1(n_60),
.B2(n_61),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_1),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_48),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_2),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_14),
.B(n_61),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_43),
.B1(n_46),
.B2(n_128),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_103),
.B1(n_185),
.B2(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_85),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_30),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_2),
.A2(n_30),
.B(n_213),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_3),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_125),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_43),
.B1(n_46),
.B2(n_125),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_125),
.Y(n_263)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_5),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_123),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_123),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_5),
.A2(n_43),
.B1(n_46),
.B2(n_123),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_43),
.B1(n_46),
.B2(n_55),
.Y(n_112)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_137),
.B(n_159),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_8),
.A2(n_35),
.B1(n_43),
.B2(n_46),
.Y(n_255)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_11),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_11),
.A2(n_43),
.B1(n_46),
.B2(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_130),
.Y(n_185)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_14),
.A2(n_43),
.B(n_58),
.C(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_43),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_92),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_90),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_76),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_68),
.C(n_71),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_20),
.A2(n_21),
.B1(n_68),
.B2(n_317),
.Y(n_323)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_38),
.B2(n_67),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_23),
.A2(n_36),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_23),
.A2(n_36),
.B1(n_143),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_23),
.A2(n_263),
.B(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_23),
.A2(n_82),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_24),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_24),
.A2(n_28),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_25),
.B(n_30),
.Y(n_134)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g127 ( 
.A(n_26),
.B(n_128),
.CON(n_127),
.SN(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_29),
.B1(n_127),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_28),
.B(n_283),
.Y(n_282)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_29),
.A2(n_43),
.A3(n_45),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_42),
.B(n_44),
.C(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_31),
.A2(n_36),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_36),
.B(n_128),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_49),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_41),
.A2(n_50),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_42),
.A2(n_51),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_42),
.A2(n_51),
.B1(n_122),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_42),
.A2(n_51),
.B1(n_155),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_42),
.A2(n_49),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_42),
.A2(n_51),
.B1(n_74),
.B2(n_279),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_44),
.B(n_46),
.Y(n_214)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_46),
.A2(n_62),
.B(n_128),
.C(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_73),
.B(n_75),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_50),
.A2(n_75),
.B(n_86),
.Y(n_265)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_66),
.C(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_56),
.A2(n_65),
.B1(n_72),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_59),
.B(n_63),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_63),
.B(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_57),
.A2(n_59),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_57),
.A2(n_59),
.B1(n_181),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_57),
.A2(n_59),
.B1(n_202),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_57),
.A2(n_220),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_57),
.A2(n_59),
.B1(n_110),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_57),
.A2(n_118),
.B(n_255),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_59),
.B(n_128),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_60),
.B(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_64),
.B(n_119),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.C(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_68),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_68),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_71),
.B(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_72),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_314),
.A3(n_324),
.B1(n_327),
.B2(n_328),
.C(n_331),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_294),
.B(n_313),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_270),
.B(n_293),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_160),
.B(n_245),
.C(n_269),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_148),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_97),
.B(n_148),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_131),
.B2(n_147),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_115),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_100),
.B(n_115),
.C(n_147),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_109),
.B2(n_114),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_101),
.B(n_114),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_105),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_103),
.A2(n_138),
.B1(n_170),
.B2(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_103),
.A2(n_173),
.B(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_103),
.A2(n_104),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_107),
.A2(n_168),
.B(n_205),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_111),
.B(n_236),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_126),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_138),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_132),
.B(n_140),
.C(n_145),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_149),
.B(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_154),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_159),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_244),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_238),
.B(n_243),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_225),
.B(n_237),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_207),
.B(n_224),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_194),
.B(n_206),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_182),
.B(n_193),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_178),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_187),
.B(n_192),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_195),
.B(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_205),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_215),
.B1(n_222),
.B2(n_223),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_227),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_234),
.C(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_267),
.B2(n_268),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_257),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_257),
.C(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_266),
.Y(n_257)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_272),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_292),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_285),
.B2(n_286),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_286),
.C(n_292),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_280),
.C(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_280),
.B1(n_281),
.B2(n_284),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_288),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_304),
.B(n_308),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_290),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_295),
.B(n_296),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_311),
.B2(n_312),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_303),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_303),
.C(n_312),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_301),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_316),
.C(n_321),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_302),
.B(n_316),
.CI(n_321),
.CON(n_326),
.SN(n_326)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_308),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_322),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_326),
.Y(n_329)
);


endmodule