module real_jpeg_28918_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_58),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_0),
.A2(n_33),
.B1(n_37),
.B2(n_58),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_77),
.B1(n_78),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_1),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_104),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_104),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_1),
.A2(n_33),
.B1(n_37),
.B2(n_104),
.Y(n_223)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_2),
.A2(n_90),
.B(n_164),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_77),
.B1(n_78),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_4),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_149),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_149),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_29),
.B1(n_77),
.B2(n_78),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_6),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_124)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_11),
.B(n_33),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_56),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_33),
.B1(n_37),
.B2(n_56),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_10),
.A2(n_44),
.B1(n_77),
.B2(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_10),
.A2(n_33),
.B1(n_37),
.B2(n_44),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_11),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_48),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_48),
.B(n_188),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_147),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_11),
.B(n_97),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_236),
.Y(n_238)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_15),
.A2(n_77),
.B1(n_78),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_15),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_129),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_129),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_15),
.A2(n_33),
.B1(n_37),
.B2(n_129),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_107),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_106),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_45),
.B(n_59),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_25),
.A2(n_41),
.B(n_196),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_26),
.Y(n_140)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_30),
.B1(n_36),
.B2(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_27),
.B(n_52),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_27),
.A2(n_36),
.B(n_147),
.C(n_215),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_30),
.A2(n_49),
.A3(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_31),
.B(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_32),
.A2(n_41),
.B1(n_69),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_32),
.A2(n_39),
.B(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_32),
.A2(n_41),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_32),
.A2(n_41),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_32),
.A2(n_41),
.B1(n_195),
.B2(n_213),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_32),
.B(n_147),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_64),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_37),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_41),
.A2(n_70),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_46),
.A2(n_51),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_46),
.A2(n_51),
.B1(n_143),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_46),
.A2(n_51),
.B1(n_173),
.B2(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_49),
.B1(n_75),
.B2(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_48),
.B(n_75),
.Y(n_161)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_49),
.A2(n_79),
.B1(n_146),
.B2(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_51),
.B(n_124),
.Y(n_158)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_72),
.B1(n_73),
.B2(n_85),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_68),
.B1(n_85),
.B2(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_63),
.A2(n_64),
.B1(n_117),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_63),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_92),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_63),
.A2(n_65),
.B1(n_228),
.B2(n_236),
.Y(n_235)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_64),
.B(n_147),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_67),
.A2(n_119),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_81),
.B(n_82),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_80),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B(n_79),
.C(n_80),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_77),
.Y(n_79)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g146 ( 
.A(n_77),
.B(n_147),
.CON(n_146),
.SN(n_146)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_102),
.B1(n_103),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_83),
.A2(n_102),
.B1(n_128),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_83),
.B(n_147),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.C(n_100),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_94),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_88),
.B(n_94),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_93),
.A2(n_185),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_105),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_114),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_112),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_114),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.C(n_126),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_115),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_121),
.A2(n_126),
.B1(n_127),
.B2(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_121),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B(n_125),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_273),
.B(n_278),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_177),
.B(n_259),
.C(n_272),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_165),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_134),
.B(n_165),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_150),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_136),
.B(n_137),
.C(n_150),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_145),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_148),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_159),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_152),
.B(n_156),
.C(n_159),
.Y(n_270)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_166),
.A2(n_167),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_171),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_175),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_172),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_201),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_258),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_251),
.B(n_257),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_206),
.B(n_250),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_197),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_181),
.B(n_197),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.C(n_193),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_182),
.A2(n_183),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_186),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_204),
.C(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_244),
.B(n_249),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_224),
.B(n_243),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_223),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_242),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_230),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_241),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_270),
.B2(n_271),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_267),
.C(n_271),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);


endmodule