module fake_jpeg_20703_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_17),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_19),
.B1(n_31),
.B2(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_51),
.B1(n_76),
.B2(n_40),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_19),
.B1(n_31),
.B2(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_56),
.B(n_34),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_69),
.Y(n_87)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_27),
.Y(n_105)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_19),
.B1(n_31),
.B2(n_33),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_73),
.B1(n_34),
.B2(n_35),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_20),
.B1(n_19),
.B2(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_47),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_84),
.B1(n_32),
.B2(n_24),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_85),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_97),
.B1(n_106),
.B2(n_108),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_28),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_92),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_52),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_46),
.C(n_43),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_98),
.C(n_39),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_45),
.B1(n_46),
.B2(n_43),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_107),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_43),
.B1(n_39),
.B2(n_30),
.Y(n_106)
);

INVx2_ASAP7_75t_R g107 ( 
.A(n_53),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_39),
.B1(n_35),
.B2(n_33),
.Y(n_108)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_53),
.A2(n_26),
.B1(n_35),
.B2(n_33),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_18),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_32),
.B1(n_18),
.B2(n_34),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_67),
.B1(n_77),
.B2(n_59),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_135),
.B1(n_81),
.B2(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_70),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_24),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_144),
.C(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_32),
.B1(n_60),
.B2(n_62),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_108),
.B(n_24),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_28),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_120),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_28),
.B1(n_22),
.B2(n_24),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_142),
.B1(n_127),
.B2(n_128),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_143),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_27),
.C(n_28),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_150),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_85),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_97),
.C(n_106),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_178),
.C(n_22),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_161),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_108),
.B(n_94),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_159),
.B(n_172),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_156),
.A2(n_164),
.B1(n_172),
.B2(n_151),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_13),
.C(n_12),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_13),
.B(n_12),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_163),
.B1(n_171),
.B2(n_173),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_113),
.B(n_81),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_111),
.B1(n_109),
.B2(n_89),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_24),
.B(n_28),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_180),
.B(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_162),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_122),
.B1(n_27),
.B2(n_2),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_118),
.A2(n_111),
.B1(n_109),
.B2(n_89),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_146),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_102),
.B1(n_100),
.B2(n_96),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_83),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_16),
.Y(n_175)
);

OAI221xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_110),
.B1(n_16),
.B2(n_22),
.C(n_100),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_R g193 ( 
.A1(n_176),
.A2(n_22),
.B1(n_27),
.B2(n_16),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_22),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_22),
.B(n_27),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_192),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_190),
.B(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_138),
.B1(n_125),
.B2(n_147),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_202),
.B1(n_206),
.B2(n_210),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_133),
.A3(n_128),
.B1(n_127),
.B2(n_140),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_176),
.B(n_177),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_121),
.B1(n_13),
.B2(n_11),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_196),
.B1(n_3),
.B2(n_4),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_195),
.B(n_207),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_22),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_27),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_149),
.A2(n_122),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_122),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_122),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_148),
.C(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_171),
.B1(n_160),
.B2(n_165),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_189),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_152),
.C(n_172),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_228),
.C(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_233),
.B1(n_234),
.B2(n_237),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_222),
.Y(n_251)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_156),
.A3(n_155),
.B1(n_161),
.B2(n_175),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_154),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_180),
.C(n_155),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_231),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_181),
.B1(n_154),
.B2(n_10),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_238),
.B1(n_210),
.B2(n_206),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_194),
.B1(n_184),
.B2(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_208),
.C(n_207),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_244),
.C(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_189),
.C(n_188),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_188),
.C(n_186),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_254),
.C(n_257),
.Y(n_269)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_228),
.A2(n_209),
.B1(n_192),
.B2(n_182),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_217),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_198),
.C(n_196),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_8),
.C(n_218),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_229),
.B1(n_215),
.B2(n_222),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_239),
.B(n_227),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_216),
.B(n_239),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_244),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_274),
.B1(n_277),
.B2(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_276),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_229),
.B(n_217),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_266),
.B(n_277),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_233),
.B1(n_234),
.B2(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_238),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_8),
.B1(n_250),
.B2(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_275),
.Y(n_290)
);

NOR2x1_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_257),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_273),
.B(n_264),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_281),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_240),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_276),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_289),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_241),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_287),
.C(n_269),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_290),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_254),
.C(n_246),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_279),
.B1(n_266),
.B2(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_293),
.C(n_285),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_298),
.B1(n_296),
.B2(n_294),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_263),
.C(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_304),
.C(n_303),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_271),
.B(n_265),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_288),
.B(n_280),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_263),
.C(n_274),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_306),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_293),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_295),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_312),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_305),
.B(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_313),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_308),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_321),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_322),
.B(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_317),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_314),
.Y(n_327)
);


endmodule