module real_jpeg_29671_n_25 (n_17, n_123, n_8, n_0, n_21, n_2, n_125, n_10, n_9, n_12, n_124, n_24, n_6, n_121, n_23, n_11, n_14, n_7, n_22, n_18, n_3, n_117, n_119, n_5, n_4, n_122, n_1, n_20, n_19, n_118, n_126, n_16, n_15, n_13, n_120, n_25);

input n_17;
input n_123;
input n_8;
input n_0;
input n_21;
input n_2;
input n_125;
input n_10;
input n_9;
input n_12;
input n_124;
input n_24;
input n_6;
input n_121;
input n_23;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_117;
input n_119;
input n_5;
input n_4;
input n_122;
input n_1;
input n_20;
input n_19;
input n_118;
input n_126;
input n_16;
input n_15;
input n_13;
input n_120;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_0),
.Y(n_111)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_1),
.B(n_67),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_2),
.B(n_38),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_41),
.C(n_106),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_6),
.B(n_32),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_7),
.B(n_26),
.CI(n_30),
.CON(n_25),
.SN(n_25)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_8),
.B(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_9),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_10),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_11),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_12),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_13),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_13),
.B(n_76),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_15),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_16),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_18),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_18),
.B(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_20),
.B(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_21),
.B(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_22),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_45),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.B(n_114),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_88),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_99),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_34),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_109),
.B(n_113),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_108),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_102),
.B(n_105),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_97),
.B(n_101),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_92),
.C(n_96),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_91),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_90),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_85),
.B(n_89),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_84),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_79),
.B(n_83),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_75),
.B(n_78),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_74),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_68),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_71),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_77),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_81),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_112),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_117),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_118),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_119),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_120),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_121),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_122),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_123),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_124),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_125),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_126),
.Y(n_95)
);


endmodule