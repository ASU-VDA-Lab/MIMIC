module real_aes_8048_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_869;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_637;
wire n_526;
wire n_653;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_371;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_0), .A2(n_86), .B1(n_483), .B2(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_1), .A2(n_48), .B1(n_370), .B2(n_406), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_2), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_3), .A2(n_276), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_4), .A2(n_114), .B1(n_559), .B2(n_815), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_5), .A2(n_34), .B1(n_557), .B2(n_559), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_6), .A2(n_138), .B1(n_406), .B2(n_648), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_7), .A2(n_29), .B1(n_343), .B2(n_882), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_8), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_9), .A2(n_493), .B1(n_524), .B2(n_525), .Y(n_492) );
INVx1_ASAP7_75t_L g524 ( .A(n_9), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_10), .Y(n_623) );
INVx1_ASAP7_75t_L g628 ( .A(n_11), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_12), .A2(n_107), .B1(n_420), .B2(n_592), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_13), .A2(n_36), .B1(n_367), .B2(n_370), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_14), .A2(n_231), .B1(n_483), .B2(n_485), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_15), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_16), .A2(n_141), .B1(n_490), .B2(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_17), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_18), .A2(n_238), .B1(n_368), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_19), .A2(n_145), .B1(n_338), .B2(n_343), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_20), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_21), .A2(n_159), .B1(n_720), .B2(n_878), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_22), .Y(n_583) );
AOI22x1_ASAP7_75t_L g397 ( .A1(n_23), .A2(n_398), .B1(n_450), .B2(n_451), .Y(n_397) );
INVx1_ASAP7_75t_L g450 ( .A(n_23), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_24), .A2(n_140), .B1(n_682), .B2(n_728), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_25), .A2(n_274), .B1(n_350), .B2(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_26), .Y(n_569) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_27), .A2(n_102), .B1(n_312), .B2(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g855 ( .A(n_27), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_28), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_30), .A2(n_248), .B1(n_370), .B2(n_406), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_31), .A2(n_186), .B1(n_513), .B2(n_606), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_32), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_33), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_35), .A2(n_267), .B1(n_559), .B2(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_37), .A2(n_164), .B1(n_382), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_38), .A2(n_147), .B1(n_606), .B2(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g837 ( .A1(n_39), .A2(n_53), .B1(n_361), .B2(n_678), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_40), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_41), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_42), .A2(n_203), .B1(n_463), .B2(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_43), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_44), .B(n_437), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_45), .Y(n_798) );
INVx1_ASAP7_75t_L g616 ( .A(n_46), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_47), .Y(n_626) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_49), .A2(n_103), .B1(n_312), .B2(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g856 ( .A(n_49), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_50), .A2(n_210), .B1(n_410), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_51), .A2(n_111), .B1(n_406), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_52), .A2(n_113), .B1(n_463), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_54), .A2(n_255), .B1(n_554), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_55), .A2(n_170), .B1(n_368), .B2(n_679), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_56), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_57), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_58), .A2(n_206), .B1(n_480), .B2(n_483), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_59), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_60), .B(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_61), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_62), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_63), .A2(n_216), .B1(n_419), .B2(n_708), .Y(n_778) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_64), .A2(n_132), .B1(n_606), .B2(n_908), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_65), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_66), .A2(n_101), .B1(n_389), .B2(n_480), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_67), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_68), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_69), .A2(n_121), .B1(n_402), .B2(n_411), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_70), .A2(n_269), .B1(n_430), .B2(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_71), .A2(n_225), .B1(n_382), .B2(n_912), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_72), .A2(n_235), .B1(n_438), .B2(n_490), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_73), .A2(n_240), .B1(n_651), .B2(n_652), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_74), .A2(n_178), .B1(n_611), .B2(n_612), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_75), .A2(n_143), .B1(n_409), .B2(n_410), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_76), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_77), .A2(n_182), .B1(n_475), .B2(n_548), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_78), .B(n_437), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_79), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_80), .A2(n_200), .B1(n_592), .B2(n_866), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_81), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_82), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_83), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_84), .A2(n_148), .B1(n_338), .B2(n_431), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_85), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_87), .Y(n_870) );
INVx1_ASAP7_75t_L g892 ( .A(n_88), .Y(n_892) );
XOR2x2_ASAP7_75t_L g894 ( .A(n_88), .B(n_895), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_89), .A2(n_139), .B1(n_389), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_90), .A2(n_228), .B1(n_545), .B2(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_91), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_92), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_93), .A2(n_196), .B1(n_485), .B2(n_557), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_94), .Y(n_380) );
AOI222xp33_ASAP7_75t_L g486 ( .A1(n_95), .A2(n_169), .B1(n_175), .B2(n_487), .C1(n_489), .C2(n_490), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_96), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_97), .A2(n_98), .B1(n_480), .B2(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_99), .A2(n_197), .B1(n_483), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_100), .A2(n_162), .B1(n_476), .B2(n_576), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_104), .A2(n_263), .B1(n_548), .B2(n_549), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_105), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_106), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_108), .A2(n_176), .B1(n_367), .B2(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g293 ( .A(n_109), .Y(n_293) );
INVx1_ASAP7_75t_L g508 ( .A(n_110), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_112), .A2(n_259), .B1(n_552), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_115), .A2(n_201), .B1(n_418), .B2(n_420), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_116), .A2(n_202), .B1(n_730), .B2(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_117), .Y(n_562) );
INVx1_ASAP7_75t_L g290 ( .A(n_118), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_119), .A2(n_179), .B1(n_387), .B2(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g506 ( .A(n_120), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_122), .A2(n_163), .B1(n_361), .B2(n_612), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_123), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_124), .A2(n_273), .B1(n_339), .B2(n_343), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_125), .A2(n_243), .B1(n_589), .B2(n_682), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_126), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_127), .A2(n_198), .B1(n_561), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_128), .A2(n_251), .B1(n_829), .B2(n_885), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_129), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_130), .A2(n_134), .B1(n_343), .B2(n_475), .Y(n_673) );
OA22x2_ASAP7_75t_L g660 ( .A1(n_131), .A2(n_661), .B1(n_662), .B2(n_684), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_131), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_133), .A2(n_233), .B1(n_736), .B2(n_737), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_135), .B(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_136), .A2(n_227), .B1(n_485), .B2(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_137), .B(n_546), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_142), .A2(n_144), .B1(n_461), .B2(n_463), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_146), .A2(n_149), .B1(n_517), .B2(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_150), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_151), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_152), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_153), .B(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_154), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_155), .A2(n_241), .B1(n_648), .B2(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g294 ( .A(n_156), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_157), .B(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_158), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_160), .A2(n_602), .B1(n_629), .B2(n_630), .Y(n_601) );
INVx1_ASAP7_75t_L g629 ( .A(n_160), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_161), .B(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_165), .A2(n_218), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_166), .Y(n_403) );
AND2x6_ASAP7_75t_L g289 ( .A(n_167), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_167), .Y(n_849) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_168), .A2(n_230), .B1(n_312), .B2(n_316), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_171), .A2(n_189), .B1(n_611), .B2(n_612), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_172), .A2(n_250), .B1(n_574), .B2(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_173), .B(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_174), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_177), .A2(n_859), .B1(n_860), .B2(n_886), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_177), .Y(n_886) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_180), .A2(n_264), .B1(n_368), .B2(n_648), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_181), .A2(n_193), .B1(n_476), .B2(n_667), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_183), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_184), .B(n_574), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_185), .A2(n_213), .B1(n_361), .B2(n_362), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_187), .A2(n_257), .B1(n_517), .B2(n_682), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_188), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_190), .A2(n_285), .B1(n_409), .B2(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g715 ( .A(n_191), .Y(n_715) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_192), .A2(n_253), .B1(n_312), .B2(n_313), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_194), .B(n_670), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_195), .A2(n_278), .B1(n_521), .B2(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_SL g710 ( .A1(n_199), .A2(n_711), .B1(n_739), .B2(n_740), .Y(n_710) );
INVx1_ASAP7_75t_L g740 ( .A(n_199), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_204), .A2(n_749), .B1(n_770), .B2(n_771), .Y(n_748) );
INVx1_ASAP7_75t_L g770 ( .A(n_204), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_205), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_207), .A2(n_232), .B1(n_678), .B2(n_679), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_208), .A2(n_244), .B1(n_378), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_209), .A2(n_256), .B1(n_338), .B2(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_211), .A2(n_229), .B1(n_338), .B2(n_343), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_212), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_214), .Y(n_416) );
INVx1_ASAP7_75t_L g718 ( .A(n_215), .Y(n_718) );
AOI22xp33_ASAP7_75t_SL g913 ( .A1(n_217), .A2(n_280), .B1(n_414), .B2(n_587), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_219), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_220), .A2(n_242), .B1(n_463), .B2(n_731), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_221), .B(n_471), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_222), .A2(n_260), .B1(n_343), .B2(n_438), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_223), .B(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_224), .Y(n_391) );
INVx1_ASAP7_75t_L g714 ( .A(n_226), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_230), .B(n_854), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_234), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_236), .A2(n_272), .B1(n_420), .B2(n_463), .Y(n_514) );
INVx1_ASAP7_75t_L g774 ( .A(n_237), .Y(n_774) );
INVx1_ASAP7_75t_L g654 ( .A(n_239), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_245), .Y(n_709) );
INVx1_ASAP7_75t_L g717 ( .A(n_246), .Y(n_717) );
OA22x2_ASAP7_75t_L g792 ( .A1(n_247), .A2(n_793), .B1(n_794), .B2(n_817), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_247), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_249), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_252), .B(n_438), .Y(n_504) );
INVx1_ASAP7_75t_L g852 ( .A(n_253), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_254), .Y(n_538) );
INVx1_ASAP7_75t_L g722 ( .A(n_258), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_261), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_262), .Y(n_376) );
INVx1_ASAP7_75t_L g312 ( .A(n_265), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_265), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_266), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_268), .Y(n_759) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_270), .A2(n_287), .B(n_295), .C(n_857), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_271), .Y(n_354) );
OA22x2_ASAP7_75t_L g300 ( .A1(n_275), .A2(n_301), .B1(n_302), .B2(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
INVx1_ASAP7_75t_L g723 ( .A(n_277), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_279), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_281), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_282), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_283), .B(n_546), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_284), .Y(n_501) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_290), .Y(n_848) );
OA21x2_ASAP7_75t_L g890 ( .A1(n_291), .A2(n_847), .B(n_891), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_656), .B1(n_842), .B2(n_843), .C(n_844), .Y(n_295) );
INVx1_ASAP7_75t_L g842 ( .A(n_296), .Y(n_842) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_529), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_396), .B2(n_528), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_358), .Y(n_303) );
NOR3xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_329), .C(n_347), .Y(n_304) );
OAI22xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_322), .B1(n_323), .B2(n_328), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_306), .A2(n_637), .B1(n_714), .B2(n_715), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_306), .A2(n_323), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_308), .Y(n_426) );
BUFx3_ASAP7_75t_L g497 ( .A(n_308), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_308), .A2(n_325), .B1(n_784), .B2(n_785), .C(n_786), .Y(n_783) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
INVx2_ASAP7_75t_L g390 ( .A(n_309), .Y(n_390) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_315), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_310), .B(n_315), .Y(n_327) );
AND2x2_ASAP7_75t_L g369 ( .A(n_310), .B(n_353), .Y(n_369) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g334 ( .A(n_311), .B(n_315), .Y(n_334) );
AND2x2_ASAP7_75t_L g342 ( .A(n_311), .B(n_321), .Y(n_342) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_314), .Y(n_316) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
INVx1_ASAP7_75t_L g373 ( .A(n_315), .Y(n_373) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_318), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g368 ( .A(n_318), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g473 ( .A(n_318), .B(n_390), .Y(n_473) );
AND2x6_ASAP7_75t_L g543 ( .A(n_318), .B(n_327), .Y(n_543) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
INVx1_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
INVx1_ASAP7_75t_L g346 ( .A(n_319), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_319), .B(n_321), .Y(n_374) );
AND2x2_ASAP7_75t_L g335 ( .A(n_320), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g365 ( .A(n_321), .B(n_346), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_323), .A2(n_423), .B1(n_424), .B2(n_427), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_323), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_323), .A2(n_424), .B1(n_578), .B2(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_325), .A2(n_426), .B1(n_616), .B2(n_617), .Y(n_615) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g469 ( .A(n_326), .Y(n_469) );
AND2x4_ASAP7_75t_L g361 ( .A(n_327), .B(n_335), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_327), .B(n_365), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B(n_337), .Y(n_329) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_331), .A2(n_665), .B(n_666), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g787 ( .A1(n_331), .A2(n_788), .B(n_789), .Y(n_787) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_333), .Y(n_434) );
INVx4_ASAP7_75t_L g488 ( .A(n_333), .Y(n_488) );
INVx2_ASAP7_75t_L g500 ( .A(n_333), .Y(n_500) );
INVx2_ASAP7_75t_L g822 ( .A(n_333), .Y(n_822) );
AND2x6_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x4_ASAP7_75t_L g344 ( .A(n_334), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g448 ( .A(n_334), .Y(n_448) );
AND2x2_ASAP7_75t_L g379 ( .A(n_335), .B(n_369), .Y(n_379) );
AND2x6_ASAP7_75t_L g389 ( .A(n_335), .B(n_390), .Y(n_389) );
BUFx4f_ASAP7_75t_SL g489 ( .A(n_338), .Y(n_489) );
INVx2_ASAP7_75t_L g901 ( .A(n_338), .Y(n_901) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_339), .Y(n_438) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_339), .Y(n_571) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g352 ( .A(n_341), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g351 ( .A(n_342), .B(n_352), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_342), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g476 ( .A(n_342), .B(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_SL g490 ( .A(n_344), .Y(n_490) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_344), .Y(n_576) );
INVx1_ASAP7_75t_L g449 ( .A(n_345), .Y(n_449) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_354), .B2(n_355), .Y(n_347) );
OAI221xp5_ASAP7_75t_SL g754 ( .A1(n_349), .A2(n_619), .B1(n_755), .B2(n_756), .C(n_757), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_351), .Y(n_431) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_351), .Y(n_548) );
BUFx2_ASAP7_75t_L g622 ( .A(n_351), .Y(n_622) );
BUFx4f_ASAP7_75t_SL g667 ( .A(n_351), .Y(n_667) );
INVx1_ASAP7_75t_L g357 ( .A(n_353), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_355), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_580) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx4_ASAP7_75t_L g443 ( .A(n_356), .Y(n_443) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_356), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_356), .A2(n_502), .B1(n_642), .B2(n_643), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_356), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
AND2x2_ASAP7_75t_L g708 ( .A(n_357), .B(n_384), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_375), .C(n_385), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_366), .Y(n_359) );
BUFx3_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
INVx6_ASAP7_75t_L g462 ( .A(n_361), .Y(n_462) );
BUFx3_ASAP7_75t_L g611 ( .A(n_361), .Y(n_611) );
BUFx3_ASAP7_75t_L g781 ( .A(n_361), .Y(n_781) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx5_ASAP7_75t_L g419 ( .A(n_363), .Y(n_419) );
BUFx3_ASAP7_75t_L g464 ( .A(n_363), .Y(n_464) );
INVx3_ASAP7_75t_L g652 ( .A(n_363), .Y(n_652) );
INVx4_ASAP7_75t_L g678 ( .A(n_363), .Y(n_678) );
INVx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_365), .B(n_369), .Y(n_395) );
AND2x2_ASAP7_75t_L g481 ( .A(n_365), .B(n_369), .Y(n_481) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_368), .Y(n_523) );
BUFx3_ASAP7_75t_L g594 ( .A(n_368), .Y(n_594) );
INVx2_ASAP7_75t_L g607 ( .A(n_368), .Y(n_607) );
AND2x4_ASAP7_75t_L g383 ( .A(n_369), .B(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_371), .Y(n_420) );
BUFx2_ASAP7_75t_L g554 ( .A(n_371), .Y(n_554) );
BUFx2_ASAP7_75t_L g731 ( .A(n_371), .Y(n_731) );
BUFx2_ASAP7_75t_L g866 ( .A(n_371), .Y(n_866) );
INVx6_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g679 ( .A(n_372), .Y(n_679) );
INVx1_ASAP7_75t_SL g812 ( .A(n_372), .Y(n_812) );
OR2x6_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g477 ( .A(n_373), .Y(n_477) );
INVx1_ASAP7_75t_L g384 ( .A(n_374), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_380), .B2(n_381), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
INVx2_ASAP7_75t_L g484 ( .A(n_379), .Y(n_484) );
BUFx2_ASAP7_75t_SL g908 ( .A(n_379), .Y(n_908) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
BUFx3_ASAP7_75t_L g485 ( .A(n_383), .Y(n_485) );
BUFx2_ASAP7_75t_SL g561 ( .A(n_383), .Y(n_561) );
BUFx2_ASAP7_75t_L g648 ( .A(n_383), .Y(n_648) );
BUFx3_ASAP7_75t_L g835 ( .A(n_383), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx4_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
INVx2_ASAP7_75t_L g734 ( .A(n_388), .Y(n_734) );
INVx5_ASAP7_75t_SL g815 ( .A(n_388), .Y(n_815) );
INVx11_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx11_ASAP7_75t_L g558 ( .A(n_389), .Y(n_558) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_393), .A2(n_413), .B1(n_415), .B2(n_416), .C(n_417), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_393), .A2(n_462), .B1(n_872), .B2(n_873), .Y(n_871) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g528 ( .A(n_396), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_452), .B1(n_453), .B2(n_527), .Y(n_396) );
INVx2_ASAP7_75t_L g527 ( .A(n_397), .Y(n_527) );
INVx1_ASAP7_75t_SL g451 ( .A(n_398), .Y(n_451) );
AND2x2_ASAP7_75t_SL g398 ( .A(n_399), .B(n_421), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_412), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B1(n_404), .B2(n_407), .C(n_408), .Y(n_400) );
INVx2_ASAP7_75t_L g810 ( .A(n_401), .Y(n_810) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx3_ASAP7_75t_L g513 ( .A(n_402), .Y(n_513) );
BUFx3_ASAP7_75t_L g728 ( .A(n_402), .Y(n_728) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_402), .Y(n_864) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g769 ( .A(n_411), .Y(n_769) );
INVx2_ASAP7_75t_L g736 ( .A(n_413), .Y(n_736) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_419), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_428), .C(n_440), .Y(n_421) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI222xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B1(n_433), .B2(n_435), .C1(n_436), .C2(n_439), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g502 ( .A(n_430), .Y(n_502) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g582 ( .A(n_431), .Y(n_582) );
OAI222xp33_ASAP7_75t_L g796 ( .A1(n_433), .A2(n_797), .B1(n_798), .B2(n_799), .C1(n_800), .C2(n_801), .Y(n_796) );
OAI21xp5_ASAP7_75t_SL g897 ( .A1(n_433), .A2(n_898), .B(n_899), .Y(n_897) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g568 ( .A(n_434), .Y(n_568) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_444), .B2(n_445), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_SL g507 ( .A(n_443), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_445), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_445), .A2(n_507), .B1(n_759), .B2(n_760), .Y(n_758) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g724 ( .A(n_446), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
OR2x6_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_455), .B1(n_492), .B2(n_526), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
XOR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_491), .Y(n_457) );
NAND4xp75_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .C(n_478), .D(n_486), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_465), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
INVx2_ASAP7_75t_L g552 ( .A(n_462), .Y(n_552) );
INVx2_ASAP7_75t_L g651 ( .A(n_462), .Y(n_651) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OA211x2_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .C(n_474), .Y(n_466) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g637 ( .A(n_469), .Y(n_637) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx5_ASAP7_75t_L g546 ( .A(n_472), .Y(n_546) );
INVx2_ASAP7_75t_L g827 ( .A(n_472), .Y(n_827) );
INVx2_ASAP7_75t_L g885 ( .A(n_472), .Y(n_885) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g549 ( .A(n_476), .Y(n_549) );
BUFx2_ASAP7_75t_L g804 ( .A(n_476), .Y(n_804) );
INVx1_ASAP7_75t_L g883 ( .A(n_476), .Y(n_883) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g519 ( .A(n_480), .Y(n_519) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g559 ( .A(n_481), .Y(n_559) );
BUFx3_ASAP7_75t_L g703 ( .A(n_481), .Y(n_703) );
BUFx3_ASAP7_75t_L g912 ( .A(n_481), .Y(n_912) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g589 ( .A(n_484), .Y(n_589) );
INVx2_ASAP7_75t_L g619 ( .A(n_487), .Y(n_619) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_488), .A2(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g526 ( .A(n_492), .Y(n_526) );
INVx2_ASAP7_75t_L g525 ( .A(n_493), .Y(n_525) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_494), .B(n_510), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .C(n_505), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_497), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_502), .B2(n_503), .C(n_504), .Y(n_499) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_500), .A2(n_538), .B(n_539), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_520), .Y(n_515) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_522), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_867) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_597), .B2(n_598), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_533), .B1(n_563), .B2(n_596), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
XOR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_562), .Y(n_534) );
NAND3x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_550), .C(n_555), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .C(n_547), .Y(n_540) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g671 ( .A(n_543), .Y(n_671) );
BUFx4f_ASAP7_75t_L g698 ( .A(n_543), .Y(n_698) );
BUFx2_ASAP7_75t_L g829 ( .A(n_543), .Y(n_829) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g797 ( .A(n_548), .Y(n_797) );
INVx4_ASAP7_75t_L g879 ( .A(n_548), .Y(n_879) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .Y(n_555) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_SL g587 ( .A(n_558), .Y(n_587) );
INVx4_ASAP7_75t_L g682 ( .A(n_558), .Y(n_682) );
BUFx3_ASAP7_75t_L g612 ( .A(n_559), .Y(n_612) );
INVx1_ASAP7_75t_L g596 ( .A(n_563), .Y(n_596) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
XOR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_595), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_584), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_577), .C(n_580), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_572), .C(n_573), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_568), .A2(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_571), .Y(n_720) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B1(n_631), .B2(n_655), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g630 ( .A(n_602), .Y(n_630) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_603), .B(n_614), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_609), .Y(n_603) );
NAND2xp33_ASAP7_75t_SL g604 ( .A(n_605), .B(n_608), .Y(n_604) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .C(n_625), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_620), .B1(n_621), .B2(n_623), .C(n_624), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g716 ( .A1(n_619), .A2(n_621), .B1(n_717), .B2(n_718), .C(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g655 ( .A(n_631), .Y(n_655) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_654), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_644), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_638), .C(n_641), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_649), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
INVx1_ASAP7_75t_L g843 ( .A(n_656), .Y(n_843) );
AOI22xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B1(n_742), .B2(n_743), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_685), .B1(n_686), .B2(n_741), .Y(n_658) );
INVx1_ASAP7_75t_L g741 ( .A(n_659), .Y(n_741) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g684 ( .A(n_662), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_674), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .C(n_673), .Y(n_668) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g806 ( .A(n_671), .Y(n_806) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_680), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_678), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx4_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
XOR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_710), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
XOR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_709), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_700), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .C(n_699), .Y(n_695) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_705), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g738 ( .A(n_703), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_SL g739 ( .A(n_711), .Y(n_739) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_712), .B(n_725), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_716), .C(n_721), .Y(n_712) );
INVx1_ASAP7_75t_L g800 ( .A(n_720), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_732), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_744), .A2(n_745), .B1(n_790), .B2(n_791), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_747), .A2(n_748), .B1(n_772), .B2(n_773), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g771 ( .A(n_749), .Y(n_771) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_761), .Y(n_749) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .C(n_758), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
XNOR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
NOR4xp75_ASAP7_75t_L g775 ( .A(n_776), .B(n_779), .C(n_783), .D(n_787), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_818), .B1(n_840), .B2(n_841), .Y(n_791) );
INVx1_ASAP7_75t_L g840 ( .A(n_792), .Y(n_840) );
INVx1_ASAP7_75t_SL g817 ( .A(n_794), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_807), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_802), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_813), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g869 ( .A(n_815), .Y(n_869) );
INVx3_ASAP7_75t_L g841 ( .A(n_818), .Y(n_841) );
XOR2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_839), .Y(n_818) );
NAND2x1_ASAP7_75t_SL g819 ( .A(n_820), .B(n_831), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_825), .Y(n_820) );
OAI21xp5_ASAP7_75t_SL g821 ( .A1(n_822), .A2(n_823), .B(n_824), .Y(n_821) );
OAI21xp5_ASAP7_75t_SL g875 ( .A1(n_822), .A2(n_876), .B(n_877), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .C(n_830), .Y(n_825) );
NOR2x1_ASAP7_75t_L g831 ( .A(n_832), .B(n_836), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx1_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
NOR2x1_ASAP7_75t_L g845 ( .A(n_846), .B(n_850), .Y(n_845) );
OR2x2_ASAP7_75t_SL g916 ( .A(n_846), .B(n_851), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_849), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
OAI322xp33_ASAP7_75t_L g857 ( .A1(n_848), .A2(n_858), .A3(n_887), .B1(n_890), .B2(n_892), .C1(n_893), .C2(n_914), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_848), .B(n_889), .Y(n_891) );
CKINVDCx16_ASAP7_75t_R g889 ( .A(n_849), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_861), .B(n_874), .Y(n_860) );
NOR3xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_867), .C(n_871), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_865), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_880), .Y(n_874) );
INVx3_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_884), .Y(n_880) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_906), .C(n_910), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_902), .Y(n_896) );
INVx3_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .C(n_905), .Y(n_902) );
AND2x2_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .Y(n_906) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_913), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_915), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
endmodule