module fake_jpeg_411_n_453 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_5),
.B(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_54),
.Y(n_148)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_23),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_75),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_29),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_89),
.Y(n_118)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_42),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_18),
.B(n_14),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_29),
.B(n_13),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_18),
.B(n_13),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_41),
.B1(n_22),
.B2(n_42),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_95),
.A2(n_47),
.B1(n_79),
.B2(n_72),
.Y(n_169)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_41),
.CON(n_105),
.SN(n_105)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_105),
.B(n_26),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_120),
.A2(n_135),
.B1(n_147),
.B2(n_57),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_55),
.B(n_21),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_123),
.B(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_48),
.B(n_21),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_41),
.B1(n_22),
.B2(n_31),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_139),
.B1(n_73),
.B2(n_78),
.Y(n_166)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_134),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_31),
.B1(n_43),
.B2(n_22),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_43),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_136),
.B(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_54),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_49),
.A2(n_22),
.B1(n_45),
.B2(n_40),
.Y(n_139)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_53),
.B(n_45),
.Y(n_144)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_50),
.Y(n_145)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_22),
.B1(n_26),
.B2(n_36),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_84),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_165),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_62),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_166),
.B(n_172),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_65),
.C(n_86),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_137),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_156),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_159),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_82),
.C(n_44),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_77),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_82),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_37),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_37),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_167),
.B(n_174),
.Y(n_242)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_169),
.A2(n_141),
.B1(n_113),
.B2(n_125),
.Y(n_230)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_117),
.A2(n_34),
.B1(n_27),
.B2(n_44),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_101),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_36),
.B(n_34),
.C(n_27),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_180),
.Y(n_233)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_108),
.B(n_14),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_106),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_190),
.Y(n_237)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_105),
.A2(n_87),
.B1(n_56),
.B2(n_81),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_194),
.B1(n_199),
.B2(n_68),
.Y(n_226)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_193),
.Y(n_209)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_94),
.B(n_12),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_195),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_139),
.A2(n_76),
.B(n_64),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_131),
.A2(n_60),
.B1(n_66),
.B2(n_51),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_142),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_61),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_198),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_78),
.B1(n_68),
.B2(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_112),
.B(n_12),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_126),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_94),
.A3(n_127),
.B1(n_17),
.B2(n_33),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_157),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_217),
.B(n_234),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_115),
.B1(n_103),
.B2(n_113),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_243),
.B1(n_194),
.B2(n_195),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_226),
.A2(n_230),
.B1(n_127),
.B2(n_163),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_115),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_231),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_103),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_153),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_119),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_239),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_152),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_155),
.B(n_119),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_189),
.A2(n_193),
.B1(n_187),
.B2(n_149),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_244),
.B(n_182),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_174),
.B(n_141),
.C(n_125),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_187),
.C(n_152),
.Y(n_247)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_247),
.B(n_215),
.Y(n_311)
);

BUFx8_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_248),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_264),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_250),
.A2(n_265),
.B1(n_266),
.B2(n_241),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_245),
.Y(n_290)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_154),
.B1(n_196),
.B2(n_176),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_253),
.A2(n_17),
.B1(n_182),
.B2(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_183),
.B(n_156),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_254),
.A2(n_259),
.B(n_274),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_165),
.B(n_161),
.C(n_167),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_255),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_220),
.A2(n_196),
.B(n_168),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_242),
.B(n_184),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_262),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_202),
.B(n_181),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g309 ( 
.A1(n_263),
.A2(n_203),
.B1(n_215),
.B2(n_241),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_229),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_170),
.B1(n_186),
.B2(n_175),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_177),
.B1(n_150),
.B2(n_158),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_205),
.B1(n_231),
.B2(n_240),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_269),
.B(n_272),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_278),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_190),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_273),
.B(n_277),
.Y(n_319)
);

AND2x4_ASAP7_75t_SL g274 ( 
.A(n_207),
.B(n_158),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_209),
.A2(n_173),
.B(n_171),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_210),
.B(n_235),
.Y(n_292)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_212),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_150),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_0),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_253),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_217),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_224),
.B(n_188),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_202),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_211),
.C(n_219),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_286),
.A2(n_312),
.B1(n_249),
.B2(n_250),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_311),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_297),
.B(n_271),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_295),
.B(n_299),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_227),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_304),
.C(n_305),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_210),
.B(n_214),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_216),
.A3(n_235),
.B1(n_234),
.B2(n_232),
.C1(n_211),
.C2(n_221),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_228),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_219),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_218),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_315),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_309),
.A2(n_248),
.B1(n_278),
.B2(n_265),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_223),
.C(n_218),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_203),
.C(n_232),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_252),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_1),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_276),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_274),
.B1(n_256),
.B2(n_246),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_275),
.A2(n_1),
.B(n_2),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_266),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_297),
.A2(n_248),
.B(n_259),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_321),
.A2(n_328),
.B(n_288),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_327),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_264),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_335),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_281),
.B1(n_255),
.B2(n_247),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_339),
.A2(n_315),
.B1(n_294),
.B2(n_295),
.Y(n_359)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_342),
.B(n_343),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_291),
.A2(n_269),
.B1(n_277),
.B2(n_273),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_318),
.B1(n_317),
.B2(n_320),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_314),
.Y(n_342)
);

AOI32xp33_ASAP7_75t_L g343 ( 
.A1(n_306),
.A2(n_274),
.A3(n_248),
.B1(n_258),
.B2(n_257),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_330),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_345),
.A2(n_346),
.B1(n_349),
.B2(n_298),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_310),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_286),
.A2(n_279),
.B1(n_4),
.B2(n_5),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_304),
.C(n_311),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_357),
.C(n_360),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_358),
.B1(n_373),
.B2(n_374),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_356),
.A2(n_333),
.B(n_338),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_308),
.B1(n_312),
.B2(n_290),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_345),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_305),
.C(n_307),
.Y(n_360)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_296),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_366),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_313),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_288),
.C(n_292),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_344),
.C(n_322),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_339),
.A2(n_302),
.B1(n_287),
.B2(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_323),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_301),
.B1(n_287),
.B2(n_318),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_366),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_385),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_378),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_367),
.A2(n_325),
.B1(n_324),
.B2(n_321),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_379),
.B(n_381),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_368),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_367),
.A2(n_335),
.B1(n_329),
.B2(n_322),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_384),
.A2(n_390),
.B1(n_374),
.B2(n_377),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_368),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_386),
.B(n_6),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_320),
.C(n_346),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_391),
.C(n_394),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_309),
.C(n_327),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_352),
.A2(n_327),
.B1(n_309),
.B2(n_6),
.Y(n_392)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_392),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_3),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_3),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_3),
.C(n_5),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_369),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_398),
.Y(n_413)
);

OAI31xp33_ASAP7_75t_SL g396 ( 
.A1(n_388),
.A2(n_365),
.A3(n_356),
.B(n_373),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_378),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_358),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_380),
.A2(n_354),
.B(n_355),
.Y(n_400)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_408),
.Y(n_418)
);

OAI321xp33_ASAP7_75t_L g405 ( 
.A1(n_384),
.A2(n_359),
.A3(n_370),
.B1(n_362),
.B2(n_371),
.C(n_351),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_405),
.B(n_387),
.Y(n_414)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_362),
.C(n_353),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_410),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_411),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_380),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_416),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_414),
.A2(n_403),
.B1(n_8),
.B2(n_9),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_404),
.B(n_375),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_375),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_417),
.B(n_395),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_420),
.A2(n_421),
.B(n_396),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_402),
.A2(n_391),
.B(n_385),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_389),
.C(n_393),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_423),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_394),
.C(n_8),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_426),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_409),
.C(n_406),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_406),
.C(n_402),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_433),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_397),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_428),
.B(n_434),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_420),
.Y(n_438)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_7),
.C(n_9),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_7),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_423),
.Y(n_443)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_432),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_440),
.B(n_415),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_427),
.A2(n_418),
.B(n_424),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_426),
.B(n_430),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_443),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_445),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_435),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_442),
.Y(n_447)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g449 ( 
.A1(n_447),
.A2(n_438),
.B(n_441),
.C(n_439),
.D(n_433),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_446),
.B(n_448),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_437),
.C(n_436),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_415),
.Y(n_453)
);


endmodule