module fake_netlist_6_4412_n_2035 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2035);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2035;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_76),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_12),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_58),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_8),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_147),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_105),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_77),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_100),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_93),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_26),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_43),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_28),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_131),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_3),
.Y(n_227)
);

CKINVDCx11_ASAP7_75t_R g228 ( 
.A(n_30),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_28),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_36),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_63),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_164),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_95),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_62),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_167),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_187),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_2),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_65),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_85),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_96),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_143),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_5),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_39),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_62),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_159),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_90),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_189),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_182),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_29),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_8),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_68),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_184),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_70),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_80),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_26),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_174),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_103),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_121),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_113),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_59),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_109),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_51),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_129),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_165),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_125),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_92),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_179),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_171),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_46),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_18),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_73),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_74),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_120),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_66),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_38),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_110),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_139),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_117),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_56),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_106),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_115),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_94),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_192),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_40),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_1),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_108),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_38),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_10),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_146),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_83),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_87),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_173),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_57),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_193),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_145),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_86),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_19),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_41),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_124),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_37),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_69),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_14),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_149),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_7),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_154),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_4),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_155),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_175),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_89),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_4),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_11),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_190),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_183),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_3),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_18),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_48),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_5),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_114),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_130),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_102),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_79),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_172),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_185),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_63),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_111),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_10),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_23),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_107),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_144),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_54),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_9),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_178),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_152),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_34),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_123),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_133),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_97),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_47),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_58),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_42),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_40),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_13),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_61),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_24),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_162),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_166),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_198),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_33),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_51),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_53),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_53),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_75),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_157),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_50),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_37),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_168),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_35),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_65),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_98),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_116),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_21),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_141),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_140),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_104),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_151),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_52),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_136),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_7),
.Y(n_389)
);

CKINVDCx11_ASAP7_75t_R g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_46),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_11),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_160),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_169),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_68),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_43),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_204),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_211),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_226),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_243),
.B(n_218),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_228),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_0),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_274),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_309),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_279),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_214),
.B(n_0),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_390),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_214),
.B(n_1),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_234),
.B(n_14),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_333),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_242),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_267),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_333),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_267),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_383),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_245),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_267),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_224),
.B(n_15),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_267),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_274),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_250),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_267),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_300),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_252),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_300),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_300),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_300),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_300),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_387),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_254),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

BUFx6f_ASAP7_75t_SL g443 ( 
.A(n_374),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_199),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_199),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_206),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_234),
.B(n_258),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_248),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_262),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_266),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_248),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_310),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_269),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_387),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_272),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_206),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_275),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_310),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_229),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_278),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_259),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_259),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_281),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_338),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_302),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_282),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_302),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_286),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_287),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_322),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_290),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_256),
.B(n_15),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_291),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_320),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_292),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_294),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_297),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_298),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_320),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_306),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_308),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_314),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_200),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_227),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_317),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_230),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_327),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_337),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_202),
.B(n_16),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_237),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_340),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_258),
.B(n_16),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_466),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_201),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_424),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_401),
.B(n_331),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_399),
.A2(n_241),
.B1(n_392),
.B2(n_376),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_430),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_405),
.B(n_322),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_404),
.A2(n_409),
.B(n_402),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_398),
.B(n_248),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

BUFx8_ASAP7_75t_L g522 ( 
.A(n_443),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_236),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_417),
.B(n_201),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_417),
.B(n_236),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_409),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_441),
.B(n_307),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_434),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_435),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_435),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_499),
.B(n_205),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_408),
.B(n_342),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_436),
.B(n_307),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

BUFx8_ASAP7_75t_SL g541 ( 
.A(n_403),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_419),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_437),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_412),
.B(n_205),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_428),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_419),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_420),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_413),
.B(n_207),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_428),
.B(n_311),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_454),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_457),
.B(n_311),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_452),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_452),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_457),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_411),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_420),
.B(n_207),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_459),
.Y(n_565)
);

AND3x2_ASAP7_75t_L g566 ( 
.A(n_496),
.B(n_381),
.C(n_332),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_400),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_489),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_463),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_480),
.B(n_208),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_490),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_480),
.B(n_208),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_464),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_460),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_509),
.B(n_445),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_548),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_538),
.B(n_548),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_502),
.Y(n_586)
);

XOR2x2_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_444),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_509),
.B(n_332),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_538),
.B(n_416),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_506),
.B(n_423),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_510),
.B(n_407),
.C(n_418),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_543),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_559),
.A2(n_453),
.B1(n_474),
.B2(n_449),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_548),
.B(n_429),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_541),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_559),
.B(n_446),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_508),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_566),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_563),
.B(n_381),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_533),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_502),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_559),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_508),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_433),
.Y(n_608)
);

CKINVDCx6p67_ASAP7_75t_R g609 ( 
.A(n_562),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_567),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_533),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_575),
.B(n_577),
.C(n_546),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_519),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_533),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_503),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_537),
.B(n_440),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_524),
.B(n_450),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_563),
.B(n_524),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_503),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_556),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_503),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_518),
.A2(n_496),
.B1(n_431),
.B2(n_442),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_560),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_544),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_503),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_540),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_518),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_560),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_556),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_556),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_544),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_541),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_560),
.B(n_456),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_537),
.B(n_455),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_524),
.B(n_490),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_519),
.A2(n_443),
.B1(n_406),
.B2(n_422),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_544),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_521),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_521),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_521),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_567),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_570),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_570),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_549),
.Y(n_652)
);

BUFx6f_ASAP7_75t_SL g653 ( 
.A(n_568),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_562),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_570),
.B(n_458),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_579),
.A2(n_487),
.B1(n_492),
.B2(n_481),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_579),
.B(n_448),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_579),
.B(n_517),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_568),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_518),
.A2(n_202),
.B1(n_425),
.B2(n_255),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_549),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_549),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_528),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_517),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_546),
.B(n_233),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_518),
.A2(n_249),
.B1(n_270),
.B2(n_268),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_522),
.B(n_494),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_508),
.Y(n_669)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_512),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_551),
.B(n_517),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_549),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_551),
.B(n_233),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_518),
.B(n_462),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_527),
.A2(n_389),
.B1(n_351),
.B2(n_316),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_549),
.B(n_465),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_522),
.B(n_498),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_575),
.B(n_473),
.C(n_468),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_530),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_526),
.B(n_477),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_526),
.B(n_233),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_530),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_512),
.A2(n_486),
.B1(n_495),
.B2(n_482),
.Y(n_684)
);

XOR2xp5_ASAP7_75t_L g685 ( 
.A(n_577),
.B(n_479),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_540),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_527),
.B(n_233),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_530),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_562),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_528),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_530),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_562),
.B(n_289),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_522),
.B(n_374),
.Y(n_693)
);

BUFx4f_ASAP7_75t_L g694 ( 
.A(n_540),
.Y(n_694)
);

INVx6_ASAP7_75t_L g695 ( 
.A(n_522),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_540),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_500),
.B(n_483),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_527),
.B(n_233),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_508),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_528),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_500),
.B(n_484),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_572),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_540),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_572),
.A2(n_361),
.B1(n_280),
.B2(n_334),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_576),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_522),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_540),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_527),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_576),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_505),
.B(n_488),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_528),
.B(n_343),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_529),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_529),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_529),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_529),
.B(n_534),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_505),
.B(n_443),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_534),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_539),
.B(n_263),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_540),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_539),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_534),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_534),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_550),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_550),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_539),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_539),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_550),
.B(n_345),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_550),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_540),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_507),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_539),
.B(n_263),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_621),
.B(n_558),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_667),
.B(n_338),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_658),
.B(n_451),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_682),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_621),
.B(n_558),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_674),
.B(n_263),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_683),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_614),
.B(n_263),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_665),
.B(n_263),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_692),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_641),
.B(n_558),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_588),
.A2(n_370),
.B(n_284),
.C(n_301),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_580),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_603),
.B(n_273),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_581),
.B(n_273),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_588),
.A2(n_288),
.B(n_330),
.C(n_304),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_641),
.B(n_558),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_704),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_660),
.A2(n_271),
.B1(n_209),
.B2(n_212),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_581),
.A2(n_341),
.B1(n_239),
.B2(n_238),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_704),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_590),
.B(n_558),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_709),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_504),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_597),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_655),
.B(n_485),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_504),
.Y(n_759)
);

AO22x2_ASAP7_75t_L g760 ( 
.A1(n_607),
.A2(n_329),
.B1(n_344),
.B2(n_339),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_589),
.A2(n_377),
.B1(n_239),
.B2(n_238),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_608),
.B(n_504),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_651),
.B(n_485),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_589),
.B(n_617),
.C(n_591),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_653),
.B(n_222),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_671),
.B(n_504),
.Y(n_766)
);

BUFx5_ASAP7_75t_L g767 ( 
.A(n_612),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_688),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_671),
.B(n_210),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_709),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_585),
.B(n_504),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_623),
.B(n_507),
.Y(n_772)
);

HB1xp67_ASAP7_75t_SL g773 ( 
.A(n_597),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_691),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_640),
.B(n_491),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_623),
.B(n_511),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_625),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_649),
.B(n_478),
.C(n_426),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_L g779 ( 
.A(n_628),
.B(n_493),
.C(n_491),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_583),
.B(n_511),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_625),
.B(n_513),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_627),
.B(n_253),
.C(n_247),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_580),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_586),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_636),
.B(n_513),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_679),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_679),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_657),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_607),
.B(n_273),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_670),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_636),
.B(n_514),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_637),
.B(n_514),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_637),
.B(n_515),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_586),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_622),
.B(n_515),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_607),
.B(n_273),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_604),
.Y(n_797)
);

BUFx8_ASAP7_75t_L g798 ( 
.A(n_653),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_680),
.B(n_516),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_604),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_721),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_619),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_634),
.A2(n_335),
.B1(n_336),
.B2(n_350),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_721),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_642),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_634),
.A2(n_283),
.B1(n_273),
.B2(n_303),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_642),
.B(n_493),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_642),
.A2(n_367),
.B1(n_219),
.B2(n_215),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_706),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_634),
.A2(n_221),
.B1(n_313),
.B2(n_220),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_605),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_605),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_598),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_702),
.B(n_497),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_726),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_676),
.B(n_283),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_666),
.A2(n_283),
.B1(n_303),
.B2(n_338),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_611),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_727),
.A2(n_295),
.B1(n_217),
.B2(n_216),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_697),
.B(n_701),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_710),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_605),
.B(n_697),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_701),
.B(n_516),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_711),
.B(n_283),
.Y(n_825)
);

AOI221xp5_ASAP7_75t_L g826 ( 
.A1(n_705),
.A2(n_395),
.B1(n_362),
.B2(n_360),
.C(n_359),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_678),
.B(n_210),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_666),
.A2(n_283),
.B1(n_303),
.B2(n_338),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_711),
.B(n_582),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_584),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_613),
.B(n_303),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_635),
.B(n_497),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_592),
.B(n_520),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_596),
.B(n_520),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_687),
.B(n_203),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_731),
.B(n_532),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_703),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_615),
.B(n_303),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_639),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_601),
.B(n_532),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_650),
.B(n_670),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_685),
.A2(n_215),
.B1(n_348),
.B2(n_349),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_656),
.B(n_222),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_601),
.B(n_536),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_593),
.B(n_225),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_673),
.A2(n_338),
.B1(n_276),
.B2(n_394),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_695),
.B(n_374),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_620),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_618),
.B(n_338),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_629),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_624),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_692),
.B(n_213),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_624),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_639),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_631),
.B(n_536),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_626),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_626),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_659),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_633),
.B(n_542),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_638),
.B(n_338),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_673),
.A2(n_338),
.B1(n_264),
.B2(n_277),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_L g862 ( 
.A(n_594),
.B(n_219),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_717),
.B(n_574),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_703),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_645),
.B(n_542),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_611),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_652),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_661),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_717),
.B(n_574),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_599),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_663),
.Y(n_871)
);

OR2x6_ASAP7_75t_SL g872 ( 
.A(n_654),
.B(n_225),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_630),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_672),
.B(n_223),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_684),
.B(n_235),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_692),
.B(n_231),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_630),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_720),
.A2(n_547),
.B(n_545),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_712),
.B(n_244),
.Y(n_879)
);

OAI22xp33_ASAP7_75t_L g880 ( 
.A1(n_693),
.A2(n_359),
.B1(n_240),
.B2(n_232),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_609),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_681),
.A2(n_246),
.B1(n_388),
.B2(n_380),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_643),
.Y(n_883)
);

AO22x2_ASAP7_75t_L g884 ( 
.A1(n_587),
.A2(n_324),
.B1(n_326),
.B2(n_328),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_675),
.A2(n_574),
.B(n_564),
.C(n_571),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_687),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_643),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_728),
.B(n_545),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_595),
.B(n_600),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_703),
.B(n_348),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_646),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_698),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_668),
.A2(n_362),
.B1(n_232),
.B2(n_240),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_602),
.B(n_547),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_698),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_644),
.B(n_285),
.C(n_296),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_703),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_692),
.B(n_265),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_599),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_599),
.B(n_251),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_595),
.B(n_600),
.Y(n_901)
);

AND2x2_ASAP7_75t_SL g902 ( 
.A(n_677),
.B(n_260),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_599),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_595),
.B(n_265),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_786),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_733),
.A2(n_694),
.B(n_716),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_737),
.A2(n_694),
.B(n_681),
.Y(n_907)
);

O2A1O1Ixp5_ASAP7_75t_L g908 ( 
.A1(n_747),
.A2(n_732),
.B(n_719),
.C(n_602),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_789),
.A2(n_715),
.B(n_713),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_820),
.A2(n_352),
.B(n_356),
.C(n_366),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_743),
.A2(n_719),
.B(n_732),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_749),
.A2(n_754),
.B(n_789),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_796),
.A2(n_738),
.B(n_766),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_796),
.A2(n_708),
.B(n_696),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_829),
.B(n_602),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_786),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_742),
.B(n_695),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_738),
.A2(n_723),
.B(n_722),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_799),
.B(n_729),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_756),
.A2(n_708),
.B(n_696),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_841),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_824),
.B(n_646),
.Y(n_922)
);

BUFx10_ASAP7_75t_L g923 ( 
.A(n_757),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_805),
.B(n_777),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_827),
.A2(n_654),
.B1(n_689),
.B2(n_347),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_786),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_759),
.A2(n_708),
.B(n_696),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_769),
.A2(n_700),
.B(n_725),
.C(n_724),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_736),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_795),
.B(n_647),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_769),
.B(n_647),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_805),
.B(n_600),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_777),
.B(n_707),
.Y(n_933)
);

NOR2x1_ASAP7_75t_L g934 ( 
.A(n_823),
.B(n_707),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_818),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_762),
.A2(n_664),
.B(n_648),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_790),
.B(n_659),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_806),
.B(n_648),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_806),
.B(n_664),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_740),
.A2(n_700),
.B(n_690),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_739),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_815),
.B(n_606),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_758),
.B(n_690),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_739),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_747),
.A2(n_714),
.B(n_725),
.C(n_724),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_815),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_786),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_823),
.B(n_349),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_787),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_771),
.A2(n_714),
.B(n_718),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_735),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_825),
.A2(n_718),
.B(n_501),
.C(n_535),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_809),
.B(n_606),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_751),
.A2(n_553),
.B(n_554),
.C(n_555),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_768),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_821),
.B(n_606),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_816),
.A2(n_557),
.B(n_501),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_787),
.B(n_353),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_807),
.B(n_804),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_866),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_888),
.A2(n_610),
.B(n_699),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_815),
.B(n_606),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_787),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_750),
.A2(n_587),
.B1(n_695),
.B2(n_699),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_740),
.A2(n_730),
.B(n_686),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_790),
.B(n_609),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_768),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_815),
.B(n_610),
.Y(n_968)
);

AO21x1_ASAP7_75t_L g969 ( 
.A1(n_825),
.A2(n_535),
.B(n_501),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_787),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_772),
.A2(n_616),
.B(n_699),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_866),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_781),
.B(n_610),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_785),
.B(n_610),
.Y(n_974)
);

AND2x2_ASAP7_75t_SL g975 ( 
.A(n_902),
.B(n_847),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_791),
.B(n_616),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_792),
.B(n_616),
.Y(n_977)
);

CKINVDCx6p67_ASAP7_75t_R g978 ( 
.A(n_872),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_798),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_793),
.B(n_616),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_863),
.B(n_662),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_782),
.A2(n_730),
.B(n_686),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_776),
.A2(n_699),
.B(n_669),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_L g984 ( 
.A1(n_827),
.A2(n_845),
.B(n_889),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_886),
.A2(n_730),
.B(n_686),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_788),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_734),
.A2(n_669),
.B(n_662),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_813),
.B(n_761),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_774),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_889),
.B(n_662),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_901),
.B(n_662),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_863),
.B(n_669),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_774),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_763),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_816),
.A2(n_669),
.B(n_686),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_869),
.B(n_830),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_803),
.A2(n_810),
.B1(n_875),
.B2(n_892),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_894),
.A2(n_632),
.B(n_730),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_780),
.A2(n_632),
.B(n_730),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_869),
.B(n_564),
.Y(n_1000)
);

INVx8_ASAP7_75t_L g1001 ( 
.A(n_742),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_840),
.A2(n_632),
.B(n_552),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_814),
.B(n_564),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_844),
.A2(n_632),
.B(n_552),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_814),
.B(n_807),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_753),
.A2(n_353),
.B1(n_355),
.B2(n_373),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_811),
.B(n_355),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_850),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_803),
.B(n_801),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_741),
.A2(n_561),
.B(n_553),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_755),
.B(n_564),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_770),
.B(n_564),
.Y(n_1012)
);

OAI321xp33_ASAP7_75t_L g1013 ( 
.A1(n_880),
.A2(n_469),
.A3(n_464),
.B1(n_467),
.B2(n_470),
.C(n_471),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_775),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_812),
.B(n_357),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_741),
.A2(n_554),
.B(n_555),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_832),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_804),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_870),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_836),
.B(n_569),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_901),
.B(n_357),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_837),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_867),
.Y(n_1023)
);

AO21x1_ASAP7_75t_L g1024 ( 
.A1(n_875),
.A2(n_525),
.B(n_535),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_895),
.B(n_569),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_822),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_849),
.A2(n_561),
.B(n_525),
.Y(n_1027)
);

AND2x6_ASAP7_75t_L g1028 ( 
.A(n_898),
.B(n_525),
.Y(n_1028)
);

NOR2x1p5_ASAP7_75t_SL g1029 ( 
.A(n_767),
.B(n_557),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_849),
.A2(n_860),
.B(n_859),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_868),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_764),
.A2(n_879),
.B1(n_862),
.B2(n_871),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_843),
.B(n_231),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_882),
.A2(n_752),
.B1(n_808),
.B2(n_861),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_822),
.B(n_569),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_852),
.B(n_467),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_744),
.A2(n_569),
.B(n_571),
.C(n_367),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_853),
.B(n_569),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_837),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_833),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_853),
.B(n_571),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_904),
.B(n_265),
.Y(n_1042)
);

AND3x2_ASAP7_75t_L g1043 ( 
.A(n_858),
.B(n_476),
.C(n_472),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_860),
.A2(n_557),
.B(n_565),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_880),
.B(n_377),
.C(n_373),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_873),
.A2(n_877),
.B(n_878),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_873),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_877),
.B(n_571),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_855),
.A2(n_578),
.B(n_565),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_879),
.B(n_571),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_865),
.A2(n_578),
.B(n_565),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_834),
.A2(n_899),
.B(n_874),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_767),
.B(n_368),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_745),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_767),
.B(n_368),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_783),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_882),
.A2(n_385),
.B1(n_386),
.B2(n_384),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_899),
.A2(n_578),
.B(n_565),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_900),
.A2(n_578),
.B(n_531),
.C(n_469),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_767),
.B(n_784),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_899),
.A2(n_874),
.B(n_797),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_902),
.B(n_384),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_870),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_794),
.Y(n_1064)
);

CKINVDCx10_ASAP7_75t_R g1065 ( 
.A(n_773),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_876),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_767),
.B(n_385),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_899),
.A2(n_523),
.B(n_531),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_852),
.B(n_531),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_767),
.B(n_386),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_800),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_885),
.A2(n_476),
.B(n_472),
.C(n_471),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_802),
.B(n_393),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_778),
.B(n_470),
.Y(n_1074)
);

CKINVDCx11_ASAP7_75t_R g1075 ( 
.A(n_742),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_765),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_848),
.A2(n_523),
.B(n_531),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_779),
.B(n_346),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_851),
.B(n_393),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_748),
.A2(n_257),
.B(n_261),
.C(n_293),
.Y(n_1080)
);

AO21x1_ASAP7_75t_L g1081 ( 
.A1(n_900),
.A2(n_17),
.B(n_19),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_837),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_842),
.B(n_299),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_852),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_893),
.B(n_305),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_839),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_856),
.A2(n_523),
.B(n_531),
.Y(n_1087)
);

AO21x1_ASAP7_75t_L g1088 ( 
.A1(n_835),
.A2(n_17),
.B(n_20),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_SL g1089 ( 
.A(n_854),
.B(n_346),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_857),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_883),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_887),
.A2(n_523),
.B(n_312),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_837),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_893),
.B(n_315),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_884),
.B(n_573),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1014),
.B(n_896),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_941),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_1086),
.B(n_881),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_960),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_929),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_984),
.B(n_864),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_SL g1102 ( 
.A1(n_910),
.A2(n_885),
.B(n_838),
.C(n_831),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_951),
.B(n_819),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_975),
.A2(n_884),
.B1(n_890),
.B2(n_760),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_905),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_959),
.B(n_903),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_986),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_912),
.A2(n_913),
.B(n_907),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1040),
.B(n_760),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_997),
.A2(n_1034),
.B1(n_1095),
.B2(n_1009),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_905),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1085),
.A2(n_861),
.B(n_846),
.C(n_826),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_972),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1001),
.B(n_884),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_935),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_967),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_SL g1117 ( 
.A(n_1083),
.B(n_391),
.C(n_395),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1095),
.A2(n_828),
.B1(n_817),
.B2(n_760),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_912),
.A2(n_897),
.B(n_864),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_996),
.B(n_891),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1095),
.A2(n_817),
.B1(n_828),
.B2(n_846),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_988),
.A2(n_835),
.B1(n_903),
.B2(n_897),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_917),
.B(n_916),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_907),
.A2(n_864),
.B(n_838),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_SL g1125 ( 
.A1(n_938),
.A2(n_831),
.B(n_864),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_973),
.A2(n_523),
.B(n_573),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_959),
.B(n_798),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_994),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_974),
.A2(n_523),
.B(n_573),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_944),
.Y(n_1130)
);

NOR2x1p5_ASAP7_75t_SL g1131 ( 
.A(n_918),
.B(n_746),
.Y(n_1131)
);

AND3x1_ASAP7_75t_SL g1132 ( 
.A(n_1008),
.B(n_360),
.C(n_382),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_1075),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_976),
.A2(n_523),
.B(n_573),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1094),
.A2(n_746),
.B1(n_573),
.B2(n_318),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1005),
.B(n_71),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1082),
.Y(n_1137)
);

AND3x2_ASAP7_75t_L g1138 ( 
.A(n_1045),
.B(n_347),
.C(n_354),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_923),
.B(n_354),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_922),
.B(n_573),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_977),
.A2(n_523),
.B(n_573),
.Y(n_1141)
);

AOI21x1_ASAP7_75t_L g1142 ( 
.A1(n_931),
.A2(n_906),
.B(n_920),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_955),
.Y(n_1143)
);

CKINVDCx10_ASAP7_75t_R g1144 ( 
.A(n_1065),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1017),
.B(n_319),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_990),
.A2(n_746),
.B(n_72),
.C(n_81),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1032),
.A2(n_321),
.B(n_323),
.C(n_379),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_980),
.A2(n_911),
.B(n_914),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_909),
.A2(n_985),
.B(n_906),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_905),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_911),
.A2(n_523),
.B(n_573),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_921),
.B(n_391),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1062),
.A2(n_382),
.B(n_379),
.C(n_371),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_914),
.A2(n_746),
.B(n_156),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1030),
.A2(n_371),
.B(n_369),
.C(n_365),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_948),
.A2(n_369),
.B(n_365),
.C(n_22),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_989),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1042),
.B(n_20),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_919),
.B(n_746),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_993),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_920),
.A2(n_197),
.B(n_196),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_SL g1162 ( 
.A1(n_1080),
.A2(n_195),
.B(n_194),
.C(n_180),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_939),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1021),
.B(n_25),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_936),
.A2(n_170),
.B(n_163),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_930),
.B(n_150),
.Y(n_1166)
);

XOR2x2_ASAP7_75t_SL g1167 ( 
.A(n_1057),
.B(n_27),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_958),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1066),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1033),
.B(n_31),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_923),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1013),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_927),
.A2(n_134),
.B(n_127),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1082),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_964),
.B(n_947),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1001),
.B(n_122),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1036),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_917),
.B(n_112),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1023),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_969),
.A2(n_101),
.B(n_91),
.C(n_88),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_947),
.B(n_84),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1076),
.B(n_32),
.Y(n_1182)
);

BUFx4f_ASAP7_75t_SL g1183 ( 
.A(n_979),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1030),
.A2(n_35),
.B(n_36),
.C(n_39),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_SL g1185 ( 
.A(n_1018),
.B(n_41),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1026),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1031),
.Y(n_1187)
);

CKINVDCx16_ASAP7_75t_R g1188 ( 
.A(n_1089),
.Y(n_1188)
);

OR2x6_ASAP7_75t_SL g1189 ( 
.A(n_1073),
.B(n_42),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1043),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1082),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_947),
.Y(n_1192)
);

AO21x1_ASAP7_75t_L g1193 ( 
.A1(n_961),
.A2(n_44),
.B(n_45),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_927),
.A2(n_82),
.B(n_47),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1047),
.Y(n_1195)
);

AO21x1_ASAP7_75t_L g1196 ( 
.A1(n_961),
.A2(n_44),
.B(n_49),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_943),
.B(n_49),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_917),
.B(n_916),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_937),
.B(n_52),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_962),
.A2(n_70),
.B(n_56),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_991),
.B(n_55),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_968),
.A2(n_915),
.B(n_1060),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_963),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_971),
.A2(n_57),
.B(n_59),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_908),
.A2(n_60),
.B(n_64),
.C(n_67),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1074),
.Y(n_1206)
);

CKINVDCx10_ASAP7_75t_R g1207 ( 
.A(n_978),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1007),
.A2(n_60),
.B(n_64),
.C(n_67),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1003),
.A2(n_1029),
.B(n_1000),
.C(n_1067),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_963),
.B(n_69),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_971),
.A2(n_983),
.B(n_987),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_963),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_946),
.B(n_1018),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1054),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1020),
.B(n_981),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1093),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1056),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1001),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1015),
.A2(n_1037),
.B(n_932),
.C(n_1079),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_992),
.B(n_970),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_936),
.A2(n_957),
.B(n_1052),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_966),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1078),
.B(n_933),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_983),
.A2(n_987),
.B(n_1092),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1084),
.Y(n_1225)
);

OR2x4_ASAP7_75t_L g1226 ( 
.A(n_1093),
.B(n_925),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1093),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_924),
.A2(n_1072),
.B(n_1088),
.C(n_1053),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_970),
.B(n_1090),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1052),
.A2(n_1046),
.B(n_942),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1055),
.B(n_1070),
.Y(n_1231)
);

OR2x6_ASAP7_75t_SL g1232 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_R g1233 ( 
.A(n_1019),
.B(n_1063),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_942),
.A2(n_956),
.B(n_953),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_982),
.A2(n_965),
.B(n_950),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_SL g1236 ( 
.A(n_926),
.B(n_949),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1036),
.B(n_934),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1028),
.B(n_926),
.Y(n_1238)
);

BUFx4f_ASAP7_75t_L g1239 ( 
.A(n_1028),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_949),
.A2(n_1006),
.B1(n_1025),
.B2(n_1091),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1028),
.A2(n_1081),
.B1(n_1069),
.B2(n_1024),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1019),
.Y(n_1242)
);

AOI21xp33_ASAP7_75t_L g1243 ( 
.A1(n_954),
.A2(n_1050),
.B(n_1011),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_950),
.A2(n_1022),
.B(n_1039),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1028),
.B(n_1063),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1012),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_928),
.A2(n_1039),
.B1(n_1022),
.B2(n_1041),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1028),
.A2(n_1027),
.B1(n_1044),
.B2(n_1035),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_999),
.A2(n_1061),
.B(n_940),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1061),
.B(n_1038),
.Y(n_1250)
);

INVxp67_ASAP7_75t_SL g1251 ( 
.A(n_1048),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_999),
.A2(n_998),
.B(n_995),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1027),
.A2(n_1016),
.B1(n_1010),
.B2(n_1002),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_952),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1002),
.B(n_1004),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1049),
.B(n_1051),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1059),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1231),
.A2(n_995),
.B(n_945),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1223),
.B(n_1004),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1211),
.A2(n_945),
.B(n_1058),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1115),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1110),
.B(n_1051),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1230),
.A2(n_998),
.B(n_1049),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_SL g1264 ( 
.A1(n_1112),
.A2(n_1077),
.B(n_1087),
.C(n_1010),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1107),
.B(n_1016),
.Y(n_1265)
);

AOI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1110),
.A2(n_1044),
.B(n_1087),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1164),
.A2(n_1077),
.B(n_1058),
.C(n_1068),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1099),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1144),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1165),
.A2(n_1068),
.B1(n_1163),
.B2(n_1184),
.C(n_1108),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1235),
.A2(n_1148),
.B(n_1249),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1169),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1255),
.A2(n_1253),
.A3(n_1224),
.B(n_1252),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1215),
.B(n_1120),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1206),
.A2(n_1117),
.B1(n_1237),
.B2(n_1222),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1142),
.A2(n_1256),
.B(n_1221),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1170),
.A2(n_1147),
.B(n_1199),
.C(n_1158),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1165),
.A2(n_1202),
.B(n_1124),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1119),
.A2(n_1215),
.B(n_1166),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1246),
.B(n_1109),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1253),
.A2(n_1196),
.A3(n_1193),
.B(n_1205),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1125),
.A2(n_1209),
.B(n_1243),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1188),
.B(n_1128),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1187),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1177),
.B(n_1145),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1243),
.A2(n_1228),
.B(n_1166),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1113),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_L g1288 ( 
.A1(n_1201),
.A2(n_1101),
.B(n_1175),
.C(n_1185),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1247),
.A2(n_1118),
.A3(n_1155),
.B(n_1121),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1109),
.B(n_1103),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1232),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_SL g1292 ( 
.A1(n_1181),
.A2(n_1118),
.B(n_1121),
.C(n_1172),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1244),
.A2(n_1250),
.B(n_1234),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1225),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1152),
.B(n_1182),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1219),
.A2(n_1153),
.B(n_1104),
.C(n_1156),
.Y(n_1296)
);

AOI221xp5_ASAP7_75t_L g1297 ( 
.A1(n_1163),
.A2(n_1208),
.B1(n_1168),
.B2(n_1139),
.C(n_1200),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1096),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1197),
.B(n_1251),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1100),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1116),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1210),
.A2(n_1204),
.B(n_1162),
.C(n_1240),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1136),
.B(n_1106),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1149),
.A2(n_1140),
.B(n_1213),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1239),
.B(n_1123),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1123),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1220),
.B(n_1097),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1140),
.A2(n_1248),
.B(n_1159),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1137),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1194),
.A2(n_1136),
.B(n_1122),
.C(n_1239),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1247),
.A2(n_1240),
.A3(n_1151),
.B(n_1159),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1154),
.A2(n_1161),
.A3(n_1173),
.B(n_1220),
.Y(n_1313)
);

O2A1O1Ixp5_ASAP7_75t_SL g1314 ( 
.A1(n_1254),
.A2(n_1130),
.B(n_1157),
.C(n_1143),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1254),
.A2(n_1129),
.B(n_1134),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1126),
.A2(n_1141),
.B(n_1238),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1180),
.A2(n_1102),
.B(n_1241),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1229),
.A2(n_1149),
.B(n_1245),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1146),
.A2(n_1203),
.B(n_1257),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1186),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1257),
.A2(n_1198),
.B(n_1106),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1257),
.A2(n_1198),
.B(n_1178),
.Y(n_1322)
);

AO21x2_ASAP7_75t_L g1323 ( 
.A1(n_1233),
.A2(n_1195),
.B(n_1160),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1218),
.B(n_1178),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1214),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1217),
.Y(n_1326)
);

OAI22x1_ASAP7_75t_L g1327 ( 
.A1(n_1167),
.A2(n_1127),
.B1(n_1190),
.B2(n_1242),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1150),
.A2(n_1212),
.B(n_1192),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1150),
.A2(n_1212),
.B(n_1192),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1226),
.A2(n_1114),
.B1(n_1176),
.B2(n_1135),
.Y(n_1330)
);

BUFx2_ASAP7_75t_SL g1331 ( 
.A(n_1171),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1176),
.A2(n_1105),
.B(n_1111),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1131),
.A2(n_1236),
.B(n_1105),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1132),
.A2(n_1226),
.B(n_1138),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1176),
.B(n_1111),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1174),
.A2(n_1216),
.B(n_1191),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1114),
.B(n_1189),
.Y(n_1337)
);

OR2x6_ASAP7_75t_L g1338 ( 
.A(n_1133),
.B(n_1114),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1174),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1191),
.A2(n_1216),
.B(n_1227),
.C(n_1098),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1227),
.A2(n_912),
.B(n_1231),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1207),
.B(n_820),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1110),
.A2(n_912),
.B(n_1108),
.Y(n_1343)
);

O2A1O1Ixp5_ASAP7_75t_L g1344 ( 
.A1(n_1255),
.A2(n_820),
.B(n_747),
.C(n_589),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1164),
.A2(n_820),
.B(n_984),
.C(n_581),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1255),
.A2(n_1110),
.A3(n_1108),
.B(n_1235),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1099),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1255),
.A2(n_1110),
.A3(n_1108),
.B(n_1235),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1183),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1223),
.A2(n_581),
.B1(n_399),
.B2(n_406),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1188),
.B(n_984),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1110),
.A2(n_912),
.B(n_1108),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1206),
.B(n_820),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_SL g1357 ( 
.A(n_1188),
.B(n_975),
.Y(n_1357)
);

NOR2x1_ASAP7_75t_R g1358 ( 
.A(n_1133),
.B(n_597),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1110),
.B(n_820),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1218),
.B(n_1198),
.Y(n_1360)
);

AO21x1_ASAP7_75t_L g1361 ( 
.A1(n_1110),
.A2(n_820),
.B(n_1165),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1164),
.A2(n_820),
.B(n_984),
.C(n_581),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1118),
.A2(n_806),
.B1(n_820),
.B2(n_1121),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1255),
.A2(n_1110),
.A3(n_1108),
.B(n_1235),
.Y(n_1364)
);

AOI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1170),
.A2(n_581),
.B1(n_509),
.B2(n_401),
.C(n_1085),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1115),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1231),
.A2(n_912),
.B(n_1230),
.Y(n_1367)
);

AO32x2_ASAP7_75t_L g1368 ( 
.A1(n_1110),
.A2(n_1163),
.A3(n_1118),
.B1(n_1253),
.B2(n_1240),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1110),
.B(n_820),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1179),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1110),
.B(n_820),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1179),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1183),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1112),
.A2(n_820),
.B(n_1205),
.C(n_1184),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1110),
.B(n_820),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1198),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1179),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1198),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1110),
.B(n_820),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1110),
.B(n_820),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1218),
.B(n_1198),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1188),
.B(n_984),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_SL g1384 ( 
.A1(n_1112),
.A2(n_820),
.B(n_1205),
.C(n_1184),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1231),
.A2(n_912),
.B(n_1230),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1231),
.A2(n_912),
.B(n_1230),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1099),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1206),
.B(n_820),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1223),
.B(n_994),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1179),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1226),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1164),
.A2(n_820),
.B(n_984),
.C(n_581),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1198),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1206),
.B(n_1086),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1172),
.A2(n_1163),
.B1(n_1110),
.B2(n_1109),
.C(n_588),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1255),
.A2(n_1110),
.A3(n_1108),
.B(n_1235),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1110),
.A2(n_1163),
.B1(n_1118),
.B2(n_1121),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_SL g1399 ( 
.A1(n_1112),
.A2(n_820),
.B(n_1205),
.C(n_1184),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1183),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1223),
.B(n_820),
.Y(n_1403)
);

AOI31xp67_ASAP7_75t_L g1404 ( 
.A1(n_1101),
.A2(n_825),
.A3(n_1256),
.B(n_1250),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1206),
.B(n_820),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1211),
.A2(n_1252),
.B(n_1230),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1206),
.B(n_820),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1113),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1231),
.A2(n_912),
.B(n_1230),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1110),
.B(n_820),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1198),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1218),
.B(n_1198),
.Y(n_1412)
);

BUFx24_ASAP7_75t_L g1413 ( 
.A(n_1178),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1231),
.A2(n_912),
.B(n_1230),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1117),
.A2(n_820),
.B(n_581),
.C(n_984),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1365),
.A2(n_1295),
.B1(n_1403),
.B2(n_1297),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1372),
.Y(n_1417)
);

AOI22x1_ASAP7_75t_SL g1418 ( 
.A1(n_1298),
.A2(n_1306),
.B1(n_1351),
.B2(n_1373),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1361),
.A2(n_1398),
.B1(n_1382),
.B2(n_1353),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1274),
.B(n_1359),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1352),
.A2(n_1357),
.B1(n_1298),
.B2(n_1275),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1363),
.A2(n_1393),
.B1(n_1362),
.B2(n_1345),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1274),
.B(n_1359),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1401),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1269),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1284),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1273),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1326),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1363),
.A2(n_1357),
.B1(n_1398),
.B2(n_1330),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1327),
.A2(n_1369),
.B1(n_1410),
.B2(n_1371),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1261),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1370),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1377),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1378),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1330),
.A2(n_1342),
.B1(n_1395),
.B2(n_1337),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1369),
.A2(n_1371),
.B1(n_1375),
.B2(n_1379),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1391),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1378),
.Y(n_1438)
);

INVx8_ASAP7_75t_L g1439 ( 
.A(n_1310),
.Y(n_1439)
);

BUFx2_ASAP7_75t_SL g1440 ( 
.A(n_1366),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1375),
.A2(n_1410),
.B1(n_1380),
.B2(n_1379),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1380),
.A2(n_1259),
.B1(n_1285),
.B2(n_1389),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1265),
.A2(n_1334),
.B1(n_1290),
.B2(n_1299),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1376),
.B(n_1394),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1305),
.A2(n_1291),
.B1(n_1282),
.B2(n_1317),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1376),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1394),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1294),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1355),
.A2(n_1405),
.B1(n_1388),
.B2(n_1407),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_SL g1450 ( 
.A(n_1272),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1287),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1305),
.A2(n_1291),
.B1(n_1282),
.B2(n_1317),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1334),
.A2(n_1286),
.B1(n_1354),
.B2(n_1343),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1283),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1286),
.A2(n_1354),
.B1(n_1343),
.B2(n_1387),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1277),
.A2(n_1415),
.B1(n_1296),
.B2(n_1280),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1360),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1268),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1324),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1268),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1324),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1325),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1300),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1280),
.A2(n_1322),
.B1(n_1301),
.B2(n_1413),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1392),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1360),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1320),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1381),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1411),
.B(n_1349),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1307),
.Y(n_1470)
);

BUFx10_ASAP7_75t_L g1471 ( 
.A(n_1381),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1310),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1412),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1344),
.A2(n_1288),
.B(n_1270),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1338),
.A2(n_1303),
.B1(n_1335),
.B2(n_1408),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1338),
.A2(n_1335),
.B1(n_1323),
.B2(n_1341),
.Y(n_1476)
);

INVx8_ASAP7_75t_L g1477 ( 
.A(n_1310),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1412),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1339),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1338),
.A2(n_1262),
.B1(n_1308),
.B2(n_1321),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1336),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1262),
.A2(n_1308),
.B1(n_1278),
.B2(n_1266),
.Y(n_1482)
);

CKINVDCx6p67_ASAP7_75t_R g1483 ( 
.A(n_1331),
.Y(n_1483)
);

BUFx10_ASAP7_75t_L g1484 ( 
.A(n_1358),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1278),
.A2(n_1266),
.B1(n_1409),
.B2(n_1386),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1367),
.A2(n_1414),
.B1(n_1385),
.B2(n_1279),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1340),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1332),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1336),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1374),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1333),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1293),
.A2(n_1318),
.B1(n_1271),
.B2(n_1319),
.Y(n_1492)
);

BUFx8_ASAP7_75t_L g1493 ( 
.A(n_1368),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1328),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1329),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1264),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1271),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1396),
.A2(n_1292),
.B1(n_1311),
.B2(n_1384),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1289),
.B(n_1368),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1293),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1396),
.A2(n_1368),
.B1(n_1304),
.B2(n_1399),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1276),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1258),
.Y(n_1503)
);

INVx8_ASAP7_75t_L g1504 ( 
.A(n_1267),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1302),
.A2(n_1289),
.B1(n_1263),
.B2(n_1281),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1314),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1289),
.A2(n_1281),
.B1(n_1350),
.B2(n_1348),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1404),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1348),
.B(n_1397),
.Y(n_1509)
);

CKINVDCx11_ASAP7_75t_R g1510 ( 
.A(n_1312),
.Y(n_1510)
);

INVx6_ASAP7_75t_L g1511 ( 
.A(n_1316),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1348),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1350),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1346),
.A2(n_1406),
.B1(n_1402),
.B2(n_1400),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1347),
.A2(n_1356),
.B1(n_1390),
.B2(n_1383),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1350),
.A2(n_1364),
.B1(n_1397),
.B2(n_1260),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1397),
.B(n_1364),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1312),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1313),
.A2(n_1365),
.B(n_581),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1313),
.A2(n_1363),
.B1(n_806),
.B2(n_820),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1315),
.B(n_1313),
.Y(n_1521)
);

BUFx10_ASAP7_75t_L g1522 ( 
.A(n_1269),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1365),
.A2(n_581),
.B1(n_399),
.B2(n_406),
.Y(n_1523)
);

BUFx4f_ASAP7_75t_SL g1524 ( 
.A(n_1351),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1372),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1378),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1365),
.A2(n_1117),
.B1(n_975),
.B2(n_1295),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1365),
.A2(n_1117),
.B1(n_975),
.B2(n_1295),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1363),
.A2(n_975),
.B1(n_884),
.B2(n_519),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1378),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1365),
.A2(n_581),
.B(n_820),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1365),
.A2(n_1117),
.B1(n_975),
.B2(n_1295),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1365),
.A2(n_1117),
.B1(n_975),
.B2(n_1295),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1272),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1365),
.A2(n_1117),
.B1(n_975),
.B2(n_1295),
.Y(n_1535)
);

CKINVDCx11_ASAP7_75t_R g1536 ( 
.A(n_1351),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1274),
.B(n_1359),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1363),
.A2(n_975),
.B1(n_884),
.B2(n_519),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1372),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1372),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1363),
.A2(n_975),
.B1(n_884),
.B2(n_519),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1269),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1378),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1351),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1327),
.A2(n_1403),
.B1(n_1295),
.B2(n_1330),
.Y(n_1545)
);

BUFx4_ASAP7_75t_SL g1546 ( 
.A(n_1351),
.Y(n_1546)
);

INVx8_ASAP7_75t_L g1547 ( 
.A(n_1309),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1372),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1372),
.Y(n_1549)
);

NAND2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1378),
.B(n_1376),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1365),
.A2(n_1117),
.B1(n_975),
.B2(n_1295),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1309),
.Y(n_1552)
);

INVx3_ASAP7_75t_SL g1553 ( 
.A(n_1269),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1352),
.A2(n_820),
.B1(n_617),
.B2(n_1365),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_SL g1555 ( 
.A1(n_1363),
.A2(n_975),
.B1(n_884),
.B2(n_519),
.Y(n_1555)
);

CKINVDCx11_ASAP7_75t_R g1556 ( 
.A(n_1351),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1363),
.A2(n_975),
.B1(n_884),
.B2(n_519),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1460),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1499),
.B(n_1455),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1509),
.B(n_1507),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1508),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1511),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1489),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1493),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1509),
.B(n_1507),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1481),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1512),
.Y(n_1567)
);

NAND2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1517),
.B(n_1429),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1513),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1518),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1416),
.A2(n_1557),
.B1(n_1541),
.B2(n_1555),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1427),
.B(n_1518),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1458),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1511),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1451),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1429),
.B(n_1453),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1463),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1497),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1534),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1424),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1505),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1434),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1474),
.A2(n_1519),
.B(n_1485),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1505),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1531),
.B(n_1421),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1511),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1493),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1491),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1521),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1474),
.A2(n_1486),
.B(n_1492),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1426),
.Y(n_1592)
);

NAND3x1_ASAP7_75t_L g1593 ( 
.A(n_1435),
.B(n_1537),
.C(n_1423),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1448),
.B(n_1449),
.Y(n_1594)
);

AO31x2_ASAP7_75t_L g1595 ( 
.A1(n_1422),
.A2(n_1520),
.A3(n_1502),
.B(n_1456),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1451),
.Y(n_1596)
);

AO21x1_ASAP7_75t_SL g1597 ( 
.A1(n_1443),
.A2(n_1480),
.B(n_1430),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1503),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1432),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1496),
.Y(n_1600)
);

AO31x2_ASAP7_75t_L g1601 ( 
.A1(n_1422),
.A2(n_1520),
.A3(n_1502),
.B(n_1456),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1419),
.B(n_1482),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1488),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1494),
.B(n_1495),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1449),
.B(n_1420),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1524),
.B(n_1418),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1487),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1529),
.A2(n_1557),
.B1(n_1555),
.B2(n_1538),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1536),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1504),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1510),
.B(n_1436),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1420),
.B(n_1423),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1433),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1437),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1514),
.A2(n_1515),
.B(n_1476),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1467),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1501),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1469),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1501),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1516),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1462),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1434),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1516),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1417),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1441),
.B(n_1470),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1464),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1442),
.B(n_1554),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1445),
.B(n_1452),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1445),
.B(n_1452),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1454),
.B(n_1487),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1444),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1525),
.Y(n_1632)
);

NOR4xp25_ASAP7_75t_SL g1633 ( 
.A(n_1539),
.B(n_1540),
.C(n_1549),
.D(n_1541),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1434),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1548),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1487),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1490),
.Y(n_1637)
);

INVx11_ASAP7_75t_L g1638 ( 
.A(n_1459),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1479),
.Y(n_1639)
);

OA21x2_ASAP7_75t_L g1640 ( 
.A1(n_1506),
.A2(n_1464),
.B(n_1428),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1450),
.B(n_1473),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1444),
.A2(n_1475),
.B(n_1447),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1459),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1446),
.A2(n_1447),
.B(n_1550),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1446),
.B(n_1438),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1545),
.B(n_1538),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1550),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1478),
.Y(n_1648)
);

BUFx2_ASAP7_75t_SL g1649 ( 
.A(n_1431),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1529),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1478),
.B(n_1527),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1528),
.A2(n_1551),
.B(n_1533),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_SL g1653 ( 
.A1(n_1483),
.A2(n_1535),
.B(n_1532),
.C(n_1465),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1526),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1457),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1457),
.B(n_1468),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1468),
.A2(n_1440),
.B1(n_1461),
.B2(n_1526),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1530),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1468),
.B(n_1471),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1530),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1472),
.B(n_1552),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1543),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1543),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1466),
.B(n_1439),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1439),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1615),
.A2(n_1619),
.B(n_1617),
.Y(n_1666)
);

OA21x2_ASAP7_75t_L g1667 ( 
.A1(n_1615),
.A2(n_1547),
.B(n_1477),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1618),
.B(n_1553),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1608),
.A2(n_1572),
.B1(n_1586),
.B2(n_1652),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1594),
.A2(n_1547),
.B(n_1477),
.C(n_1546),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1592),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1611),
.B(n_1544),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1566),
.B(n_1542),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1617),
.A2(n_1477),
.B(n_1547),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1650),
.A2(n_1553),
.B1(n_1546),
.B2(n_1484),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1564),
.B(n_1556),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1646),
.A2(n_1484),
.B(n_1425),
.C(n_1522),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1571),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1638),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1564),
.B(n_1425),
.Y(n_1680)
);

INVx5_ASAP7_75t_L g1681 ( 
.A(n_1645),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1650),
.A2(n_1522),
.B1(n_1629),
.B2(n_1628),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1628),
.A2(n_1629),
.B1(n_1646),
.B2(n_1577),
.Y(n_1683)
);

O2A1O1Ixp33_ASAP7_75t_SL g1684 ( 
.A1(n_1627),
.A2(n_1581),
.B(n_1605),
.C(n_1639),
.Y(n_1684)
);

CKINVDCx6p67_ASAP7_75t_R g1685 ( 
.A(n_1643),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1603),
.B(n_1598),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1588),
.B(n_1559),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1559),
.B(n_1579),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1637),
.A2(n_1588),
.B1(n_1593),
.B2(n_1603),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1569),
.B(n_1651),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1625),
.B(n_1612),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1651),
.B(n_1626),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1577),
.A2(n_1597),
.B1(n_1626),
.B2(n_1636),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1643),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1625),
.B(n_1574),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1603),
.B(n_1636),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1637),
.A2(n_1593),
.B1(n_1607),
.B2(n_1636),
.Y(n_1697)
);

NOR3xp33_ASAP7_75t_SL g1698 ( 
.A(n_1609),
.B(n_1606),
.C(n_1657),
.Y(n_1698)
);

O2A1O1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1653),
.A2(n_1602),
.B(n_1607),
.C(n_1576),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1638),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1602),
.A2(n_1584),
.B(n_1604),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1637),
.A2(n_1607),
.B1(n_1636),
.B2(n_1633),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1630),
.B(n_1558),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1561),
.A2(n_1644),
.B(n_1589),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1640),
.B(n_1568),
.Y(n_1705)
);

INVx5_ASAP7_75t_SL g1706 ( 
.A(n_1637),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1616),
.B(n_1599),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1620),
.A2(n_1623),
.B1(n_1637),
.B2(n_1619),
.C(n_1582),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1597),
.A2(n_1610),
.B1(n_1604),
.B2(n_1584),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1613),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1584),
.A2(n_1604),
.B(n_1568),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1614),
.B(n_1582),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1637),
.A2(n_1596),
.B1(n_1585),
.B2(n_1580),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1590),
.B(n_1614),
.Y(n_1714)
);

AO32x2_ASAP7_75t_L g1715 ( 
.A1(n_1583),
.A2(n_1654),
.A3(n_1634),
.B1(n_1622),
.B2(n_1565),
.Y(n_1715)
);

AO32x2_ASAP7_75t_L g1716 ( 
.A1(n_1583),
.A2(n_1654),
.A3(n_1634),
.B1(n_1622),
.B2(n_1565),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1610),
.B(n_1563),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1640),
.B(n_1568),
.Y(n_1718)
);

NAND2x1_ASAP7_75t_L g1719 ( 
.A(n_1645),
.B(n_1562),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1563),
.B(n_1631),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1624),
.B(n_1578),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1656),
.A2(n_1641),
.B1(n_1643),
.B2(n_1649),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1642),
.A2(n_1649),
.B(n_1631),
.C(n_1560),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1584),
.A2(n_1640),
.B1(n_1600),
.B2(n_1635),
.Y(n_1725)
);

A2O1A1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1631),
.A2(n_1659),
.B(n_1663),
.C(n_1660),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1704),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1711),
.B(n_1717),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1678),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1703),
.B(n_1655),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1669),
.A2(n_1631),
.B1(n_1640),
.B2(n_1647),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1678),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1701),
.B(n_1590),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1671),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1701),
.B(n_1563),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1690),
.B(n_1567),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1686),
.B(n_1658),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1681),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1711),
.B(n_1562),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1687),
.B(n_1695),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1691),
.B(n_1595),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1666),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1710),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1691),
.B(n_1595),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1688),
.B(n_1573),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1669),
.A2(n_1591),
.B1(n_1662),
.B2(n_1648),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1689),
.B(n_1575),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1715),
.B(n_1591),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1715),
.B(n_1591),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1666),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1716),
.B(n_1591),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1717),
.B(n_1720),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1716),
.B(n_1570),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1689),
.B(n_1587),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1681),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1707),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1601),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1692),
.B(n_1705),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1712),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1705),
.B(n_1718),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1729),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1748),
.B(n_1718),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1738),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1734),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1760),
.B(n_1712),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1746),
.A2(n_1683),
.B1(n_1682),
.B2(n_1693),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1749),
.B(n_1667),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1754),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1749),
.B(n_1667),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1749),
.B(n_1718),
.Y(n_1772)
);

INVx5_ASAP7_75t_SL g1773 ( 
.A(n_1739),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1734),
.Y(n_1774)
);

OR2x6_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1719),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1750),
.B(n_1725),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1731),
.A2(n_1683),
.B1(n_1699),
.B2(n_1708),
.C(n_1677),
.Y(n_1777)
);

INVx5_ASAP7_75t_L g1778 ( 
.A(n_1738),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1761),
.Y(n_1779)
);

INVx4_ASAP7_75t_L g1780 ( 
.A(n_1738),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1727),
.Y(n_1781)
);

OAI33xp33_ASAP7_75t_L g1782 ( 
.A1(n_1741),
.A2(n_1682),
.A3(n_1713),
.B1(n_1675),
.B2(n_1697),
.B3(n_1702),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1739),
.B(n_1681),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1729),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1741),
.A2(n_1684),
.B1(n_1699),
.B2(n_1713),
.C(n_1697),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1761),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1750),
.B(n_1714),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1750),
.B(n_1723),
.Y(n_1788)
);

NAND2x1_ASAP7_75t_L g1789 ( 
.A(n_1756),
.B(n_1674),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1732),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1739),
.B(n_1756),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1752),
.A2(n_1702),
.B1(n_1706),
.B2(n_1675),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1752),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1752),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1733),
.B(n_1709),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1733),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1733),
.B(n_1595),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1760),
.B(n_1721),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1761),
.B(n_1736),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1739),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1728),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1764),
.B(n_1747),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1768),
.B(n_1787),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1798),
.B(n_1744),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1802),
.B(n_1759),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_R g1807 ( 
.A(n_1767),
.B(n_1685),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1768),
.B(n_1787),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1802),
.B(n_1759),
.Y(n_1809)
);

NAND2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1778),
.B(n_1756),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1801),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1802),
.B(n_1728),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1762),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1798),
.B(n_1744),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1801),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1768),
.B(n_1758),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1779),
.B(n_1786),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1801),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1801),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1779),
.B(n_1728),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1779),
.B(n_1728),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1795),
.B(n_1740),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1783),
.B(n_1747),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1765),
.Y(n_1824)
);

AND2x2_ASAP7_75t_SL g1825 ( 
.A(n_1785),
.B(n_1767),
.Y(n_1825)
);

NOR2x1p5_ASAP7_75t_L g1826 ( 
.A(n_1764),
.B(n_1694),
.Y(n_1826)
);

AND2x2_ASAP7_75t_SL g1827 ( 
.A(n_1785),
.B(n_1756),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_1758),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_SL g1829 ( 
.A(n_1775),
.B(n_1735),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1786),
.B(n_1740),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1765),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1786),
.B(n_1735),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1763),
.B(n_1753),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_L g1834 ( 
.A(n_1764),
.B(n_1755),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1796),
.B(n_1770),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1796),
.B(n_1745),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1765),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1781),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1783),
.B(n_1755),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1795),
.B(n_1757),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1777),
.A2(n_1696),
.B(n_1726),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1792),
.B(n_1783),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1774),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1803),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1817),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1817),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1824),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1840),
.B(n_1796),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1829),
.B(n_1788),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1804),
.B(n_1808),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1804),
.B(n_1796),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1825),
.B(n_1795),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1824),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1831),
.Y(n_1854)
);

BUFx2_ASAP7_75t_SL g1855 ( 
.A(n_1826),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1835),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1829),
.B(n_1788),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1825),
.B(n_1788),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1831),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1837),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1808),
.B(n_1766),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1837),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1834),
.B(n_1764),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1843),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1823),
.B(n_1788),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1823),
.B(n_1772),
.Y(n_1866)
);

OR2x6_ASAP7_75t_L g1867 ( 
.A(n_1810),
.B(n_1764),
.Y(n_1867)
);

NOR2x1p5_ASAP7_75t_SL g1868 ( 
.A(n_1838),
.B(n_1781),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1843),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1813),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1835),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1838),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1799),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_L g1874 ( 
.A(n_1826),
.B(n_1764),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1811),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1827),
.A2(n_1782),
.B1(n_1792),
.B2(n_1783),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1822),
.B(n_1841),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1805),
.B(n_1799),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1811),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1815),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1823),
.B(n_1772),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1839),
.B(n_1772),
.Y(n_1882)
);

NAND2x1_ASAP7_75t_L g1883 ( 
.A(n_1839),
.B(n_1800),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1839),
.B(n_1773),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1810),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1820),
.B(n_1791),
.Y(n_1886)
);

OAI21xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1842),
.A2(n_1799),
.B(n_1776),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1827),
.B(n_1679),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1816),
.B(n_1766),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1858),
.B(n_1830),
.Y(n_1890)
);

NOR2x1p5_ASAP7_75t_L g1891 ( 
.A(n_1852),
.B(n_1679),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1847),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1877),
.B(n_1830),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1873),
.B(n_1814),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1850),
.B(n_1836),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1876),
.A2(n_1827),
.B1(n_1782),
.B2(n_1791),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1874),
.B(n_1820),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1855),
.B(n_1821),
.Y(n_1898)
);

NOR2x1_ASAP7_75t_L g1899 ( 
.A(n_1863),
.B(n_1676),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1850),
.B(n_1861),
.Y(n_1900)
);

OAI31xp33_ASAP7_75t_SL g1901 ( 
.A1(n_1844),
.A2(n_1821),
.A3(n_1807),
.B(n_1812),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1847),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1859),
.Y(n_1903)
);

OR2x6_ASAP7_75t_L g1904 ( 
.A(n_1855),
.B(n_1810),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1870),
.B(n_1832),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1859),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1867),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1860),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1851),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1860),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1862),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1851),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1883),
.Y(n_1913)
);

OA21x2_ASAP7_75t_L g1914 ( 
.A1(n_1872),
.A2(n_1818),
.B(n_1815),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1861),
.B(n_1878),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1862),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1864),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1849),
.A2(n_1777),
.B1(n_1773),
.B2(n_1706),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1849),
.B(n_1812),
.Y(n_1919)
);

AND3x2_ASAP7_75t_L g1920 ( 
.A(n_1888),
.B(n_1672),
.C(n_1680),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1857),
.B(n_1865),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1889),
.B(n_1836),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1867),
.B(n_1885),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1889),
.B(n_1816),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1857),
.B(n_1806),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1865),
.B(n_1806),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1887),
.A2(n_1867),
.B(n_1883),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1921),
.B(n_1866),
.Y(n_1928)
);

OAI22xp33_ASAP7_75t_L g1929 ( 
.A1(n_1896),
.A2(n_1867),
.B1(n_1778),
.B2(n_1722),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1899),
.B(n_1885),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1893),
.B(n_1845),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1926),
.B(n_1845),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1918),
.A2(n_1884),
.B1(n_1886),
.B2(n_1882),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1901),
.A2(n_1884),
.B1(n_1846),
.B2(n_1848),
.C(n_1881),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1902),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_L g1936 ( 
.A(n_1907),
.B(n_1890),
.C(n_1927),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1902),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1892),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1903),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1906),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1926),
.B(n_1846),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1920),
.B(n_1832),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1908),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_SL g1944 ( 
.A1(n_1898),
.A2(n_1886),
.B1(n_1882),
.B2(n_1881),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1921),
.Y(n_1945)
);

NOR2xp67_ASAP7_75t_SL g1946 ( 
.A(n_1898),
.B(n_1700),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1925),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1910),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1920),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1904),
.A2(n_1730),
.B(n_1886),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1925),
.B(n_1866),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1891),
.A2(n_1698),
.B(n_1868),
.C(n_1670),
.Y(n_1952)
);

OAI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1904),
.A2(n_1923),
.B1(n_1894),
.B2(n_1900),
.Y(n_1953)
);

OR4x1_ASAP7_75t_L g1954 ( 
.A(n_1911),
.B(n_1869),
.C(n_1854),
.D(n_1853),
.Y(n_1954)
);

OAI32xp33_ASAP7_75t_L g1955 ( 
.A1(n_1949),
.A2(n_1936),
.A3(n_1930),
.B1(n_1942),
.B2(n_1945),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1945),
.B(n_1919),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1946),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1930),
.Y(n_1958)
);

NAND2xp33_ASAP7_75t_SL g1959 ( 
.A(n_1947),
.B(n_1897),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1947),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1935),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1937),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1929),
.A2(n_1904),
.B(n_1923),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1953),
.B(n_1923),
.C(n_1904),
.Y(n_1964)
);

OAI322xp33_ASAP7_75t_L g1965 ( 
.A1(n_1929),
.A2(n_1924),
.A3(n_1916),
.B1(n_1917),
.B2(n_1905),
.C1(n_1909),
.C2(n_1912),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1944),
.A2(n_1897),
.B1(n_1923),
.B2(n_1919),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1931),
.Y(n_1967)
);

NOR2x1_ASAP7_75t_L g1968 ( 
.A(n_1953),
.B(n_1952),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1933),
.A2(n_1928),
.B1(n_1951),
.B2(n_1897),
.Y(n_1969)
);

AOI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1934),
.A2(n_1924),
.B(n_1915),
.C(n_1912),
.Y(n_1970)
);

AOI222xp33_ASAP7_75t_L g1971 ( 
.A1(n_1938),
.A2(n_1909),
.B1(n_1868),
.B2(n_1776),
.C1(n_1864),
.C2(n_1797),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1939),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1940),
.Y(n_1973)
);

OAI31xp33_ASAP7_75t_L g1974 ( 
.A1(n_1952),
.A2(n_1950),
.A3(n_1932),
.B(n_1941),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1943),
.Y(n_1975)
);

AOI222xp33_ASAP7_75t_L g1976 ( 
.A1(n_1955),
.A2(n_1948),
.B1(n_1954),
.B2(n_1913),
.C1(n_1776),
.C2(n_1871),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1956),
.B(n_1895),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1960),
.Y(n_1978)
);

OAI321xp33_ASAP7_75t_L g1979 ( 
.A1(n_1964),
.A2(n_1954),
.A3(n_1922),
.B1(n_1848),
.B2(n_1871),
.C(n_1856),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1960),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1968),
.A2(n_1974),
.B1(n_1965),
.B2(n_1957),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1958),
.A2(n_1913),
.B(n_1914),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1959),
.A2(n_1913),
.B(n_1914),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1961),
.Y(n_1984)
);

O2A1O1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1962),
.A2(n_1856),
.B(n_1872),
.C(n_1668),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1967),
.B(n_1828),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1972),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1981),
.B(n_1969),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1978),
.B(n_1980),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1977),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1982),
.Y(n_1991)
);

NAND4xp25_ASAP7_75t_L g1992 ( 
.A(n_1976),
.B(n_1966),
.C(n_1970),
.D(n_1963),
.Y(n_1992)
);

A2O1A1Ixp33_ASAP7_75t_L g1993 ( 
.A1(n_1979),
.A2(n_1975),
.B(n_1973),
.C(n_1698),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1982),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1984),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1986),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1987),
.B(n_1700),
.Y(n_1997)
);

AND4x1_ASAP7_75t_L g1998 ( 
.A(n_1985),
.B(n_1971),
.C(n_1809),
.D(n_1737),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1983),
.B(n_1809),
.Y(n_1999)
);

AOI222xp33_ASAP7_75t_L g2000 ( 
.A1(n_1994),
.A2(n_1971),
.B1(n_1776),
.B2(n_1769),
.C1(n_1771),
.C2(n_1880),
.Y(n_2000)
);

NAND4xp75_ASAP7_75t_L g2001 ( 
.A(n_1988),
.B(n_1989),
.C(n_1996),
.D(n_1995),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1992),
.A2(n_1706),
.B1(n_1791),
.B2(n_1780),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1990),
.B(n_1997),
.Y(n_2003)
);

O2A1O1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1991),
.A2(n_1914),
.B(n_1880),
.C(n_1879),
.Y(n_2004)
);

AOI322xp5_ASAP7_75t_L g2005 ( 
.A1(n_1994),
.A2(n_1771),
.A3(n_1769),
.B1(n_1797),
.B2(n_1794),
.C1(n_1793),
.C2(n_1742),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_SL g2006 ( 
.A1(n_2002),
.A2(n_1991),
.B(n_1993),
.Y(n_2006)
);

OAI211xp5_ASAP7_75t_SL g2007 ( 
.A1(n_2003),
.A2(n_1998),
.B(n_1999),
.C(n_1879),
.Y(n_2007)
);

OAI31xp33_ASAP7_75t_L g2008 ( 
.A1(n_2004),
.A2(n_1673),
.A3(n_1791),
.B(n_1800),
.Y(n_2008)
);

NOR3xp33_ASAP7_75t_L g2009 ( 
.A(n_2001),
.B(n_1780),
.C(n_1673),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_L g2010 ( 
.A(n_2000),
.B(n_1875),
.Y(n_2010)
);

AOI222xp33_ASAP7_75t_L g2011 ( 
.A1(n_2005),
.A2(n_1769),
.B1(n_1771),
.B2(n_1751),
.C1(n_1875),
.C2(n_1797),
.Y(n_2011)
);

OAI21x1_ASAP7_75t_L g2012 ( 
.A1(n_2004),
.A2(n_1819),
.B(n_1818),
.Y(n_2012)
);

INVxp67_ASAP7_75t_SL g2013 ( 
.A(n_2006),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_2008),
.B(n_1828),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_2009),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_2012),
.Y(n_2016)
);

O2A1O1Ixp5_ASAP7_75t_SL g2017 ( 
.A1(n_2007),
.A2(n_1819),
.B(n_1800),
.C(n_1762),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2010),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2018),
.B(n_2013),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_2013),
.B(n_2011),
.C(n_1780),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2016),
.Y(n_2021)
);

AOI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_2015),
.A2(n_1780),
.B1(n_1800),
.B2(n_1751),
.C(n_1769),
.Y(n_2022)
);

NOR3xp33_ASAP7_75t_L g2023 ( 
.A(n_2019),
.B(n_2014),
.C(n_2017),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2023),
.A2(n_2020),
.B1(n_2022),
.B2(n_2021),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_2024),
.A2(n_1778),
.B1(n_1780),
.B2(n_1793),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2024),
.B(n_1833),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_SL g2027 ( 
.A1(n_2025),
.A2(n_1778),
.B1(n_1780),
.B2(n_1789),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2026),
.A2(n_1778),
.B1(n_1793),
.B2(n_1794),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_2027),
.A2(n_1778),
.B1(n_1793),
.B2(n_1794),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_2028),
.A2(n_1791),
.B1(n_1794),
.B2(n_1800),
.Y(n_2030)
);

OR2x6_ASAP7_75t_L g2031 ( 
.A(n_2029),
.B(n_1664),
.Y(n_2031)
);

OA21x2_ASAP7_75t_L g2032 ( 
.A1(n_2031),
.A2(n_2030),
.B(n_1665),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2032),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_2033),
.A2(n_1790),
.B1(n_1784),
.B2(n_1791),
.C(n_1800),
.Y(n_2034)
);

AOI211xp5_ASAP7_75t_L g2035 ( 
.A1(n_2034),
.A2(n_1665),
.B(n_1664),
.C(n_1661),
.Y(n_2035)
);


endmodule