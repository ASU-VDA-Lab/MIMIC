module real_aes_10993_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g167 ( .A(n_0), .Y(n_167) );
AND2x2_ASAP7_75t_L g504 ( .A(n_1), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_1), .B(n_59), .Y(n_510) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_1), .Y(n_519) );
INVx1_ASAP7_75t_L g566 ( .A(n_1), .Y(n_566) );
INVxp67_ASAP7_75t_L g552 ( .A(n_2), .Y(n_552) );
OAI222xp33_ASAP7_75t_L g601 ( .A1(n_2), .A2(n_12), .B1(n_72), .B2(n_602), .C1(n_606), .C2(n_612), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_3), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_4), .B(n_117), .Y(n_217) );
INVx2_ASAP7_75t_L g582 ( .A(n_5), .Y(n_582) );
OR2x2_ASAP7_75t_L g616 ( .A(n_5), .B(n_580), .Y(n_616) );
INVx1_ASAP7_75t_L g555 ( .A(n_6), .Y(n_555) );
INVx1_ASAP7_75t_L g503 ( .A(n_7), .Y(n_503) );
OR2x2_ASAP7_75t_L g509 ( .A(n_7), .B(n_510), .Y(n_509) );
BUFx2_ASAP7_75t_L g521 ( .A(n_7), .Y(n_521) );
INVx1_ASAP7_75t_L g478 ( .A(n_8), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_9), .Y(n_191) );
INVx1_ASAP7_75t_L g528 ( .A(n_10), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_11), .Y(n_199) );
INVxp67_ASAP7_75t_L g550 ( .A(n_12), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_13), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_14), .B(n_139), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_15), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_16), .A2(n_489), .B1(n_669), .B2(n_689), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_16), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_17), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_18), .B(n_132), .Y(n_247) );
BUFx2_ASAP7_75t_SL g476 ( .A(n_19), .Y(n_476) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_21), .B(n_134), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_22), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_23), .B(n_139), .Y(n_216) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_24), .Y(n_91) );
OAI21xp33_ASAP7_75t_L g113 ( .A1(n_25), .A2(n_114), .B(n_115), .Y(n_113) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_26), .A2(n_44), .B1(n_642), .B2(n_644), .C(n_646), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_26), .A2(n_50), .B1(n_653), .B2(n_658), .C(n_662), .Y(n_652) );
INVx1_ASAP7_75t_L g580 ( .A(n_27), .Y(n_580) );
INVx1_ASAP7_75t_L g630 ( .A(n_27), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_28), .B(n_132), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_29), .Y(n_159) );
OAI21x1_ASAP7_75t_L g107 ( .A1(n_30), .A2(n_54), .B(n_108), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_31), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_32), .B(n_132), .Y(n_131) );
INVxp67_ASAP7_75t_L g523 ( .A(n_33), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_33), .A2(n_51), .B1(n_625), .B2(n_626), .C(n_627), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_34), .Y(n_194) );
AND2x6_ASAP7_75t_L g83 ( .A(n_35), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_35), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_35), .B(n_674), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_36), .A2(n_63), .B1(n_117), .B2(n_119), .Y(n_116) );
BUFx2_ASAP7_75t_L g701 ( .A(n_36), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_37), .B(n_105), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_38), .Y(n_152) );
INVx1_ASAP7_75t_L g84 ( .A(n_39), .Y(n_84) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_39), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_40), .Y(n_226) );
OAI222xp33_ASAP7_75t_L g492 ( .A1(n_41), .A2(n_52), .B1(n_73), .B2(n_493), .C1(n_506), .C2(n_511), .Y(n_492) );
INVx1_ASAP7_75t_L g588 ( .A(n_41), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_42), .B(n_119), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_43), .B(n_119), .Y(n_245) );
OAI332xp33_ASAP7_75t_L g516 ( .A1(n_44), .A2(n_517), .A3(n_522), .B1(n_533), .B2(n_542), .B3(n_551), .C1(n_560), .C2(n_567), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_45), .B(n_145), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_46), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_47), .B(n_105), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_48), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g178 ( .A(n_49), .Y(n_178) );
INVx1_ASAP7_75t_L g640 ( .A(n_50), .Y(n_640) );
INVx1_ASAP7_75t_L g534 ( .A(n_51), .Y(n_534) );
INVx1_ASAP7_75t_L g634 ( .A(n_52), .Y(n_634) );
INVx2_ASAP7_75t_L g501 ( .A(n_53), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_55), .B(n_140), .Y(n_141) );
INVx1_ASAP7_75t_L g171 ( .A(n_56), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_57), .Y(n_202) );
BUFx10_ASAP7_75t_L g684 ( .A(n_58), .Y(n_684) );
INVx2_ASAP7_75t_L g505 ( .A(n_59), .Y(n_505) );
INVx1_ASAP7_75t_L g196 ( .A(n_60), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_61), .B(n_140), .Y(n_230) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_62), .Y(n_486) );
INVx1_ASAP7_75t_L g704 ( .A(n_63), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_64), .B(n_105), .Y(n_249) );
INVx1_ASAP7_75t_L g181 ( .A(n_65), .Y(n_181) );
INVx2_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
INVx1_ASAP7_75t_L g595 ( .A(n_67), .Y(n_595) );
INVx1_ASAP7_75t_L g539 ( .A(n_68), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_69), .Y(n_488) );
NOR2xp67_ASAP7_75t_L g110 ( .A(n_70), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g498 ( .A(n_71), .Y(n_498) );
INVxp67_ASAP7_75t_L g543 ( .A(n_72), .Y(n_543) );
INVx1_ASAP7_75t_L g599 ( .A(n_73), .Y(n_599) );
BUFx3_ASAP7_75t_L g585 ( .A(n_74), .Y(n_585) );
INVx1_ASAP7_75t_L g610 ( .A(n_74), .Y(n_610) );
BUFx3_ASAP7_75t_L g587 ( .A(n_75), .Y(n_587) );
INVx1_ASAP7_75t_L g605 ( .A(n_75), .Y(n_605) );
NAND2xp33_ASAP7_75t_L g221 ( .A(n_76), .B(n_105), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_471), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx8_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
INVx2_ASAP7_75t_SL g143 ( .A(n_82), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_82), .A2(n_145), .B(n_204), .Y(n_203) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g156 ( .A(n_83), .Y(n_156) );
AOI21xp33_ASAP7_75t_L g182 ( .A1(n_83), .A2(n_146), .B(n_180), .Y(n_182) );
INVx1_ASAP7_75t_L g233 ( .A(n_83), .Y(n_233) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g706 ( .A1(n_86), .A2(n_707), .B(n_708), .Y(n_706) );
NAND2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_90), .Y(n_114) );
INVx2_ASAP7_75t_L g119 ( .A(n_90), .Y(n_119) );
INVx2_ASAP7_75t_L g176 ( .A(n_90), .Y(n_176) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g118 ( .A(n_91), .Y(n_118) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
INVx1_ASAP7_75t_L g193 ( .A(n_91), .Y(n_193) );
OAI21xp33_ASAP7_75t_L g150 ( .A1(n_92), .A2(n_151), .B(n_155), .Y(n_150) );
INVx1_ASAP7_75t_L g218 ( .A(n_92), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_92), .A2(n_247), .B(n_248), .Y(n_246) );
INVx5_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
BUFx12f_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
INVx5_ASAP7_75t_L g136 ( .A(n_93), .Y(n_136) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND3x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_367), .C(n_434), .Y(n_96) );
NOR3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_315), .C(n_337), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g98 ( .A(n_99), .B(n_288), .Y(n_98) );
AOI221xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_183), .B1(n_252), .B2(n_270), .C(n_271), .Y(n_99) );
AND2x4_ASAP7_75t_SL g100 ( .A(n_101), .B(n_147), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_101), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_101), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g333 ( .A(n_101), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_101), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_124), .Y(n_101) );
AND2x4_ASAP7_75t_L g331 ( .A(n_102), .B(n_262), .Y(n_331) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g275 ( .A(n_103), .Y(n_275) );
AND2x4_ASAP7_75t_L g303 ( .A(n_103), .B(n_124), .Y(n_303) );
AND2x2_ASAP7_75t_L g308 ( .A(n_103), .B(n_292), .Y(n_308) );
AND2x2_ASAP7_75t_L g319 ( .A(n_103), .B(n_274), .Y(n_319) );
INVx2_ASAP7_75t_SL g346 ( .A(n_103), .Y(n_346) );
AO31x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_109), .A3(n_120), .B(n_121), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2x1p5_ASAP7_75t_SL g232 ( .A(n_105), .B(n_233), .Y(n_232) );
BUFx5_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g123 ( .A(n_106), .Y(n_123) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_113), .B1(n_115), .B2(n_116), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_115), .B(n_158), .Y(n_157) );
BUFx2_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_115), .Y(n_179) );
INVx3_ASAP7_75t_L g214 ( .A(n_115), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g151 ( .A1(n_117), .A2(n_152), .B1(n_153), .B2(n_154), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_117), .A2(n_139), .B1(n_225), .B2(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
INVx2_ASAP7_75t_L g244 ( .A(n_118), .Y(n_244) );
OAI21x1_ASAP7_75t_SL g209 ( .A1(n_120), .A2(n_210), .B(n_215), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_120), .A2(n_242), .B(n_246), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_124), .Y(n_270) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g292 ( .A(n_125), .Y(n_292) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B(n_144), .Y(n_125) );
OAI21x1_ASAP7_75t_SL g208 ( .A1(n_126), .A2(n_209), .B(n_219), .Y(n_208) );
BUFx4f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_127), .B(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g240 ( .A(n_127), .Y(n_240) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g146 ( .A(n_128), .Y(n_146) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_143), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_136), .Y(n_130) );
INVx2_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
INVx2_ASAP7_75t_L g213 ( .A(n_132), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_134), .B(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_134), .B(n_202), .Y(n_201) );
INVxp67_ASAP7_75t_L g229 ( .A(n_134), .Y(n_229) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g153 ( .A(n_135), .Y(n_153) );
INVx2_ASAP7_75t_SL g142 ( .A(n_136), .Y(n_142) );
CKINVDCx6p67_ASAP7_75t_R g223 ( .A(n_136), .Y(n_223) );
INVx2_ASAP7_75t_SL g231 ( .A(n_136), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_141), .B(n_142), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_139), .A2(n_175), .B1(n_177), .B2(n_178), .Y(n_174) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g198 ( .A(n_140), .B(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_146), .B(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_146), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g342 ( .A(n_147), .Y(n_342) );
AND2x2_ASAP7_75t_L g382 ( .A(n_147), .B(n_270), .Y(n_382) );
AND2x2_ASAP7_75t_L g408 ( .A(n_147), .B(n_379), .Y(n_408) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_163), .Y(n_147) );
AND2x2_ASAP7_75t_L g291 ( .A(n_148), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g261 ( .A(n_149), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g269 ( .A(n_149), .B(n_263), .Y(n_269) );
INVx1_ASAP7_75t_L g274 ( .A(n_149), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_149), .B(n_263), .Y(n_283) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_149), .Y(n_302) );
AND2x2_ASAP7_75t_L g332 ( .A(n_149), .B(n_292), .Y(n_332) );
AND2x4_ASAP7_75t_L g345 ( .A(n_149), .B(n_346), .Y(n_345) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_157), .B(n_162), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_153), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_158) );
AND2x2_ASAP7_75t_L g296 ( .A(n_163), .B(n_186), .Y(n_296) );
INVx2_ASAP7_75t_L g314 ( .A(n_163), .Y(n_314) );
AND2x2_ASAP7_75t_L g318 ( .A(n_163), .B(n_292), .Y(n_318) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g263 ( .A(n_164), .Y(n_263) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_173), .B(n_182), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_170), .B(n_172), .Y(n_165) );
NOR2x1_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_169), .A2(n_191), .B1(n_192), .B2(n_194), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_179), .B(n_180), .Y(n_173) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_177), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_177), .Y(n_479) );
AO21x1_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_190), .B(n_195), .Y(n_189) );
AOI21x1_ASAP7_75t_L g197 ( .A1(n_179), .A2(n_198), .B(n_200), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_184), .B(n_234), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_205), .Y(n_184) );
OR2x2_ASAP7_75t_L g268 ( .A(n_185), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g411 ( .A(n_185), .B(n_299), .Y(n_411) );
AND2x2_ASAP7_75t_L g446 ( .A(n_185), .B(n_425), .Y(n_446) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_185), .Y(n_455) );
AND2x2_ASAP7_75t_L g460 ( .A(n_185), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x4_ASAP7_75t_L g304 ( .A(n_187), .B(n_237), .Y(n_304) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
INVx1_ASAP7_75t_L g280 ( .A(n_188), .Y(n_280) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_197), .B(n_203), .Y(n_188) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_L g204 ( .A(n_195), .Y(n_204) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g277 ( .A(n_205), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g370 ( .A(n_205), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_206), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_206), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g458 ( .A(n_206), .B(n_254), .Y(n_458) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_220), .Y(n_206) );
AND2x4_ASAP7_75t_L g355 ( .A(n_207), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_207), .B(n_255), .Y(n_430) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx3_ASAP7_75t_L g267 ( .A(n_208), .Y(n_267) );
AOI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_214), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
INVx2_ASAP7_75t_L g251 ( .A(n_220), .Y(n_251) );
INVx1_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
AND2x2_ASAP7_75t_L g324 ( .A(n_220), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g356 ( .A(n_220), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_220), .B(n_259), .Y(n_419) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_227), .C(n_232), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_223), .A2(n_243), .B(n_245), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .C(n_231), .Y(n_227) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_250), .Y(n_234) );
OR2x2_ASAP7_75t_L g390 ( .A(n_235), .B(n_376), .Y(n_390) );
AND2x4_ASAP7_75t_L g461 ( .A(n_235), .B(n_355), .Y(n_461) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g265 ( .A(n_236), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_236), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_236), .B(n_251), .Y(n_287) );
AND2x4_ASAP7_75t_L g299 ( .A(n_236), .B(n_267), .Y(n_299) );
INVx1_ASAP7_75t_L g396 ( .A(n_236), .Y(n_396) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g255 ( .A(n_238), .Y(n_255) );
OAI21x1_ASAP7_75t_SL g238 ( .A1(n_239), .A2(n_241), .B(n_249), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x4_ASAP7_75t_SL g335 ( .A(n_250), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_251), .B(n_325), .Y(n_376) );
AND2x2_ASAP7_75t_L g425 ( .A(n_251), .B(n_267), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_260), .B1(n_264), .B2(n_268), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x4_ASAP7_75t_L g322 ( .A(n_254), .B(n_257), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_254), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
AND2x2_ASAP7_75t_L g420 ( .A(n_254), .B(n_418), .Y(n_420) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_254), .A2(n_465), .B(n_467), .C(n_469), .Y(n_464) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g365 ( .A(n_255), .B(n_267), .Y(n_365) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_256), .Y(n_293) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_257), .Y(n_361) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
AND2x2_ASAP7_75t_L g336 ( .A(n_259), .B(n_267), .Y(n_336) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g468 ( .A(n_261), .B(n_303), .Y(n_468) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_262), .Y(n_452) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_264), .A2(n_436), .B(n_440), .Y(n_435) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx2_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
INVx1_ASAP7_75t_L g276 ( .A(n_269), .Y(n_276) );
INVx2_ASAP7_75t_L g334 ( .A(n_269), .Y(n_334) );
INVx2_ASAP7_75t_L g379 ( .A(n_270), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_270), .Y(n_381) );
AND2x4_ASAP7_75t_L g421 ( .A(n_270), .B(n_334), .Y(n_421) );
OR2x2_ASAP7_75t_L g439 ( .A(n_270), .B(n_353), .Y(n_439) );
AND2x2_ASAP7_75t_L g449 ( .A(n_270), .B(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_277), .B1(n_281), .B2(n_284), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
AND2x2_ASAP7_75t_L g378 ( .A(n_273), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g393 ( .A(n_273), .B(n_313), .Y(n_393) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g386 ( .A(n_275), .Y(n_386) );
AND2x2_ASAP7_75t_L g380 ( .A(n_276), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g348 ( .A(n_279), .Y(n_348) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g325 ( .A(n_280), .Y(n_325) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g320 ( .A(n_282), .B(n_303), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_282), .B(n_303), .Y(n_328) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_283), .B(n_351), .Y(n_445) );
NAND2xp33_ASAP7_75t_L g416 ( .A(n_284), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g347 ( .A(n_285), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x4_ASAP7_75t_L g400 ( .A(n_286), .B(n_304), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_287), .B(n_310), .Y(n_309) );
AOI221x1_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_297), .B1(n_300), .B2(n_304), .C(n_305), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B(n_294), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g359 ( .A(n_291), .B(n_331), .Y(n_359) );
AND2x4_ASAP7_75t_L g413 ( .A(n_291), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g352 ( .A(n_292), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_292), .B(n_314), .Y(n_463) );
AND2x2_ASAP7_75t_L g437 ( .A(n_295), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_298), .A2(n_306), .B1(n_309), .B2(n_311), .Y(n_305) );
AOI332xp33_ASAP7_75t_L g392 ( .A1(n_298), .A2(n_375), .A3(n_382), .B1(n_393), .B2(n_394), .B3(n_397), .C1(n_399), .C2(n_400), .Y(n_392) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g407 ( .A(n_299), .B(n_324), .Y(n_407) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g399 ( .A(n_301), .Y(n_399) );
OR2x2_ASAP7_75t_L g432 ( .A(n_301), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g373 ( .A(n_302), .Y(n_373) );
INVx2_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
INVx1_ASAP7_75t_L g391 ( .A(n_303), .Y(n_391) );
INVx1_ASAP7_75t_L g466 ( .A(n_303), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_304), .B(n_355), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_304), .A2(n_423), .B(n_426), .C(n_431), .Y(n_422) );
INVx2_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g433 ( .A(n_308), .Y(n_433) );
INVx1_ASAP7_75t_L g371 ( .A(n_310), .Y(n_371) );
INVx1_ASAP7_75t_L g428 ( .A(n_310), .Y(n_428) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g384 ( .A1(n_313), .A2(n_385), .B(n_387), .C(n_389), .Y(n_384) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g414 ( .A(n_314), .B(n_398), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_321), .B1(n_326), .B2(n_328), .C(n_329), .Y(n_315) );
NOR2x1_ASAP7_75t_SL g316 ( .A(n_317), .B(n_320), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_317), .A2(n_359), .B1(n_360), .B2(n_362), .Y(n_358) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NOR2xp33_ASAP7_75t_SL g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_323), .A2(n_454), .B(n_456), .C(n_458), .Y(n_453) );
INVx2_ASAP7_75t_L g366 ( .A(n_325), .Y(n_366) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI332xp33_ASAP7_75t_L g401 ( .A1(n_327), .A2(n_374), .A3(n_402), .B1(n_403), .B2(n_404), .B3(n_406), .C1(n_407), .C2(n_408), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B(n_335), .Y(n_329) );
AND2x2_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x4_ASAP7_75t_L g403 ( .A(n_331), .B(n_351), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_334), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_335), .B(n_339), .Y(n_338) );
NAND3xp33_ASAP7_75t_SL g337 ( .A(n_338), .B(n_343), .C(n_358), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_347), .B1(n_349), .B2(n_354), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g353 ( .A(n_345), .Y(n_353) );
AND2x2_ASAP7_75t_L g450 ( .A(n_345), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_350), .Y(n_369) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI31xp33_ASAP7_75t_L g377 ( .A1(n_354), .A2(n_378), .A3(n_380), .B(n_382), .Y(n_377) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g457 ( .A(n_355), .Y(n_457) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
BUFx2_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_365), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g443 ( .A(n_366), .Y(n_443) );
NOR3xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_383), .C(n_409), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_372), .B2(n_374), .C(n_377), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_370), .A2(n_390), .B(n_391), .Y(n_389) );
OR2x2_ASAP7_75t_L g465 ( .A(n_373), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_380), .A2(n_416), .B1(n_420), .B2(n_421), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g383 ( .A(n_384), .B(n_392), .C(n_401), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g462 ( .A(n_405), .B(n_463), .Y(n_462) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_415), .C(n_422), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g470 ( .A(n_419), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_421), .A2(n_441), .B1(n_444), .B2(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g442 ( .A(n_424), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_447), .C(n_464), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_453), .B1(n_459), .B2(n_462), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_670), .B1(n_688), .B2(n_690), .C(n_695), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_489), .B1(n_668), .B2(n_669), .Y(n_472) );
INVx1_ASAP7_75t_L g668 ( .A(n_473), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_483), .B2(n_484), .Y(n_473) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_481), .B2(n_482), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_476), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_477), .Y(n_482) );
INVx1_ASAP7_75t_L g480 ( .A(n_478), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g669 ( .A(n_489), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_489), .A2(n_669), .B1(n_701), .B2(n_702), .Y(n_700) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_572), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_516), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_502), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g514 ( .A(n_497), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_497), .B(n_501), .Y(n_527) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_498), .B(n_501), .Y(n_508) );
AND2x4_ASAP7_75t_L g531 ( .A(n_498), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
INVx1_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
AND2x2_ASAP7_75t_L g657 ( .A(n_498), .B(n_501), .Y(n_657) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g532 ( .A(n_501), .Y(n_532) );
INVx1_ASAP7_75t_L g537 ( .A(n_501), .Y(n_537) );
INVx1_ASAP7_75t_L g665 ( .A(n_501), .Y(n_665) );
AND2x2_ASAP7_75t_L g568 ( .A(n_502), .B(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g654 ( .A(n_502), .B(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g660 ( .A(n_502), .B(n_661), .Y(n_660) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
INVx1_ASAP7_75t_L g520 ( .A(n_505), .Y(n_520) );
INVx1_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx2_ASAP7_75t_SL g541 ( .A(n_507), .Y(n_541) );
INVx1_ASAP7_75t_L g554 ( .A(n_507), .Y(n_554) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g515 ( .A(n_509), .Y(n_515) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g663 ( .A(n_515), .B(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g666 ( .A(n_515), .B(n_667), .Y(n_666) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
BUFx2_ASAP7_75t_L g651 ( .A(n_521), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B1(n_528), .B2(n_529), .Y(n_522) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g546 ( .A(n_527), .Y(n_546) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_528), .A2(n_539), .B1(n_606), .B2(n_623), .C(n_624), .Y(n_622) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g549 ( .A(n_531), .Y(n_549) );
AND2x4_ASAP7_75t_L g570 ( .A(n_532), .B(n_571), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_539), .B2(n_540), .Y(n_533) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_537), .B(n_538), .Y(n_559) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_547), .B2(n_550), .Y(n_542) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g661 ( .A(n_549), .Y(n_661) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_553), .B1(n_555), .B2(n_556), .Y(n_551) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_555), .A2(n_601), .B1(n_615), .B2(n_617), .C(n_620), .Y(n_600) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx6_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x6_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g667 ( .A(n_570), .Y(n_667) );
AOI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_648), .B(n_652), .Y(n_572) );
NAND4xp25_ASAP7_75t_SL g573 ( .A(n_574), .B(n_600), .C(n_622), .D(n_631), .Y(n_573) );
AOI222xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_588), .B1(n_589), .B2(n_595), .C1(n_596), .C2(n_599), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
AND2x4_ASAP7_75t_L g591 ( .A(n_578), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g596 ( .A(n_578), .B(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g621 ( .A(n_578), .Y(n_621) );
AND2x4_ASAP7_75t_L g687 ( .A(n_578), .B(n_592), .Y(n_687) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g647 ( .A(n_581), .B(n_630), .Y(n_647) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g629 ( .A(n_582), .B(n_630), .Y(n_629) );
INVx6_ASAP7_75t_L g645 ( .A(n_583), .Y(n_645) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_L g598 ( .A(n_584), .Y(n_598) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g604 ( .A(n_585), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g619 ( .A(n_585), .B(n_587), .Y(n_619) );
INVx1_ASAP7_75t_L g594 ( .A(n_586), .Y(n_594) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g614 ( .A(n_587), .B(n_610), .Y(n_614) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx4_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g682 ( .A(n_593), .Y(n_682) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_595), .A2(n_663), .B(n_666), .Y(n_662) );
BUFx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_604), .Y(n_625) );
INVx1_ASAP7_75t_L g611 ( .A(n_605), .Y(n_611) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g623 ( .A(n_613), .Y(n_623) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g639 ( .A(n_614), .Y(n_639) );
AND2x4_ASAP7_75t_L g617 ( .A(n_615), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g620 ( .A(n_618), .B(n_621), .Y(n_620) );
BUFx4f_ASAP7_75t_L g626 ( .A(n_618), .Y(n_626) );
INVx1_ASAP7_75t_L g643 ( .A(n_618), .Y(n_643) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx3_ASAP7_75t_L g633 ( .A(n_625), .Y(n_633) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_SL g679 ( .A(n_629), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B1(n_635), .B2(n_640), .C(n_641), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
CKINVDCx20_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x6_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
OR2x4_ASAP7_75t_L g699 ( .A(n_673), .B(n_677), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_674), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g707 ( .A(n_674), .Y(n_707) );
INVx1_ASAP7_75t_L g694 ( .A(n_675), .Y(n_694) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI31xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .A3(n_683), .B(n_685), .Y(n_677) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx6_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_700), .B1(n_703), .B2(n_705), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx8_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_701), .Y(n_702) );
CKINVDCx14_ASAP7_75t_R g703 ( .A(n_704), .Y(n_703) );
BUFx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
endmodule