module fake_jpeg_16534_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_47),
.Y(n_72)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_31),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_20),
.Y(n_88)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_32),
.B1(n_16),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_25),
.B1(n_32),
.B2(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_30),
.Y(n_82)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_73),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_90),
.B1(n_94),
.B2(n_97),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_32),
.B1(n_24),
.B2(n_17),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_79),
.B1(n_98),
.B2(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_86),
.Y(n_114)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_35),
.C(n_40),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_70),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_31),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_88),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_20),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_71),
.B1(n_56),
.B2(n_64),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_41),
.B1(n_39),
.B2(n_33),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_41),
.A3(n_39),
.B1(n_22),
.B2(n_25),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_65),
.A3(n_27),
.B1(n_33),
.B2(n_53),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_59),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_65),
.B1(n_58),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_92),
.B1(n_91),
.B2(n_49),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_106),
.B1(n_115),
.B2(n_33),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_62),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_120),
.B(n_82),
.Y(n_136)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_122),
.B(n_123),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_97),
.B(n_84),
.Y(n_140)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_72),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_22),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_88),
.B1(n_76),
.B2(n_87),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_134),
.B1(n_141),
.B2(n_144),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_137),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_84),
.B1(n_78),
.B2(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_149),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_139),
.B(n_147),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_113),
.C(n_102),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_92),
.B1(n_90),
.B2(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_154),
.B1(n_122),
.B2(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_85),
.Y(n_148)
);

NOR2x1p5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_22),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_159),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_169),
.B1(n_107),
.B2(n_19),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_118),
.B(n_110),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_132),
.B(n_29),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_171),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_124),
.B1(n_102),
.B2(n_101),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_126),
.C(n_121),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_116),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_112),
.C(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_104),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_119),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_147),
.B1(n_150),
.B2(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_150),
.B1(n_101),
.B2(n_141),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_128),
.B1(n_146),
.B2(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_107),
.B1(n_130),
.B2(n_131),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_137),
.B(n_30),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_195),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_19),
.B(n_22),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_161),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_163),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_208),
.B1(n_166),
.B2(n_179),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_13),
.B1(n_11),
.B2(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_210),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_174),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_222),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_228),
.B1(n_233),
.B2(n_236),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_177),
.B(n_172),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_160),
.C(n_182),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_193),
.C(n_185),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_170),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_170),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_173),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_196),
.Y(n_256)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

OAI221xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.C(n_205),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_208),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_241),
.B(n_229),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_186),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_259),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_255),
.C(n_260),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_257),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_203),
.B(n_209),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_184),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_253),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_203),
.C(n_211),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_214),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_188),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_181),
.C(n_197),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_189),
.Y(n_261)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_189),
.Y(n_265)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_217),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_266),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_213),
.C(n_214),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_272),
.C(n_280),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_212),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_271),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_241),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_225),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_245),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_244),
.A2(n_225),
.B1(n_233),
.B2(n_234),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_234),
.B1(n_220),
.B2(n_210),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_260),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_251),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_272),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_280),
.Y(n_300)
);

OAI221xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_242),
.B1(n_239),
.B2(n_253),
.C(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_254),
.C(n_243),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_293),
.C(n_5),
.Y(n_308)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_288),
.B(n_295),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_11),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_4),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_2),
.B(n_4),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_292),
.B(n_297),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_269),
.B1(n_263),
.B2(n_264),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_4),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_10),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_4),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_302),
.B(n_304),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_310),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_268),
.B(n_263),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_303),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_291),
.B(n_5),
.CI(n_6),
.CON(n_305),
.SN(n_305)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_6),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_283),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_308),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_296),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_309)
);

BUFx4f_ASAP7_75t_SL g310 ( 
.A(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_317),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_292),
.B(n_286),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_314),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_293),
.B(n_283),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_7),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_8),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_8),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_9),
.C(n_10),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_300),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_329),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_308),
.B(n_304),
.Y(n_327)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_310),
.Y(n_329)
);

NAND4xp25_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_305),
.C(n_9),
.D(n_10),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_333),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_330),
.B(n_328),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_10),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_316),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_324),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_323),
.C(n_331),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_342),
.C(n_338),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_340),
.B(n_334),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_325),
.B(n_315),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_332),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_318),
.Y(n_347)
);


endmodule