module fake_jpeg_23973_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_18),
.C(n_29),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_52),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_20),
.B1(n_19),
.B2(n_31),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_28),
.B(n_32),
.Y(n_55)
);

OR2x4_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_62),
.B1(n_72),
.B2(n_74),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_24),
.B(n_23),
.Y(n_106)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_73),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_16),
.B1(n_31),
.B2(n_20),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_52),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_87),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_38),
.B1(n_37),
.B2(n_19),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_16),
.B1(n_31),
.B2(n_20),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_42),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_37),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_107),
.C(n_39),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_105),
.Y(n_122)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_57),
.B1(n_51),
.B2(n_24),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_104),
.B1(n_112),
.B2(n_22),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_21),
.B1(n_17),
.B2(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_18),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_19),
.B(n_29),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_73),
.C(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_39),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_77),
.B1(n_75),
.B2(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_121),
.B1(n_124),
.B2(n_136),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_133),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_125),
.B(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_77),
.B1(n_78),
.B2(n_65),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_60),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_137),
.C(n_139),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_68),
.B1(n_67),
.B2(n_61),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_58),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_106),
.B1(n_98),
.B2(n_104),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_79),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_21),
.B(n_24),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_71),
.B1(n_69),
.B2(n_66),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_39),
.B1(n_27),
.B2(n_25),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_96),
.B1(n_115),
.B2(n_32),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_92),
.C(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_144),
.B1(n_110),
.B2(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_92),
.B(n_22),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_32),
.B1(n_26),
.B2(n_83),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_148),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_116),
.B1(n_103),
.B2(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_153),
.B1(n_157),
.B2(n_163),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_108),
.B1(n_109),
.B2(n_91),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_108),
.C(n_110),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_151),
.C(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_101),
.B1(n_89),
.B2(n_97),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

OAI22x1_ASAP7_75t_SL g165 ( 
.A1(n_117),
.A2(n_32),
.B1(n_26),
.B2(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_171),
.B1(n_10),
.B2(n_14),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_139),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_26),
.CI(n_2),
.CON(n_167),
.SN(n_167)
);

MAJIxp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_174),
.C(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_8),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_175),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_8),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_138),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_9),
.C(n_13),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_9),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_118),
.B1(n_134),
.B2(n_124),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_172),
.A2(n_119),
.B(n_127),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_162),
.B1(n_164),
.B2(n_156),
.Y(n_212)
);

AOI21x1_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_118),
.B(n_135),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_178),
.B(n_1),
.CI(n_3),
.CON(n_226),
.SN(n_226)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_194),
.C(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_200),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_191),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_120),
.B(n_126),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_197),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_144),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_167),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_132),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_149),
.C(n_171),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_162),
.B1(n_176),
.B2(n_147),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_225),
.B1(n_192),
.B2(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_226),
.C(n_192),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_149),
.C(n_155),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_163),
.C(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_185),
.C(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_223),
.C(n_182),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_150),
.C(n_158),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_177),
.A2(n_167),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_178),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_198),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_238),
.B1(n_216),
.B2(n_213),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_202),
.C(n_203),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_215),
.C(n_214),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_196),
.B1(n_197),
.B2(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_189),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_186),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_182),
.C(n_181),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_221),
.C(n_181),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_221),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_243),
.B(n_206),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_249),
.B(n_234),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_206),
.B(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_223),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_258),
.C(n_259),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_211),
.B1(n_207),
.B2(n_210),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_235),
.B1(n_226),
.B2(n_180),
.Y(n_270)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.Y(n_281)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_268),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_250),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_232),
.B1(n_230),
.B2(n_191),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_226),
.B1(n_180),
.B2(n_12),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_255),
.A3(n_257),
.B1(n_245),
.B2(n_205),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_247),
.B(n_253),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_267),
.B(n_261),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_262),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_248),
.C(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_277),
.C(n_4),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_248),
.C(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_279),
.A2(n_269),
.B1(n_11),
.B2(n_10),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_283),
.B(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_286),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_11),
.B(n_12),
.Y(n_285)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_13),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_280),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_288),
.B(n_274),
.Y(n_295)
);

OAI321xp33_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_296),
.A3(n_297),
.B1(n_294),
.B2(n_293),
.C(n_14),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_277),
.C(n_13),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_5),
.C(n_6),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_5),
.C(n_6),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_300),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_5),
.Y(n_302)
);


endmodule