module fake_jpeg_27849_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_22),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_20),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_14),
.B(n_26),
.C(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_16),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_13),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_18),
.B1(n_33),
.B2(n_17),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_54),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_29),
.C(n_28),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_32),
.C(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_33),
.B1(n_12),
.B2(n_22),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_59),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_29),
.B1(n_21),
.B2(n_23),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_36),
.B1(n_39),
.B2(n_15),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_22),
.B(n_12),
.C(n_14),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_78),
.B(n_13),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_66),
.B1(n_52),
.B2(n_48),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_15),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_46),
.C(n_45),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_59),
.C(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_58),
.B1(n_60),
.B2(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_86),
.C(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_51),
.Y(n_88)
);

AOI22x1_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_44),
.B1(n_31),
.B2(n_32),
.Y(n_89)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_78),
.A3(n_72),
.B1(n_66),
.B2(n_68),
.C(n_45),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_64),
.B1(n_71),
.B2(n_69),
.C(n_15),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_46),
.C(n_61),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_71),
.C(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_19),
.B1(n_13),
.B2(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_88),
.C(n_23),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_24),
.B(n_25),
.C(n_45),
.D(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_80),
.B1(n_91),
.B2(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_107),
.B1(n_93),
.B2(n_101),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.C(n_99),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_86),
.B(n_82),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_111),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_116),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_103),
.C(n_107),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_118),
.B(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_19),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_25),
.B1(n_6),
.B2(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_6),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_6),
.B(n_9),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_108),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_110),
.C(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_123),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_126),
.A3(n_127),
.B1(n_123),
.B2(n_5),
.C1(n_3),
.C2(n_4),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_114),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_5),
.C(n_8),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_10),
.C(n_0),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_0),
.A3(n_1),
.B1(n_10),
.B2(n_112),
.C1(n_115),
.C2(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);


endmodule