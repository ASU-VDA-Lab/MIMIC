module fake_jpeg_32199_n_527 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_20),
.A2(n_17),
.B1(n_9),
.B2(n_3),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_52),
.A2(n_45),
.B1(n_51),
.B2(n_46),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_82),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_23),
.B(n_10),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_64),
.B(n_102),
.Y(n_134)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_29),
.B(n_31),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_87),
.Y(n_138)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_36),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_10),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_29),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_101),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_100),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_31),
.B(n_11),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_105),
.Y(n_144)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_30),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_50),
.B1(n_41),
.B2(n_28),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_114),
.A2(n_121),
.B1(n_135),
.B2(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_60),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_141),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_52),
.A2(n_35),
.B1(n_34),
.B2(n_47),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_120),
.A2(n_131),
.B1(n_133),
.B2(n_80),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_50),
.B1(n_28),
.B2(n_32),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_47),
.B1(n_35),
.B2(n_50),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_59),
.A2(n_32),
.B1(n_49),
.B2(n_43),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_87),
.B(n_43),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_84),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_143),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_68),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_77),
.A2(n_45),
.B1(n_51),
.B2(n_46),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_153),
.B1(n_156),
.B2(n_162),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_49),
.B1(n_37),
.B2(n_36),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_44),
.B1(n_37),
.B2(n_30),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_75),
.A2(n_12),
.B1(n_17),
.B2(n_4),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_79),
.A2(n_44),
.B1(n_12),
.B2(n_4),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_99),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_168),
.B(n_181),
.Y(n_228)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_171),
.B(n_173),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_44),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_110),
.B(n_13),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_174),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_74),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_175),
.B(n_176),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_19),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx6_ASAP7_75t_SL g270 ( 
.A(n_180),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_97),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_184),
.Y(n_268)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_118),
.A2(n_53),
.B1(n_88),
.B2(n_85),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_189),
.A2(n_192),
.B1(n_210),
.B2(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_98),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_223),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_109),
.B(n_73),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_196),
.B(n_212),
.C(n_216),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_71),
.B1(n_70),
.B2(n_69),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_167),
.B1(n_148),
.B2(n_140),
.Y(n_237)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_106),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_200),
.B(n_209),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_204),
.B1(n_221),
.B2(n_222),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_203),
.Y(n_247)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_205),
.B(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_207),
.B(n_208),
.Y(n_272)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_118),
.A2(n_53),
.B1(n_62),
.B2(n_61),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_137),
.A2(n_57),
.B1(n_55),
.B2(n_54),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_215),
.B(n_218),
.Y(n_269)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_117),
.B(n_19),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_127),
.A2(n_11),
.B1(n_15),
.B2(n_4),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_165),
.B1(n_164),
.B2(n_158),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_117),
.B(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_156),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_113),
.B1(n_132),
.B2(n_162),
.Y(n_235)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_226),
.Y(n_260)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_112),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_135),
.B1(n_114),
.B2(n_167),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_234),
.A2(n_239),
.B(n_27),
.C(n_8),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_235),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_237),
.A2(n_246),
.B1(n_204),
.B2(n_193),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_148),
.B1(n_140),
.B2(n_158),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_172),
.A2(n_147),
.B(n_129),
.C(n_132),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_241),
.A2(n_0),
.B(n_1),
.Y(n_307)
);

AOI222xp33_ASAP7_75t_L g242 ( 
.A1(n_172),
.A2(n_179),
.B1(n_168),
.B2(n_211),
.C1(n_190),
.C2(n_181),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_242),
.A2(n_203),
.B(n_186),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_243),
.A2(n_245),
.B1(n_27),
.B2(n_8),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_177),
.A2(n_172),
.B1(n_197),
.B2(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_177),
.A2(n_165),
.B1(n_164),
.B2(n_154),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_13),
.B(n_17),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_250),
.A2(n_227),
.B(n_234),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_183),
.B(n_154),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_151),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_199),
.B(n_0),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_27),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_191),
.B(n_151),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_184),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_27),
.C(n_19),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_208),
.C(n_215),
.Y(n_278)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_281),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_289),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_226),
.C(n_195),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_284),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_225),
.C(n_223),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_185),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_287),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_286),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_178),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_288),
.B(n_297),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_251),
.B(n_188),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_291),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_267),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_264),
.B1(n_248),
.B2(n_259),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_294),
.B1(n_248),
.B2(n_253),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_270),
.A2(n_169),
.B1(n_207),
.B2(n_201),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_249),
.Y(n_295)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_19),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_298),
.A2(n_305),
.B1(n_239),
.B2(n_243),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_27),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_184),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_310),
.Y(n_328)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_227),
.B(n_170),
.C(n_184),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_302),
.B(n_313),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_265),
.C(n_230),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_303),
.B(n_252),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_304),
.A2(n_306),
.B1(n_232),
.B2(n_252),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_8),
.B1(n_15),
.B2(n_4),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_311),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_242),
.A2(n_1),
.B(n_5),
.C(n_7),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_308),
.A2(n_229),
.B(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_227),
.B(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_5),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_316),
.A2(n_329),
.B(n_302),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_274),
.B1(n_277),
.B2(n_290),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_318),
.A2(n_323),
.B1(n_349),
.B2(n_305),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_237),
.B1(n_246),
.B2(n_235),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_313),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_325),
.A2(n_333),
.B1(n_339),
.B2(n_256),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_330),
.A2(n_248),
.B1(n_258),
.B2(n_301),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_235),
.B1(n_241),
.B2(n_269),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_338),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_312),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_289),
.A2(n_235),
.B1(n_269),
.B2(n_268),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_341),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_275),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_275),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_310),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_307),
.A2(n_269),
.B(n_229),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_348),
.A2(n_308),
.B(n_305),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_291),
.A2(n_268),
.B1(n_230),
.B2(n_258),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_314),
.B(n_279),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_352),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_353),
.A2(n_371),
.B1(n_380),
.B2(n_382),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_281),
.C(n_278),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_373),
.C(n_346),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_358),
.A2(n_359),
.B1(n_366),
.B2(n_369),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_305),
.B1(n_308),
.B2(n_286),
.Y(n_359)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_361),
.B(n_368),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_296),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_374),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_284),
.Y(n_363)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_364),
.B(n_315),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_319),
.A2(n_308),
.B(n_305),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_365),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_343),
.A2(n_308),
.B(n_309),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_367),
.A2(n_375),
.B(n_354),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_314),
.B(n_283),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_318),
.A2(n_311),
.B1(n_295),
.B2(n_238),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_236),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_370),
.Y(n_409)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_238),
.B1(n_255),
.B2(n_236),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_372),
.A2(n_379),
.B1(n_380),
.B2(n_382),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_257),
.C(n_233),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_257),
.B(n_233),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_343),
.A2(n_249),
.B(n_256),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_349),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_376),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_326),
.B1(n_317),
.B2(n_332),
.Y(n_390)
);

AOI22x1_ASAP7_75t_L g378 ( 
.A1(n_325),
.A2(n_333),
.B1(n_327),
.B2(n_332),
.Y(n_378)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_378),
.A2(n_339),
.B(n_327),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_330),
.A2(n_255),
.B1(n_7),
.B2(n_11),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_346),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_328),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_321),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_387),
.B(n_391),
.C(n_395),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_401),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_390),
.A2(n_398),
.B1(n_408),
.B2(n_411),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_328),
.C(n_326),
.Y(n_395)
);

OAI22x1_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_348),
.B1(n_337),
.B2(n_324),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_396),
.A2(n_355),
.B(n_352),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_317),
.C(n_344),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_402),
.C(n_403),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_377),
.A2(n_320),
.B1(n_344),
.B2(n_338),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_400),
.A2(n_353),
.B(n_365),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_320),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_315),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_412),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_334),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_407),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_334),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_322),
.B1(n_345),
.B2(n_14),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_378),
.A2(n_354),
.B1(n_355),
.B2(n_358),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_414),
.A2(n_421),
.B(n_428),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_416),
.B(n_402),
.Y(n_447)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_411),
.A2(n_392),
.B1(n_393),
.B2(n_390),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_418),
.A2(n_389),
.B1(n_399),
.B2(n_378),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_384),
.Y(n_419)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_422),
.Y(n_445)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_410),
.B(n_370),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_368),
.B1(n_397),
.B2(n_372),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_360),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_426),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_388),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_429),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_396),
.A2(n_364),
.B(n_398),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_371),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_431),
.Y(n_458)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_433),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_351),
.Y(n_433)
);

INVx13_ASAP7_75t_L g435 ( 
.A(n_388),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_435),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_369),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_436),
.A2(n_385),
.B(n_375),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_374),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_5),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_440),
.A2(n_457),
.B1(n_422),
.B2(n_438),
.Y(n_468)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_387),
.C(n_437),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_449),
.C(n_454),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_447),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_405),
.C(n_395),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_414),
.A2(n_367),
.B(n_391),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_450),
.A2(n_428),
.B(n_432),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_356),
.C(n_345),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_431),
.A2(n_379),
.B1(n_356),
.B2(n_14),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_457),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_419),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_413),
.A2(n_5),
.B1(n_7),
.B2(n_17),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_424),
.C(n_430),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_424),
.C(n_430),
.Y(n_473)
);

XOR2x1_ASAP7_75t_SL g460 ( 
.A(n_441),
.B(n_416),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_460),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_451),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_465),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_421),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_433),
.Y(n_466)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_468),
.A2(n_413),
.B1(n_436),
.B2(n_462),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_470),
.A2(n_450),
.B(n_446),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_437),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_473),
.C(n_443),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_454),
.B(n_423),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_474),
.A2(n_476),
.B1(n_427),
.B2(n_445),
.Y(n_489)
);

OA22x2_ASAP7_75t_L g475 ( 
.A1(n_440),
.A2(n_435),
.B1(n_426),
.B2(n_418),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_448),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_470),
.Y(n_495)
);

NOR3xp33_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_420),
.C(n_425),
.Y(n_478)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_489),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_435),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_449),
.C(n_458),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_488),
.C(n_471),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_485),
.A2(n_415),
.B1(n_466),
.B2(n_475),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_465),
.A2(n_445),
.B(n_453),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_472),
.B(n_444),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_429),
.C(n_452),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_463),
.A2(n_415),
.B1(n_427),
.B2(n_452),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_468),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_493),
.B(n_500),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_473),
.C(n_475),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_501),
.C(n_503),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_496),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_480),
.B1(n_486),
.B2(n_477),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_499),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_482),
.A2(n_455),
.B1(n_475),
.B2(n_427),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_447),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_480),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_464),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_508),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_R g509 ( 
.A(n_497),
.B(n_483),
.Y(n_509)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_509),
.A2(n_511),
.B(n_488),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_492),
.A2(n_481),
.B(n_491),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_494),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_513),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_506),
.A2(n_487),
.B1(n_495),
.B2(n_503),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_514),
.A2(n_510),
.B(n_502),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g515 ( 
.A(n_504),
.B(n_493),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_515),
.B(n_504),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_518),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_516),
.Y(n_520)
);

OAI311xp33_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_508),
.A3(n_500),
.B1(n_506),
.C1(n_485),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_439),
.C(n_501),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_521),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_439),
.C(n_417),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_417),
.B(n_510),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_417),
.Y(n_527)
);


endmodule