module fake_jpeg_18866_n_60 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_55;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

AO22x1_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_38),
.B1(n_42),
.B2(n_29),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_34),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_23),
.C(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_38),
.B(n_31),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_42),
.B(n_43),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_45),
.B(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_48),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.C(n_34),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.C(n_35),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_22),
.B(n_27),
.Y(n_58)
);

OAI21x1_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_20),
.B(n_26),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_33),
.Y(n_60)
);


endmodule