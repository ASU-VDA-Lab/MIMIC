module fake_aes_11532_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_7), .B(n_3), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_4), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_0), .B(n_2), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_14), .B(n_0), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_14), .B(n_0), .Y(n_21) );
OA21x2_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_15), .B(n_17), .Y(n_22) );
OAI22xp33_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_16), .B1(n_12), .B2(n_15), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_18), .B1(n_21), .B2(n_23), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_21), .B1(n_22), .B2(n_17), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_17), .B1(n_16), .B2(n_22), .Y(n_29) );
AOI221xp5_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_28), .B1(n_12), .B2(n_15), .C(n_13), .Y(n_30) );
AOI322xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_17), .A3(n_13), .B1(n_1), .B2(n_6), .C1(n_7), .C2(n_5), .Y(n_31) );
AOI211xp5_ASAP7_75t_L g32 ( .A1(n_28), .A2(n_17), .B(n_13), .C(n_8), .Y(n_32) );
OAI311xp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_13), .A3(n_5), .B1(n_9), .C1(n_10), .Y(n_33) );
AND4x1_ASAP7_75t_L g34 ( .A(n_32), .B(n_4), .C(n_9), .D(n_10), .Y(n_34) );
OAI21xp5_ASAP7_75t_L g35 ( .A1(n_30), .A2(n_17), .B(n_13), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_34), .Y(n_37) );
AOI22xp33_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_34), .B1(n_33), .B2(n_31), .Y(n_38) );
OAI22xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_11), .B1(n_36), .B2(n_37), .Y(n_39) );
endmodule