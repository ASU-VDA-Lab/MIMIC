module fake_netlist_5_1528_n_1844 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1844);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1844;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_1014;
wire n_279;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_90),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_94),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_163),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_83),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_21),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_89),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_98),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_2),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_103),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_30),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_77),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_48),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_25),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_47),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_20),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_40),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_147),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_6),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_64),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_109),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_82),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_13),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_80),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_63),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_86),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_157),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_9),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

INVx4_ASAP7_75t_R g237 ( 
.A(n_102),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_160),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_20),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_33),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_78),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_49),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_22),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_180),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_61),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_114),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_177),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_58),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_154),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_188),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_156),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_87),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_120),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_124),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_108),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_182),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_22),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_171),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_126),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_16),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_40),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_74),
.Y(n_271)
);

CKINVDCx11_ASAP7_75t_R g272 ( 
.A(n_99),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_122),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_41),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_84),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_139),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_165),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_54),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_178),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_121),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_31),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_153),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_116),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_73),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_113),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_52),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_88),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_179),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_60),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_16),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_130),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_175),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_14),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_50),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_41),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_70),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_149),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_134),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_162),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_173),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_161),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_30),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_95),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_128),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_185),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_164),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_110),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_15),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_101),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_38),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_28),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_12),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_79),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_92),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_21),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_81),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_42),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_46),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_117),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_24),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_184),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_174),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_42),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_36),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_123),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_66),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_62),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_76),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_51),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_31),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_118),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_146),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_35),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_13),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_71),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_4),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_7),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_138),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_59),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_50),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_119),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_45),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_29),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_4),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_1),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_141),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_43),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_93),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_125),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_9),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_44),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_29),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_148),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_38),
.Y(n_357)
);

BUFx8_ASAP7_75t_SL g358 ( 
.A(n_45),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_53),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_112),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_72),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_11),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_26),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_176),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_28),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_158),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_129),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_49),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_137),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_34),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_69),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_10),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_18),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_2),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_19),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_91),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_65),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_7),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_209),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_198),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_210),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_216),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_234),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_239),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_243),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_244),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_245),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_254),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_278),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_358),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_310),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_286),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_222),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_235),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_198),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_302),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_232),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_258),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_312),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_301),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_305),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_317),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_194),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_272),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_207),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_240),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_246),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_196),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_242),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_203),
.Y(n_420)
);

INVxp33_ASAP7_75t_SL g421 ( 
.A(n_203),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_270),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_206),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_196),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_207),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_241),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_241),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_248),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_252),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_207),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_233),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_309),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_324),
.Y(n_440)
);

INVxp33_ASAP7_75t_SL g441 ( 
.A(n_206),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_261),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_261),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_266),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_282),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_283),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_283),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_270),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_338),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_201),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_270),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_205),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_217),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_269),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_274),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_211),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_227),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_211),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_293),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_293),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_192),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_290),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_192),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_219),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_294),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_219),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_271),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_271),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_275),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_213),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_275),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_295),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_236),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_432),
.A2(n_331),
.B(n_280),
.Y(n_476)
);

AND3x2_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_345),
.C(n_377),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_396),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_401),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_437),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_413),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_413),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_417),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_438),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_416),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_464),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_364),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_431),
.B(n_334),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_465),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_467),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_468),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_423),
.A2(n_320),
.B1(n_260),
.B2(n_375),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_470),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_R g512 ( 
.A(n_397),
.B(n_190),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_416),
.B(n_280),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_404),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_394),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_472),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_381),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_379),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_379),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_380),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_381),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_405),
.B(n_343),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_385),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_408),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_380),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_412),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_334),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_385),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_454),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_388),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_400),
.B(n_331),
.Y(n_534)
);

NOR2x1_ASAP7_75t_L g535 ( 
.A(n_458),
.B(n_377),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_388),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_434),
.B(n_334),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_389),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_415),
.B(n_251),
.Y(n_540)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_407),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_439),
.B(n_264),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_390),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_390),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_391),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_391),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_453),
.B(n_193),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_392),
.Y(n_550)
);

BUFx12f_ASAP7_75t_L g551 ( 
.A(n_397),
.Y(n_551)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_545),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_490),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_545),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_482),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_483),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_548),
.B(n_498),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_545),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_489),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_483),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_490),
.B(n_382),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_479),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_524),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_420),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_534),
.A2(n_445),
.B1(n_446),
.B2(n_443),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_540),
.A2(n_448),
.B1(n_450),
.B2(n_447),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_545),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_481),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_532),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_513),
.B(n_414),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_527),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_476),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

CKINVDCx6p67_ASAP7_75t_R g578 ( 
.A(n_551),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_476),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_478),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_530),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_524),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_527),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_480),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_515),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_542),
.B(n_421),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_476),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

BUFx6f_ASAP7_75t_SL g589 ( 
.A(n_519),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_530),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_527),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_527),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_500),
.A2(n_457),
.B1(n_441),
.B2(n_428),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_530),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_494),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_530),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_543),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_543),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_543),
.B(n_414),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_494),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_543),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_500),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_512),
.A2(n_357),
.B1(n_212),
.B2(n_214),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_526),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_543),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_529),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_482),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_494),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_535),
.A2(n_496),
.B(n_493),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_529),
.B(n_537),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_552),
.B(n_419),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_549),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_494),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_475),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_494),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_549),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_537),
.A2(n_398),
.B1(n_471),
.B2(n_459),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_495),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_535),
.B(n_473),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_495),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_482),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_435),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_541),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_495),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_501),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_501),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_541),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_497),
.B(n_436),
.C(n_435),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_550),
.Y(n_640)
);

AND3x2_ASAP7_75t_L g641 ( 
.A(n_514),
.B(n_452),
.C(n_393),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_550),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_482),
.Y(n_644)
);

CKINVDCx6p67_ASAP7_75t_R g645 ( 
.A(n_551),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_510),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_550),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_519),
.A2(n_386),
.B1(n_383),
.B2(n_384),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_493),
.B(n_460),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_523),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_514),
.B(n_436),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_516),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_523),
.A2(n_387),
.B1(n_422),
.B2(n_418),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_525),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_484),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_509),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_509),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_503),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_511),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_503),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_525),
.Y(n_661)
);

BUFx8_ASAP7_75t_SL g662 ( 
.A(n_528),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_503),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

BUFx8_ASAP7_75t_SL g665 ( 
.A(n_516),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_475),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_541),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_541),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_484),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_505),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_531),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_503),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_SL g673 ( 
.A(n_533),
.B(n_444),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_547),
.B(n_267),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_503),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_541),
.B(n_268),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_496),
.B(n_444),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_477),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_533),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_484),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_503),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_536),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_536),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_538),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_538),
.B(n_455),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_475),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_539),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_504),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_504),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_504),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_504),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_539),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_547),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_544),
.B(n_456),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_544),
.B(n_456),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_499),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_546),
.A2(n_424),
.B1(n_425),
.B2(n_427),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_487),
.B(n_463),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_617),
.B(n_463),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_586),
.A2(n_473),
.B1(n_466),
.B2(n_289),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_683),
.B(n_466),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_650),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_572),
.A2(n_485),
.B(n_484),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_617),
.B(n_522),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_677),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_685),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_607),
.B(n_612),
.Y(n_708)
);

OAI221xp5_ASAP7_75t_L g709 ( 
.A1(n_568),
.A2(n_356),
.B1(n_349),
.B2(n_238),
.C(n_546),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_685),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_612),
.B(n_522),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_R g712 ( 
.A(n_561),
.B(n_190),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_684),
.B(n_207),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_654),
.B(n_522),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_604),
.B(n_247),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_654),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_572),
.A2(n_207),
.B1(n_215),
.B2(n_344),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_638),
.B(n_499),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_661),
.B(n_487),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_652),
.Y(n_720)
);

NAND2x1_ASAP7_75t_L g721 ( 
.A(n_572),
.B(n_487),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_559),
.B(n_411),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_664),
.B(n_487),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_566),
.B(n_429),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_553),
.B(n_215),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_671),
.Y(n_726)
);

INVx8_ASAP7_75t_L g727 ( 
.A(n_589),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_553),
.B(n_215),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_671),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_666),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_597),
.B(n_460),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_626),
.A2(n_679),
.B(n_687),
.C(n_682),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_679),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_562),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_682),
.B(n_504),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_555),
.B(n_215),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_687),
.B(n_504),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_673),
.B(n_313),
.C(n_311),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_692),
.B(n_507),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_692),
.B(n_507),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_698),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_SL g742 ( 
.A(n_589),
.B(n_213),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_646),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_693),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_574),
.B(n_507),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_696),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_576),
.A2(n_215),
.B1(n_344),
.B2(n_276),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_608),
.A2(n_430),
.B(n_399),
.C(n_402),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_696),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_576),
.B(n_507),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_576),
.B(n_507),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_555),
.B(n_344),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_578),
.B(n_191),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_579),
.B(n_507),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_624),
.B(n_336),
.C(n_326),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_649),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_579),
.B(n_511),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_579),
.B(n_511),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_589),
.B(n_214),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_564),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_587),
.B(n_502),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_563),
.B(n_461),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_649),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_676),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_587),
.B(n_502),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_560),
.B(n_344),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_560),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_570),
.B(n_344),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_570),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_618),
.B(n_629),
.Y(n_770)
);

AOI221x1_ASAP7_75t_L g771 ( 
.A1(n_581),
.A2(n_325),
.B1(n_277),
.B2(n_316),
.C(n_352),
.Y(n_771)
);

OAI221xp5_ASAP7_75t_L g772 ( 
.A1(n_569),
.A2(n_342),
.B1(n_296),
.B2(n_291),
.C(n_288),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_694),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_L g774 ( 
.A(n_631),
.B(n_506),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_631),
.B(n_506),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_587),
.B(n_508),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_616),
.B(n_298),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_554),
.B(n_508),
.Y(n_778)
);

AO221x1_ASAP7_75t_L g779 ( 
.A1(n_670),
.A2(n_304),
.B1(n_307),
.B2(n_461),
.C(n_399),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_554),
.B(n_249),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_636),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_636),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_695),
.B(n_191),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_616),
.B(n_667),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_667),
.B(n_250),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_567),
.B(n_195),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_621),
.B(n_517),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_573),
.B(n_253),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_L g789 ( 
.A(n_651),
.B(n_403),
.C(n_402),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_582),
.B(n_403),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_608),
.B(n_195),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_562),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_589),
.B(n_197),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_686),
.B(n_517),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_578),
.B(n_197),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_668),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_581),
.B(n_255),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_564),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_565),
.Y(n_799)
);

AND2x4_ASAP7_75t_SL g800 ( 
.A(n_645),
.B(n_281),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_676),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_565),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_674),
.Y(n_803)
);

O2A1O1Ixp5_ASAP7_75t_L g804 ( 
.A1(n_674),
.A2(n_518),
.B(n_521),
.C(n_520),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_665),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_666),
.B(n_520),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_577),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_580),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_565),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_571),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_571),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_571),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_613),
.A2(n_359),
.B1(n_225),
.B2(n_340),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_678),
.B(n_676),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_666),
.B(n_520),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_613),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_562),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_590),
.B(n_256),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_676),
.B(n_199),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_645),
.B(n_281),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_619),
.Y(n_821)
);

OAI221xp5_ASAP7_75t_L g822 ( 
.A1(n_648),
.A2(n_406),
.B1(n_410),
.B2(n_409),
.C(n_488),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_588),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_619),
.B(n_521),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_588),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_590),
.B(n_257),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_588),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_641),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_623),
.B(n_521),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_623),
.B(n_484),
.Y(n_830)
);

INVxp33_ASAP7_75t_L g831 ( 
.A(n_662),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_640),
.Y(n_832)
);

INVx8_ASAP7_75t_L g833 ( 
.A(n_676),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_625),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_634),
.B(n_492),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_584),
.B(n_406),
.C(n_409),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_585),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_595),
.B(n_259),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_634),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_640),
.B(n_484),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_609),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_643),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_595),
.B(n_262),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_643),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_647),
.B(n_485),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_653),
.B(n_337),
.C(n_339),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_697),
.B(n_281),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_647),
.B(n_199),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_625),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_627),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_634),
.B(n_350),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_808),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_706),
.B(n_642),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_767),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_769),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_705),
.B(n_627),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_748),
.A2(n_659),
.B(n_635),
.C(n_637),
.Y(n_857)
);

AND2x6_ASAP7_75t_L g858 ( 
.A(n_814),
.B(n_591),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_786),
.B(n_598),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_SL g860 ( 
.A(n_701),
.B(n_225),
.C(n_220),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_827),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_722),
.B(n_350),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_741),
.B(n_632),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_702),
.B(n_200),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_790),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_707),
.B(n_200),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_699),
.Y(n_867)
);

AND2x6_ASAP7_75t_L g868 ( 
.A(n_814),
.B(n_591),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_827),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_703),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_825),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_825),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_716),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_727),
.B(n_837),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_722),
.B(n_350),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_717),
.B(n_632),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_786),
.B(n_598),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_825),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_730),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_717),
.B(n_633),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_727),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_726),
.B(n_599),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_729),
.B(n_599),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_803),
.A2(n_601),
.B1(n_602),
.B2(n_603),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_712),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_841),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_733),
.B(n_601),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_756),
.B(n_410),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_763),
.B(n_486),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_770),
.A2(n_610),
.B1(n_606),
.B2(n_603),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_796),
.B(n_486),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_744),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_746),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_749),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_750),
.A2(n_606),
.B(n_602),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_710),
.B(n_202),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_730),
.Y(n_897)
);

OR2x4_ASAP7_75t_L g898 ( 
.A(n_791),
.B(n_488),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_743),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_773),
.B(n_202),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_727),
.Y(n_901)
);

CKINVDCx11_ASAP7_75t_R g902 ( 
.A(n_796),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_761),
.B(n_633),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_765),
.B(n_635),
.Y(n_904)
);

AND2x6_ASAP7_75t_SL g905 ( 
.A(n_791),
.B(n_491),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_825),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_708),
.B(n_204),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_700),
.B(n_204),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_720),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_762),
.B(n_208),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_839),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_709),
.A2(n_610),
.B1(n_656),
.B2(n_637),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_776),
.B(n_639),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_724),
.B(n_218),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_712),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_781),
.B(n_491),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_760),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_731),
.B(n_492),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_781),
.B(n_575),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_760),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_847),
.B(n_220),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_851),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_800),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_747),
.B(n_639),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_747),
.B(n_656),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_782),
.B(n_630),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_783),
.B(n_218),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_757),
.B(n_657),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_828),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_805),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_839),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_SL g932 ( 
.A1(n_813),
.A2(n_340),
.B1(n_346),
.B2(n_373),
.Y(n_932)
);

AND3x1_ASAP7_75t_L g933 ( 
.A(n_748),
.B(n_347),
.C(n_346),
.Y(n_933)
);

INVx6_ASAP7_75t_L g934 ( 
.A(n_820),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_732),
.A2(n_583),
.B(n_575),
.C(n_689),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_798),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_755),
.B(n_347),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_783),
.B(n_221),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_742),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_839),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_800),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_839),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_758),
.B(n_657),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_793),
.B(n_221),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_745),
.B(n_659),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_842),
.B(n_583),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_782),
.B(n_591),
.Y(n_947)
);

BUFx5_ASAP7_75t_L g948 ( 
.A(n_811),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_718),
.B(n_223),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_711),
.B(n_592),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_779),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_835),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_807),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_816),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_751),
.B(n_592),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_738),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_778),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_713),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_754),
.B(n_592),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_833),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_836),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_813),
.B(n_353),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_822),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_798),
.B(n_594),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_821),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_799),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_833),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_832),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_819),
.A2(n_691),
.B(n_690),
.C(n_689),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_823),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_759),
.B(n_285),
.C(n_376),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_799),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_785),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_713),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_833),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_823),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_846),
.B(n_353),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_785),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_835),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_721),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_802),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_802),
.B(n_594),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_809),
.B(n_594),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_753),
.B(n_224),
.Y(n_984)
);

OA22x2_ASAP7_75t_L g985 ( 
.A1(n_771),
.A2(n_355),
.B1(n_359),
.B2(n_373),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_788),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_784),
.A2(n_704),
.B(n_806),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_784),
.A2(n_630),
.B(n_658),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_844),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_818),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_809),
.B(n_596),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_789),
.B(n_355),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_818),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_795),
.Y(n_994)
);

OR2x6_ASAP7_75t_L g995 ( 
.A(n_764),
.B(n_596),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_810),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_787),
.B(n_596),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_838),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_794),
.B(n_600),
.Y(n_999)
);

BUFx4f_ASAP7_75t_SL g1000 ( 
.A(n_838),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_764),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_714),
.B(n_600),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_834),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_849),
.B(n_600),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_L g1005 ( 
.A(n_772),
.B(n_226),
.C(n_376),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_812),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_605),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_734),
.B(n_605),
.Y(n_1008)
);

INVx3_ASAP7_75t_SL g1009 ( 
.A(n_843),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_774),
.B(n_226),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_SL g1011 ( 
.A(n_831),
.B(n_363),
.C(n_372),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_775),
.B(n_228),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_792),
.B(n_605),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_801),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_719),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_801),
.B(n_691),
.Y(n_1016)
);

INVx6_ASAP7_75t_L g1017 ( 
.A(n_780),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_988),
.A2(n_815),
.B(n_658),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_927),
.A2(n_848),
.B1(n_777),
.B2(n_843),
.Y(n_1019)
);

INVx6_ASAP7_75t_L g1020 ( 
.A(n_886),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_957),
.B(n_777),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_938),
.A2(n_804),
.B(n_723),
.C(n_739),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_957),
.B(n_735),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_865),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_993),
.B(n_998),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_990),
.A2(n_737),
.B(n_740),
.C(n_715),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_967),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_SL g1028 ( 
.A1(n_939),
.A2(n_932),
.B1(n_930),
.B2(n_994),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_918),
.B(n_824),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_984),
.B(n_914),
.C(n_961),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_909),
.B(n_817),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_895),
.A2(n_829),
.B(n_840),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_859),
.B(n_830),
.Y(n_1033)
);

AND2x6_ASAP7_75t_L g1034 ( 
.A(n_967),
.B(n_615),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_898),
.B(n_797),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_826),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_860),
.A2(n_768),
.B(n_766),
.C(n_752),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_877),
.B(n_845),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_853),
.B(n_556),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_981),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_987),
.A2(n_660),
.B(n_630),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_921),
.B(n_725),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_867),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_922),
.B(n_973),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_SL g1045 ( 
.A1(n_971),
.A2(n_622),
.B(n_620),
.C(n_663),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_970),
.A2(n_658),
.B(n_660),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_902),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_929),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_870),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_899),
.B(n_728),
.Y(n_1050)
);

AO32x2_ASAP7_75t_L g1051 ( 
.A1(n_951),
.A2(n_681),
.A3(n_660),
.B1(n_658),
.B2(n_736),
.Y(n_1051)
);

AO32x2_ASAP7_75t_L g1052 ( 
.A1(n_958),
.A2(n_681),
.A3(n_766),
.B1(n_752),
.B2(n_736),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_863),
.B(n_873),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_945),
.A2(n_681),
.B(n_644),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_863),
.B(n_556),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_945),
.A2(n_681),
.B(n_644),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_978),
.B(n_363),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_852),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_891),
.B(n_229),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_891),
.B(n_229),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_967),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_874),
.B(n_768),
.Y(n_1062)
);

AND2x6_ASAP7_75t_L g1063 ( 
.A(n_975),
.B(n_615),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1000),
.B(n_230),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_974),
.A2(n_361),
.B1(n_366),
.B2(n_369),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_903),
.A2(n_669),
.B(n_611),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1017),
.A2(n_231),
.B1(n_371),
.B2(n_369),
.Y(n_1067)
);

BUFx4_ASAP7_75t_SL g1068 ( 
.A(n_874),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_962),
.A2(n_372),
.B(n_284),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_904),
.A2(n_611),
.B(n_644),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1001),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_872),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_872),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_910),
.A2(n_688),
.B(n_620),
.C(n_675),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_861),
.B(n_230),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_904),
.A2(n_669),
.B(n_611),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_892),
.B(n_593),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_986),
.A2(n_622),
.B(n_620),
.C(n_675),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_960),
.B(n_622),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1017),
.A2(n_371),
.B1(n_366),
.B2(n_361),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_893),
.B(n_593),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_SL g1082 ( 
.A1(n_1005),
.A2(n_663),
.B(n_672),
.C(n_655),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_937),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_894),
.B(n_680),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_862),
.B(n_680),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_913),
.A2(n_669),
.B(n_611),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_875),
.B(n_680),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_913),
.A2(n_669),
.B(n_611),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_955),
.A2(n_669),
.B(n_644),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_963),
.A2(n_672),
.B(n_663),
.C(n_655),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_1014),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_955),
.A2(n_644),
.B(n_485),
.Y(n_1092)
);

AO21x1_ASAP7_75t_L g1093 ( 
.A1(n_895),
.A2(n_557),
.B(n_558),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_959),
.A2(n_644),
.B(n_485),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_861),
.B(n_341),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_885),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_992),
.B(n_341),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_L g1098 ( 
.A(n_881),
.B(n_614),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_959),
.A2(n_485),
.B(n_628),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_871),
.A2(n_485),
.B(n_628),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_888),
.B(n_351),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_888),
.B(n_351),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_861),
.B(n_360),
.Y(n_1103)
);

BUFx4f_ASAP7_75t_L g1104 ( 
.A(n_975),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_915),
.B(n_360),
.C(n_273),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_908),
.B(n_628),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_944),
.A2(n_558),
.B(n_557),
.C(n_655),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_SL g1108 ( 
.A(n_923),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_871),
.A2(n_237),
.B(n_330),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_953),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_954),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_956),
.Y(n_1112)
);

BUFx4f_ASAP7_75t_L g1113 ( 
.A(n_934),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_1009),
.B(n_263),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_872),
.Y(n_1115)
);

CKINVDCx11_ASAP7_75t_R g1116 ( 
.A(n_905),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_916),
.B(n_265),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_916),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_864),
.B(n_934),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_965),
.B(n_279),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_871),
.A2(n_335),
.B(n_329),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_968),
.B(n_989),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1015),
.A2(n_328),
.B(n_322),
.C(n_319),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_976),
.B(n_315),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_976),
.B(n_314),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_969),
.A2(n_306),
.B(n_303),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_977),
.A2(n_300),
.B(n_299),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_854),
.A2(n_297),
.B(n_292),
.C(n_287),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_976),
.B(n_172),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_878),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_855),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_858),
.A2(n_169),
.B1(n_167),
.B2(n_166),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_933),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_949),
.A2(n_0),
.B(n_5),
.C(n_6),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_878),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_906),
.A2(n_159),
.B(n_145),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_901),
.B(n_144),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_906),
.A2(n_143),
.B(n_136),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_858),
.A2(n_5),
.B1(n_8),
.B2(n_11),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_906),
.A2(n_135),
.B(n_127),
.Y(n_1140)
);

AOI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_907),
.A2(n_14),
.B(n_15),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_901),
.B(n_115),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1016),
.B(n_111),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_906),
.A2(n_106),
.B(n_100),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_857),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_931),
.A2(n_97),
.B(n_96),
.Y(n_1146)
);

BUFx4_ASAP7_75t_SL g1147 ( 
.A(n_874),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_L g1148 ( 
.A(n_1011),
.B(n_17),
.C(n_23),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_889),
.B(n_23),
.Y(n_1149)
);

BUFx8_ASAP7_75t_L g1150 ( 
.A(n_941),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_881),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1016),
.B(n_75),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_996),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_960),
.B(n_24),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1021),
.A2(n_952),
.B1(n_869),
.B2(n_979),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1019),
.A2(n_935),
.B(n_856),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1022),
.A2(n_856),
.B(n_997),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1041),
.A2(n_950),
.B(n_964),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1033),
.A2(n_931),
.B(n_942),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1018),
.A2(n_1099),
.B(n_1094),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1092),
.A2(n_991),
.B(n_964),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1027),
.B(n_889),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1054),
.A2(n_991),
.B(n_982),
.Y(n_1163)
);

OAI22x1_ASAP7_75t_L g1164 ( 
.A1(n_1030),
.A2(n_900),
.B1(n_896),
.B2(n_866),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1071),
.Y(n_1165)
);

BUFx5_ASAP7_75t_L g1166 ( 
.A(n_1034),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1029),
.A2(n_979),
.B(n_1026),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1043),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1057),
.B(n_1010),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1023),
.B(n_858),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_SL g1171 ( 
.A(n_1020),
.B(n_1047),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1037),
.A2(n_884),
.B(n_882),
.C(n_887),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1038),
.A2(n_931),
.B(n_942),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1093),
.A2(n_999),
.B(n_997),
.Y(n_1174)
);

AO32x2_ASAP7_75t_L g1175 ( 
.A1(n_1133),
.A2(n_985),
.A3(n_933),
.B1(n_911),
.B2(n_858),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1042),
.A2(n_883),
.B(n_1006),
.C(n_999),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1104),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1106),
.A2(n_890),
.B(n_1012),
.C(n_880),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1104),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1069),
.A2(n_880),
.B(n_876),
.C(n_925),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1039),
.A2(n_1002),
.B(n_928),
.Y(n_1181)
);

AO21x1_ASAP7_75t_L g1182 ( 
.A1(n_1134),
.A2(n_1087),
.B(n_1085),
.Y(n_1182)
);

INVx3_ASAP7_75t_SL g1183 ( 
.A(n_1020),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1056),
.A2(n_983),
.B(n_982),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1053),
.B(n_868),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1097),
.B(n_868),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1089),
.A2(n_983),
.B(n_1002),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1112),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1027),
.B(n_995),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1148),
.A2(n_985),
.B1(n_925),
.B2(n_924),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1058),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1122),
.B(n_868),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1049),
.B(n_868),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1110),
.A2(n_979),
.B1(n_879),
.B2(n_897),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1061),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1111),
.B(n_919),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1032),
.A2(n_942),
.B(n_943),
.Y(n_1197)
);

AND2x6_ASAP7_75t_L g1198 ( 
.A(n_1154),
.B(n_897),
.Y(n_1198)
);

OAI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1025),
.A2(n_1083),
.B1(n_1044),
.B2(n_1060),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1131),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1118),
.B(n_919),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1034),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1046),
.A2(n_942),
.B(n_943),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1090),
.A2(n_928),
.B(n_924),
.Y(n_1204)
);

AOI221x1_ASAP7_75t_L g1205 ( 
.A1(n_1126),
.A2(n_946),
.B1(n_1007),
.B2(n_1004),
.C(n_1008),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1031),
.B(n_947),
.Y(n_1206)
);

AOI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1066),
.A2(n_1013),
.B(n_1007),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1024),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_SL g1209 ( 
.A(n_1113),
.B(n_911),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1120),
.B(n_947),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1153),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1055),
.A2(n_926),
.B(n_879),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1101),
.B(n_995),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1109),
.A2(n_926),
.B(n_980),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1113),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_1051),
.A2(n_912),
.A3(n_948),
.B1(n_995),
.B2(n_972),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_1076),
.B(n_1088),
.Y(n_1217)
);

AND2x6_ASAP7_75t_L g1218 ( 
.A(n_1154),
.B(n_940),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1078),
.A2(n_966),
.A3(n_936),
.B(n_920),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1086),
.A2(n_917),
.B(n_1003),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1143),
.A2(n_940),
.B(n_948),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1141),
.B(n_948),
.C(n_32),
.Y(n_1222)
);

OAI22x1_ASAP7_75t_L g1223 ( 
.A1(n_1059),
.A2(n_1117),
.B1(n_1119),
.B2(n_1064),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1107),
.A2(n_948),
.B(n_35),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1152),
.A2(n_26),
.B(n_36),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1048),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1091),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_SL g1228 ( 
.A(n_1061),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1074),
.A2(n_37),
.B(n_39),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1102),
.B(n_1149),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1136),
.A2(n_37),
.B(n_39),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1067),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1050),
.B(n_52),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1082),
.A2(n_53),
.B(n_55),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1045),
.A2(n_55),
.B(n_56),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1100),
.A2(n_56),
.B(n_57),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1123),
.A2(n_57),
.B(n_58),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1124),
.A2(n_1125),
.B(n_1129),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1137),
.A2(n_1142),
.B(n_1077),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1028),
.B(n_1114),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1128),
.A2(n_1081),
.B(n_1084),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1127),
.B(n_1095),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1075),
.B(n_1103),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1034),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1139),
.A2(n_1105),
.B1(n_1065),
.B2(n_1080),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1132),
.A2(n_1138),
.B(n_1144),
.C(n_1146),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1098),
.A2(n_1140),
.B(n_1040),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1079),
.A2(n_1062),
.B(n_1121),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_1034),
.Y(n_1249)
);

AOI221x1_ASAP7_75t_L g1250 ( 
.A1(n_1051),
.A2(n_1130),
.B1(n_1073),
.B2(n_1072),
.C(n_1052),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1052),
.A2(n_1063),
.B(n_1130),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1063),
.A2(n_1073),
.B(n_1151),
.Y(n_1252)
);

AOI221x1_ASAP7_75t_L g1253 ( 
.A1(n_1115),
.A2(n_1135),
.B1(n_1068),
.B2(n_1147),
.C(n_1116),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1063),
.A2(n_1135),
.A3(n_1108),
.B(n_1150),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1096),
.B(n_1063),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1108),
.A2(n_1150),
.B(n_1019),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1043),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1041),
.A2(n_1018),
.B(n_987),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1023),
.B(n_957),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_SL g1260 ( 
.A(n_1048),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1019),
.A2(n_938),
.B(n_927),
.C(n_706),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1096),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1023),
.B(n_957),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1023),
.B(n_957),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1023),
.B(n_957),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1043),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_1020),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1043),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1093),
.A2(n_1090),
.A3(n_1019),
.B(n_1078),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1030),
.A2(n_938),
.B1(n_927),
.B2(n_707),
.Y(n_1270)
);

AO32x2_ASAP7_75t_L g1271 ( 
.A1(n_1133),
.A2(n_1019),
.A3(n_951),
.B1(n_1051),
.B2(n_990),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_1024),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1043),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1034),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1023),
.B(n_957),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1019),
.A2(n_1038),
.B(n_1033),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1149),
.A2(n_1087),
.B(n_1085),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1022),
.A2(n_1019),
.B(n_969),
.Y(n_1278)
);

NOR3xp33_ASAP7_75t_L g1279 ( 
.A(n_1030),
.B(n_938),
.C(n_927),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1104),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1027),
.B(n_960),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1019),
.A2(n_1038),
.B(n_1033),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1023),
.B(n_957),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1023),
.B(n_957),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_R g1285 ( 
.A(n_1096),
.B(n_561),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1019),
.A2(n_1038),
.B(n_1033),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1021),
.A2(n_938),
.B1(n_927),
.B2(n_706),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1058),
.B(n_865),
.Y(n_1288)
);

NOR3xp33_ASAP7_75t_L g1289 ( 
.A(n_1030),
.B(n_938),
.C(n_927),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1020),
.Y(n_1290)
);

AOI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_1057),
.A2(n_791),
.B1(n_962),
.B2(n_932),
.C(n_938),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1019),
.A2(n_938),
.B(n_927),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1035),
.A2(n_938),
.B(n_927),
.C(n_1036),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1214),
.A2(n_1174),
.B(n_1197),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1250),
.A2(n_1278),
.B(n_1217),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1278),
.A2(n_1160),
.B(n_1258),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1292),
.A2(n_1279),
.B(n_1289),
.C(n_1261),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1189),
.B(n_1252),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1168),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1291),
.A2(n_1270),
.B1(n_1287),
.B2(n_1293),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1270),
.A2(n_1169),
.B1(n_1245),
.B2(n_1264),
.Y(n_1301)
);

BUFx4f_ASAP7_75t_SL g1302 ( 
.A(n_1183),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1230),
.B(n_1165),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1200),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1290),
.B(n_1262),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1213),
.B(n_1255),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1158),
.A2(n_1220),
.B(n_1187),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1203),
.A2(n_1207),
.B(n_1247),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1259),
.B(n_1263),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1222),
.A2(n_1240),
.B1(n_1286),
.B2(n_1237),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1265),
.B(n_1275),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1222),
.A2(n_1284),
.B1(n_1283),
.B2(n_1206),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1208),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1257),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1266),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1268),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1273),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1212),
.A2(n_1204),
.B(n_1277),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1191),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1211),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1165),
.B(n_1188),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1201),
.B(n_1188),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1224),
.A2(n_1156),
.B(n_1232),
.C(n_1225),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1224),
.A2(n_1157),
.B(n_1181),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1237),
.A2(n_1190),
.B1(n_1164),
.B2(n_1199),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1219),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1178),
.A2(n_1172),
.B(n_1176),
.C(n_1256),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1248),
.A2(n_1229),
.B(n_1241),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1219),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1205),
.A2(n_1251),
.B(n_1234),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1235),
.A2(n_1236),
.B(n_1182),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1241),
.A2(n_1180),
.B(n_1246),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1185),
.A2(n_1239),
.A3(n_1194),
.B(n_1192),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_SL g1334 ( 
.A1(n_1242),
.A2(n_1186),
.B(n_1193),
.C(n_1170),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1221),
.A2(n_1167),
.B(n_1159),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1238),
.B(n_1155),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1223),
.B(n_1210),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1202),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1173),
.A2(n_1231),
.B(n_1244),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1233),
.A2(n_1243),
.B(n_1196),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1227),
.B(n_1288),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1272),
.B(n_1209),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

NAND2x1p5_ASAP7_75t_L g1344 ( 
.A(n_1274),
.B(n_1281),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1281),
.B(n_1171),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1215),
.B(n_1162),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1290),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1162),
.A2(n_1271),
.B(n_1216),
.C(n_1175),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1226),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1269),
.A2(n_1166),
.B(n_1253),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1166),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1166),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1269),
.A2(n_1166),
.B(n_1249),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1177),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1285),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1216),
.A2(n_1271),
.B(n_1175),
.Y(n_1356)
);

CKINVDCx16_ASAP7_75t_R g1357 ( 
.A(n_1260),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1271),
.A2(n_1175),
.B(n_1179),
.C(n_1280),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1179),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1198),
.A2(n_1218),
.B(n_1195),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1254),
.A2(n_1198),
.B(n_1218),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1254),
.A2(n_1198),
.B(n_1218),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1198),
.A2(n_1218),
.B1(n_1260),
.B2(n_1228),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1228),
.A2(n_1195),
.B(n_1280),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1280),
.A2(n_1292),
.B(n_1278),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_1279),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1285),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1214),
.A2(n_1174),
.B(n_1197),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_1279),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1250),
.A2(n_1278),
.B(n_1217),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_1291),
.C(n_1282),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1213),
.B(n_1097),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1202),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1163),
.A2(n_1184),
.B(n_1161),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1259),
.B(n_1263),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1213),
.B(n_1097),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1168),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1290),
.B(n_796),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1213),
.B(n_1097),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1163),
.A2(n_1184),
.B(n_1161),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1267),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1250),
.A2(n_1278),
.B(n_1217),
.Y(n_1382)
);

CKINVDCx11_ASAP7_75t_R g1383 ( 
.A(n_1183),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1287),
.B(n_1292),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_1291),
.C(n_1282),
.Y(n_1385)
);

AO31x2_ASAP7_75t_L g1386 ( 
.A1(n_1251),
.A2(n_1250),
.A3(n_1093),
.B(n_1217),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1291),
.A2(n_1289),
.B1(n_1279),
.B2(n_1292),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1267),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1168),
.Y(n_1389)
);

AOI21xp33_ASAP7_75t_L g1390 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_938),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_1291),
.C(n_1282),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1163),
.A2(n_1184),
.B(n_1161),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1189),
.B(n_1252),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1267),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1292),
.A2(n_1261),
.B(n_1291),
.C(n_1282),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1183),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1291),
.A2(n_1289),
.B1(n_1279),
.B2(n_1292),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1287),
.B(n_1292),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1183),
.Y(n_1399)
);

OR2x6_ASAP7_75t_L g1400 ( 
.A(n_1256),
.B(n_1167),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1260),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1168),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1292),
.A2(n_1282),
.B(n_1276),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1168),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_SL g1405 ( 
.A1(n_1292),
.A2(n_1293),
.B(n_1261),
.C(n_1145),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1251),
.A2(n_1250),
.A3(n_1093),
.B(n_1217),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1292),
.A2(n_1282),
.B(n_1276),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1168),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1259),
.B(n_1263),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1291),
.A2(n_1289),
.B1(n_1279),
.B2(n_1292),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1214),
.A2(n_1174),
.B(n_1197),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1250),
.A2(n_1278),
.B(n_1217),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1292),
.A2(n_1293),
.B(n_1261),
.C(n_1145),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1168),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1168),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1259),
.B(n_1263),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1292),
.A2(n_1282),
.B(n_1276),
.Y(n_1417)
);

AO31x2_ASAP7_75t_L g1418 ( 
.A1(n_1251),
.A2(n_1250),
.A3(n_1093),
.B(n_1217),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1321),
.B(n_1341),
.Y(n_1419)
);

CKINVDCx6p67_ASAP7_75t_R g1420 ( 
.A(n_1383),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1322),
.B(n_1309),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1387),
.A2(n_1397),
.B1(n_1410),
.B2(n_1398),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1384),
.B(n_1398),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1384),
.A2(n_1297),
.B(n_1390),
.C(n_1366),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1376),
.B(n_1379),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1303),
.B(n_1311),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1371),
.A2(n_1395),
.B(n_1385),
.C(n_1391),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1387),
.A2(n_1397),
.B1(n_1410),
.B2(n_1300),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1403),
.A2(n_1417),
.B(n_1407),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1385),
.A2(n_1391),
.B1(n_1395),
.B2(n_1301),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1303),
.B(n_1375),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1323),
.A2(n_1310),
.B1(n_1416),
.B2(n_1409),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1405),
.A2(n_1413),
.B(n_1327),
.C(n_1337),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1312),
.B(n_1365),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1348),
.A2(n_1358),
.B1(n_1325),
.B2(n_1342),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1307),
.A2(n_1318),
.B(n_1328),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1332),
.A2(n_1296),
.B(n_1405),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1314),
.Y(n_1441)
);

O2A1O1Ixp5_ASAP7_75t_L g1442 ( 
.A1(n_1294),
.A2(n_1411),
.B(n_1368),
.C(n_1351),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1383),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1365),
.B(n_1319),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1388),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1400),
.A2(n_1360),
.B(n_1345),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1351),
.A2(n_1358),
.B(n_1352),
.C(n_1348),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1325),
.B(n_1298),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1413),
.A2(n_1340),
.B(n_1334),
.C(n_1400),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1396),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1302),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1315),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1298),
.B(n_1393),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1316),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1344),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1393),
.B(n_1317),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1320),
.B(n_1334),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1353),
.A2(n_1374),
.B(n_1380),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1400),
.A2(n_1336),
.B(n_1345),
.C(n_1313),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1356),
.A2(n_1363),
.B1(n_1389),
.B2(n_1299),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1336),
.A2(n_1402),
.B(n_1377),
.C(n_1415),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1356),
.A2(n_1363),
.B1(n_1414),
.B2(n_1304),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1356),
.A2(n_1332),
.B1(n_1408),
.B2(n_1404),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1333),
.B(n_1324),
.Y(n_1464)
);

O2A1O1Ixp5_ASAP7_75t_L g1465 ( 
.A1(n_1352),
.A2(n_1326),
.B(n_1329),
.C(n_1338),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1349),
.B(n_1333),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1333),
.B(n_1324),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1346),
.B(n_1359),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1346),
.B(n_1359),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1388),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1350),
.B(n_1339),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1357),
.A2(n_1295),
.B1(n_1412),
.B2(n_1382),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1381),
.A2(n_1305),
.B(n_1347),
.C(n_1378),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1333),
.B(n_1295),
.Y(n_1474)
);

AOI21x1_ASAP7_75t_SL g1475 ( 
.A1(n_1401),
.A2(n_1339),
.B(n_1335),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1396),
.A2(n_1344),
.B(n_1331),
.C(n_1373),
.Y(n_1476)
);

INVxp33_ASAP7_75t_SL g1477 ( 
.A(n_1355),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1302),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1399),
.B(n_1367),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1370),
.B(n_1382),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1394),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1367),
.A2(n_1399),
.B(n_1354),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1370),
.A2(n_1412),
.B1(n_1343),
.B2(n_1388),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1343),
.B(n_1364),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1370),
.B(n_1330),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1401),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1386),
.B(n_1406),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1308),
.B(n_1392),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1418),
.A2(n_1292),
.B(n_1403),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1418),
.A2(n_1292),
.B(n_1261),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1418),
.B(n_1306),
.Y(n_1491)
);

NOR2xp67_ASAP7_75t_L g1492 ( 
.A(n_1399),
.B(n_1355),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1399),
.B(n_1355),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1390),
.A2(n_1292),
.B(n_1261),
.C(n_1289),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1496)
);

CKINVDCx14_ASAP7_75t_R g1497 ( 
.A(n_1383),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1298),
.B(n_1393),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1383),
.Y(n_1500)
);

NAND2x1p5_ASAP7_75t_L g1501 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1384),
.B(n_1398),
.Y(n_1502)
);

O2A1O1Ixp5_ASAP7_75t_L g1503 ( 
.A1(n_1390),
.A2(n_1292),
.B(n_1398),
.C(n_1384),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1384),
.A2(n_1292),
.B(n_1291),
.C(n_1398),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1403),
.A2(n_1292),
.B(n_1407),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1384),
.B(n_1398),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1403),
.A2(n_1292),
.B(n_1407),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_SL g1509 ( 
.A(n_1400),
.B(n_1336),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1387),
.A2(n_1291),
.B1(n_1410),
.B2(n_1397),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1511)
);

CKINVDCx6p67_ASAP7_75t_R g1512 ( 
.A(n_1383),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1371),
.A2(n_1292),
.B(n_1261),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1463),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1463),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1423),
.B(n_1502),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1474),
.B(n_1485),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1487),
.B(n_1491),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1508),
.A2(n_1505),
.B(n_1431),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1441),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1480),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1452),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1508),
.A2(n_1431),
.B(n_1489),
.Y(n_1524)
);

BUFx4f_ASAP7_75t_SL g1525 ( 
.A(n_1420),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1454),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1458),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1472),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1440),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1458),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1446),
.B(n_1459),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1498),
.B(n_1471),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1423),
.B(n_1502),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1510),
.A2(n_1422),
.B1(n_1430),
.B2(n_1504),
.Y(n_1534)
);

BUFx4f_ASAP7_75t_SL g1535 ( 
.A(n_1512),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1503),
.A2(n_1424),
.B(n_1513),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1457),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1439),
.A2(n_1490),
.B(n_1483),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1457),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1427),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1472),
.B(n_1483),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1460),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1464),
.B(n_1467),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1456),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1477),
.B(n_1428),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1464),
.A2(n_1467),
.B(n_1506),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1460),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1456),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1436),
.B(n_1466),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1475),
.A2(n_1442),
.B(n_1495),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1495),
.A2(n_1501),
.B(n_1465),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1436),
.B(n_1444),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1471),
.B(n_1447),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1448),
.B(n_1453),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1448),
.B(n_1453),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1509),
.B(n_1488),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1484),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1462),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1427),
.A2(n_1432),
.B(n_1437),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1437),
.B(n_1501),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1438),
.B(n_1488),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1449),
.A2(n_1476),
.B(n_1435),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1429),
.B(n_1461),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1422),
.A2(n_1430),
.B(n_1494),
.Y(n_1564)
);

OR2x6_ASAP7_75t_SL g1565 ( 
.A(n_1549),
.B(n_1510),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1521),
.Y(n_1566)
);

INVx5_ASAP7_75t_L g1567 ( 
.A(n_1529),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1522),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1521),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1561),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1546),
.B(n_1544),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1518),
.B(n_1552),
.Y(n_1572)
);

BUFx2_ASAP7_75t_SL g1573 ( 
.A(n_1529),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1546),
.B(n_1434),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1523),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1518),
.B(n_1419),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1546),
.B(n_1434),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1518),
.B(n_1421),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1561),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1519),
.B(n_1425),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1534),
.B(n_1433),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1519),
.B(n_1514),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1534),
.A2(n_1426),
.B1(n_1511),
.B2(n_1499),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1556),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1526),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1507),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1543),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1532),
.B(n_1455),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1564),
.A2(n_1497),
.B1(n_1450),
.B2(n_1486),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1549),
.B(n_1528),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1469),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1537),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1468),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1536),
.A2(n_1540),
.B1(n_1517),
.B2(n_1533),
.C1(n_1525),
.C2(n_1535),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1553),
.B(n_1455),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1565),
.A2(n_1536),
.B1(n_1559),
.B2(n_1563),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1589),
.B(n_1532),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1566),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1572),
.B(n_1537),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1567),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1565),
.A2(n_1559),
.B1(n_1563),
.B2(n_1533),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1586),
.A2(n_1563),
.B1(n_1559),
.B2(n_1531),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

AOI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1581),
.A2(n_1577),
.B1(n_1574),
.B2(n_1540),
.C(n_1583),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1567),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1591),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1581),
.B(n_1545),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1575),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1571),
.A2(n_1551),
.B(n_1550),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_R g1614 ( 
.A(n_1583),
.B(n_1443),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1590),
.A2(n_1531),
.B1(n_1559),
.B2(n_1563),
.C(n_1473),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1590),
.A2(n_1563),
.B1(n_1531),
.B2(n_1542),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1574),
.A2(n_1564),
.B1(n_1547),
.B2(n_1542),
.C(n_1558),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1586),
.A2(n_1531),
.B1(n_1547),
.B2(n_1588),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1577),
.A2(n_1527),
.B(n_1530),
.Y(n_1620)
);

BUFx10_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1594),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1596),
.A2(n_1531),
.B1(n_1560),
.B2(n_1528),
.C(n_1558),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1586),
.A2(n_1531),
.B1(n_1560),
.B2(n_1555),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1576),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_SL g1626 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1626)
);

AOI331xp33_ASAP7_75t_L g1627 ( 
.A1(n_1585),
.A2(n_1564),
.A3(n_1548),
.B1(n_1544),
.B2(n_1539),
.B3(n_1515),
.C1(n_1516),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1593),
.B(n_1557),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_R g1630 ( 
.A(n_1597),
.B(n_1500),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1594),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1571),
.A2(n_1527),
.B(n_1530),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1596),
.A2(n_1525),
.B1(n_1451),
.B2(n_1450),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1578),
.B(n_1555),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1578),
.B(n_1555),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1568),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1600),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1630),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1632),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_SL g1640 ( 
.A(n_1608),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1617),
.B(n_1606),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1602),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1632),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1610),
.B(n_1570),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1602),
.B(n_1562),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1622),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1623),
.A2(n_1562),
.B(n_1560),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1621),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1612),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1608),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1620),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1628),
.B(n_1579),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1601),
.Y(n_1659)
);

NOR2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1625),
.B(n_1584),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1631),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1621),
.Y(n_1662)
);

INVx4_ASAP7_75t_SL g1663 ( 
.A(n_1633),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1613),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1637),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1660),
.B(n_1644),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1637),
.Y(n_1668)
);

NOR3xp33_ASAP7_75t_L g1669 ( 
.A(n_1641),
.B(n_1623),
.C(n_1615),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1659),
.B(n_1587),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1599),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1599),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1642),
.B(n_1629),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1642),
.B(n_1592),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1661),
.B(n_1634),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1638),
.B(n_1611),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1616),
.C(n_1598),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1663),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1646),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1649),
.B(n_1636),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1660),
.B(n_1595),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1653),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1644),
.B(n_1597),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1661),
.B(n_1635),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1597),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1644),
.B(n_1592),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1658),
.B(n_1619),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1640),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1653),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1648),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1653),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

NAND2xp33_ASAP7_75t_L g1695 ( 
.A(n_1650),
.B(n_1614),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1663),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1648),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1652),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1651),
.B(n_1580),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1651),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1669),
.A2(n_1663),
.B1(n_1616),
.B2(n_1564),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1679),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1669),
.B(n_1580),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1701),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1656),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1670),
.A2(n_1598),
.B1(n_1603),
.B2(n_1604),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_1580),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1701),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1679),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1682),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1674),
.B(n_1696),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1690),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1666),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1666),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1682),
.B(n_1656),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1674),
.B(n_1582),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1668),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1676),
.B(n_1652),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1696),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1690),
.B(n_1694),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1685),
.B(n_1656),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1674),
.B(n_1678),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1678),
.B(n_1582),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1655),
.Y(n_1726)
);

NOR2xp67_ASAP7_75t_L g1727 ( 
.A(n_1690),
.B(n_1694),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.B(n_1663),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1668),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1694),
.B(n_1665),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1687),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1683),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1694),
.B(n_1663),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1686),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1687),
.B(n_1654),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1680),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1673),
.B(n_1654),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1729),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1729),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1728),
.B(n_1711),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1734),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1710),
.B(n_1677),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1728),
.B(n_1711),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1720),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1736),
.Y(n_1745)
);

AND2x4_ASAP7_75t_SL g1746 ( 
.A(n_1724),
.B(n_1733),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1717),
.B(n_1699),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1723),
.B(n_1672),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1713),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1706),
.B(n_1737),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1712),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1704),
.B(n_1686),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1702),
.A2(n_1671),
.B1(n_1662),
.B2(n_1654),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1707),
.A2(n_1671),
.B1(n_1624),
.B2(n_1673),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1724),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1736),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1714),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1725),
.A2(n_1695),
.B1(n_1524),
.B2(n_1520),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1706),
.B(n_1673),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1719),
.B(n_1699),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1713),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1737),
.B(n_1724),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1733),
.A2(n_1624),
.B1(n_1688),
.B2(n_1618),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1715),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1758),
.A2(n_1733),
.B1(n_1727),
.B2(n_1708),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1738),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1758),
.A2(n_1721),
.B1(n_1731),
.B2(n_1719),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1740),
.B(n_1721),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1740),
.B(n_1721),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1753),
.B(n_1730),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1739),
.Y(n_1771)
);

AOI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1754),
.A2(n_1705),
.B1(n_1709),
.B2(n_1718),
.C(n_1716),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1743),
.B(n_1735),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1746),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1746),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1745),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1743),
.B(n_1735),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1742),
.Y(n_1778)
);

OAI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1763),
.A2(n_1647),
.B1(n_1662),
.B2(n_1689),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1756),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1741),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1750),
.Y(n_1782)
);

AOI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1751),
.A2(n_1726),
.B(n_1716),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1750),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1759),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1778),
.B(n_1755),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1784),
.B(n_1762),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1773),
.B(n_1762),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1785),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1773),
.B(n_1744),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1777),
.B(n_1748),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_SL g1792 ( 
.A(n_1774),
.B(n_1451),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_SL g1793 ( 
.A(n_1775),
.B(n_1759),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1777),
.B(n_1749),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1782),
.B(n_1749),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1768),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1769),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1793),
.A2(n_1772),
.B1(n_1770),
.B2(n_1782),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1789),
.Y(n_1799)
);

O2A1O1Ixp33_ASAP7_75t_SL g1800 ( 
.A1(n_1787),
.A2(n_1770),
.B(n_1785),
.C(n_1783),
.Y(n_1800)
);

NOR4xp25_ASAP7_75t_L g1801 ( 
.A(n_1796),
.B(n_1781),
.C(n_1766),
.D(n_1780),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1792),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1797),
.B(n_1761),
.Y(n_1803)
);

NAND4xp25_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1765),
.C(n_1767),
.D(n_1771),
.Y(n_1804)
);

OAI211xp5_ASAP7_75t_L g1805 ( 
.A1(n_1794),
.A2(n_1776),
.B(n_1766),
.C(n_1761),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1788),
.A2(n_1779),
.B1(n_1790),
.B2(n_1791),
.C(n_1795),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1789),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1786),
.A2(n_1764),
.B1(n_1757),
.B2(n_1752),
.C(n_1760),
.Y(n_1808)
);

AOI211x1_ASAP7_75t_SL g1809 ( 
.A1(n_1787),
.A2(n_1732),
.B(n_1693),
.C(n_1697),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1803),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1799),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_SL g1812 ( 
.A(n_1802),
.B(n_1478),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1798),
.A2(n_1760),
.B1(n_1747),
.B2(n_1726),
.Y(n_1813)
);

XOR2xp5_ASAP7_75t_L g1814 ( 
.A(n_1804),
.B(n_1747),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1807),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1810),
.B(n_1801),
.Y(n_1816)
);

NOR2xp67_ASAP7_75t_L g1817 ( 
.A(n_1813),
.B(n_1805),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1814),
.B(n_1806),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1812),
.B(n_1800),
.Y(n_1819)
);

AOI221x1_ASAP7_75t_L g1820 ( 
.A1(n_1815),
.A2(n_1732),
.B1(n_1809),
.B2(n_1722),
.C(n_1683),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1812),
.B(n_1808),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1811),
.B(n_1722),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1821),
.Y(n_1823)
);

NOR2xp67_ASAP7_75t_L g1824 ( 
.A(n_1819),
.B(n_1479),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1816),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1817),
.A2(n_1818),
.B(n_1822),
.Y(n_1826)
);

AOI332xp33_ASAP7_75t_L g1827 ( 
.A1(n_1820),
.A2(n_1683),
.A3(n_1693),
.B1(n_1691),
.B2(n_1697),
.B3(n_1664),
.C1(n_1643),
.C2(n_1684),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1824),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1823),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1826),
.Y(n_1830)
);

NAND2x1_ASAP7_75t_L g1831 ( 
.A(n_1830),
.B(n_1827),
.Y(n_1831)
);

NOR3xp33_ASAP7_75t_L g1832 ( 
.A(n_1831),
.B(n_1830),
.C(n_1829),
.Y(n_1832)
);

AO22x2_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1825),
.B1(n_1828),
.B2(n_1697),
.Y(n_1833)
);

AOI31xp67_ASAP7_75t_L g1834 ( 
.A1(n_1832),
.A2(n_1691),
.A3(n_1693),
.B(n_1664),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1833),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1834),
.Y(n_1836)
);

XNOR2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1835),
.B(n_1492),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1836),
.A2(n_1481),
.B1(n_1445),
.B2(n_1470),
.Y(n_1838)
);

OAI22x1_ASAP7_75t_L g1839 ( 
.A1(n_1837),
.A2(n_1665),
.B1(n_1691),
.B2(n_1664),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1838),
.B1(n_1665),
.B2(n_1684),
.C(n_1680),
.Y(n_1840)
);

OA21x2_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1681),
.B(n_1665),
.Y(n_1841)
);

OAI222xp33_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1664),
.B1(n_1643),
.B2(n_1639),
.C1(n_1657),
.C2(n_1698),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1493),
.B1(n_1675),
.B2(n_1688),
.Y(n_1843)
);

AOI211xp5_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1482),
.B(n_1692),
.C(n_1698),
.Y(n_1844)
);


endmodule