module fake_jpeg_10971_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_31),
.B(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_52),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_25),
.B(n_1),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_28),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_29),
.C(n_23),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_70),
.CI(n_76),
.CON(n_96),
.SN(n_96)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_13),
.B(n_23),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_61),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_13),
.B1(n_24),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_73),
.B1(n_77),
.B2(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_64),
.B(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_9),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_28),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_85),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_3),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_43),
.C(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_49),
.Y(n_85)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_92),
.Y(n_109)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_56),
.B1(n_55),
.B2(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_94),
.B1(n_104),
.B2(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_72),
.B1(n_78),
.B2(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_104),
.C(n_101),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_98),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_68),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_105),
.Y(n_126)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_84),
.CON(n_115),
.SN(n_115)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_79),
.B1(n_57),
.B2(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_68),
.Y(n_117)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_68),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_115),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_118),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_94),
.B(n_97),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_112),
.B(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_125),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_83),
.B1(n_107),
.B2(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_86),
.B1(n_89),
.B2(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_122),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_120),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_91),
.B1(n_114),
.B2(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_141),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_134),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_110),
.B(n_117),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_122),
.C(n_111),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_110),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_145),
.C(n_146),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_136),
.C(n_134),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_111),
.B(n_124),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_151),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_128),
.B(n_129),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.Y(n_163)
);

XNOR2x2_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_133),
.B1(n_138),
.B2(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_164),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_144),
.C(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_158),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_154),
.C(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_159),
.C(n_155),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_156),
.C(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_157),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_147),
.B(n_121),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_175),
.Y(n_176)
);


endmodule