module fake_jpeg_29112_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx11_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_40),
.B1(n_39),
.B2(n_41),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_58),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_35),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_76)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_76),
.B1(n_5),
.B2(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_1),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_3),
.B(n_4),
.Y(n_81)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_6),
.CI(n_7),
.CON(n_83),
.SN(n_83)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_16),
.C(n_32),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_14),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_62),
.B1(n_63),
.B2(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_82),
.B1(n_76),
.B2(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_87),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_7),
.B(n_8),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_95),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_19),
.B1(n_21),
.B2(n_25),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_88),
.C(n_83),
.Y(n_100)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_11),
.B(n_17),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_10),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_34),
.B(n_13),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_104),
.C(n_98),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_90),
.B1(n_98),
.B2(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_105),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_99),
.B(n_96),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_26),
.B(n_27),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_28),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_31),
.C(n_94),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_91),
.C(n_112),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_114),
.Y(n_115)
);


endmodule