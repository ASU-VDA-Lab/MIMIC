module real_aes_16422_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AND2x4_ASAP7_75t_L g117 ( .A(n_0), .B(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_1), .A2(n_4), .B1(n_270), .B2(n_271), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_2), .A2(n_42), .B1(n_171), .B2(n_219), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_3), .A2(n_24), .B1(n_219), .B2(n_253), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_5), .A2(n_16), .B1(n_520), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_6), .A2(n_59), .B1(n_156), .B2(n_157), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_7), .A2(n_17), .B1(n_171), .B2(n_172), .Y(n_170) );
INVx1_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_9), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_10), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_11), .A2(n_18), .B1(n_521), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_12), .A2(n_132), .B1(n_796), .B2(n_797), .Y(n_131) );
INVx1_ASAP7_75t_L g796 ( .A(n_12), .Y(n_796) );
BUFx2_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
OR2x2_ASAP7_75t_L g130 ( .A(n_13), .B(n_37), .Y(n_130) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_14), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_15), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_19), .A2(n_96), .B1(n_271), .B2(n_520), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_20), .A2(n_38), .B1(n_149), .B2(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_21), .B(n_147), .Y(n_581) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_22), .A2(n_57), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_23), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_25), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_26), .B(n_144), .Y(n_211) );
INVx4_ASAP7_75t_R g195 ( .A(n_27), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_28), .A2(n_46), .B1(n_175), .B2(n_268), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_29), .A2(n_53), .B1(n_175), .B2(n_520), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_30), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_31), .B(n_545), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_32), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_33), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g275 ( .A(n_34), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_SL g250 ( .A1(n_35), .A2(n_143), .B(n_171), .C(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_36), .A2(n_54), .B1(n_171), .B2(n_175), .Y(n_259) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_37), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_39), .A2(n_84), .B1(n_171), .B2(n_512), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_40), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_40), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_41), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_43), .A2(n_45), .B1(n_171), .B2(n_172), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_44), .A2(n_58), .B1(n_520), .B2(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g215 ( .A(n_47), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_48), .B(n_171), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_49), .Y(n_229) );
INVx2_ASAP7_75t_L g125 ( .A(n_50), .Y(n_125) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
BUFx3_ASAP7_75t_L g128 ( .A(n_51), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_52), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_55), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_56), .A2(n_85), .B1(n_171), .B2(n_175), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_60), .A2(n_73), .B1(n_268), .B2(n_537), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_61), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_62), .A2(n_76), .B1(n_171), .B2(n_172), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_63), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_64), .A2(n_95), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g162 ( .A(n_65), .Y(n_162) );
AND2x4_ASAP7_75t_L g165 ( .A(n_66), .B(n_166), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_67), .A2(n_87), .B1(n_175), .B2(n_268), .Y(n_267) );
AO22x1_ASAP7_75t_L g145 ( .A1(n_68), .A2(n_74), .B1(n_146), .B2(n_149), .Y(n_145) );
INVx1_ASAP7_75t_L g166 ( .A(n_69), .Y(n_166) );
AND2x2_ASAP7_75t_L g254 ( .A(n_70), .B(n_207), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_71), .B(n_156), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_72), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_75), .B(n_219), .Y(n_230) );
INVx2_ASAP7_75t_L g144 ( .A(n_77), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_78), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_79), .B(n_207), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_80), .A2(n_94), .B1(n_156), .B2(n_175), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_81), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_82), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_83), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_86), .B(n_207), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_88), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_89), .B(n_207), .Y(n_226) );
INVx1_ASAP7_75t_L g116 ( .A(n_90), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_90), .B(n_805), .Y(n_804) );
NAND2xp33_ASAP7_75t_L g584 ( .A(n_91), .B(n_147), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_92), .A2(n_156), .B(n_177), .C(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g200 ( .A(n_93), .B(n_201), .Y(n_200) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_97), .B(n_196), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_98), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_119), .B(n_828), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx4_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx4_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx5_ASAP7_75t_L g830 ( .A(n_104), .Y(n_830) );
OR2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_110), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR2x1p5_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
AND3x2_ASAP7_75t_L g819 ( .A(n_111), .B(n_115), .C(n_129), .Y(n_819) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g805 ( .A(n_112), .Y(n_805) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g492 ( .A(n_116), .Y(n_492) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_806), .Y(n_119) );
OAI21xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_131), .B(n_798), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
BUFx12f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x6_ASAP7_75t_SL g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g809 ( .A(n_125), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_125), .B(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2x1_ASAP7_75t_L g827 ( .A(n_128), .B(n_130), .Y(n_827) );
AND2x6_ASAP7_75t_SL g803 ( .A(n_129), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g797 ( .A(n_132), .Y(n_797) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_490), .B1(n_493), .B2(n_795), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_400), .Y(n_134) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_329), .C(n_371), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_303), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_202), .B1(n_278), .B2(n_289), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_183), .Y(n_139) );
AOI21xp33_ASAP7_75t_L g322 ( .A1(n_140), .A2(n_323), .B(n_325), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_140), .A2(n_396), .B(n_397), .Y(n_395) );
OR2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_167), .Y(n_140) );
INVx2_ASAP7_75t_L g315 ( .A(n_141), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_141), .B(n_168), .Y(n_345) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_151), .C(n_163), .Y(n_142) );
INVx6_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_143), .A2(n_234), .B(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_143), .B(n_145), .Y(n_287) );
O2A1O1Ixp5_ASAP7_75t_L g579 ( .A1(n_143), .A2(n_172), .B(n_580), .C(n_581), .Y(n_579) );
BUFx8_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx1_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
INVx1_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
INVxp67_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g520 ( .A(n_147), .Y(n_520) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g150 ( .A(n_148), .Y(n_150) );
INVx1_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
INVx3_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_148), .Y(n_197) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_148), .Y(n_219) );
INVx1_ASAP7_75t_L g247 ( .A(n_148), .Y(n_247) );
INVx2_ASAP7_75t_L g253 ( .A(n_148), .Y(n_253) );
OAI21xp33_ASAP7_75t_SL g210 ( .A1(n_149), .A2(n_211), .B(n_212), .Y(n_210) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g286 ( .A(n_151), .Y(n_286) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_159), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_152), .A2(n_217), .B(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_152), .A2(n_173), .B1(n_258), .B2(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g503 ( .A(n_153), .Y(n_503) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
INVx1_ASAP7_75t_L g565 ( .A(n_157), .Y(n_565) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_158), .B(n_192), .Y(n_191) );
OAI21xp33_ASAP7_75t_L g163 ( .A1(n_159), .A2(n_160), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g178 ( .A(n_160), .Y(n_178) );
INVx2_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
INVx2_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
INVx1_ASAP7_75t_L g288 ( .A(n_163), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_164), .A2(n_243), .B(n_250), .Y(n_242) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx10_ASAP7_75t_L g179 ( .A(n_165), .Y(n_179) );
BUFx10_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
INVx1_ASAP7_75t_L g273 ( .A(n_165), .Y(n_273) );
AND2x2_ASAP7_75t_L g385 ( .A(n_167), .B(n_224), .Y(n_385) );
INVx1_ASAP7_75t_L g418 ( .A(n_167), .Y(n_418) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g280 ( .A(n_168), .B(n_225), .Y(n_280) );
AND2x2_ASAP7_75t_L g311 ( .A(n_168), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g320 ( .A(n_168), .Y(n_320) );
OR2x2_ASAP7_75t_L g339 ( .A(n_168), .B(n_185), .Y(n_339) );
AND2x2_ASAP7_75t_L g354 ( .A(n_168), .B(n_185), .Y(n_354) );
AO31x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_178), .A3(n_179), .B(n_180), .Y(n_168) );
OAI22x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B1(n_174), .B2(n_176), .Y(n_169) );
INVx4_ASAP7_75t_L g172 ( .A(n_171), .Y(n_172) );
INVx1_ASAP7_75t_L g521 ( .A(n_171), .Y(n_521) );
INVx1_ASAP7_75t_L g537 ( .A(n_171), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_172), .A2(n_229), .B(n_230), .C(n_231), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_173), .A2(n_176), .B1(n_267), .B2(n_269), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_173), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_173), .A2(n_176), .B1(n_511), .B2(n_513), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_173), .A2(n_519), .B1(n_522), .B2(n_523), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_173), .A2(n_503), .B1(n_535), .B2(n_536), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_173), .A2(n_503), .B1(n_544), .B2(n_546), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_173), .A2(n_503), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_173), .A2(n_523), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_173), .A2(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_175), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g270 ( .A(n_175), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_176), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_SL g523 ( .A(n_177), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_178), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_178), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g199 ( .A(n_179), .Y(n_199) );
AO31x2_ASAP7_75t_L g500 ( .A1(n_179), .A2(n_260), .A3(n_501), .B(n_505), .Y(n_500) );
AO31x2_ASAP7_75t_L g542 ( .A1(n_179), .A2(n_509), .A3(n_543), .B(n_548), .Y(n_542) );
AO31x2_ASAP7_75t_L g562 ( .A1(n_179), .A2(n_241), .A3(n_563), .B(n_567), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx2_ASAP7_75t_L g201 ( .A(n_182), .Y(n_201) );
BUFx2_ASAP7_75t_L g241 ( .A(n_182), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_182), .B(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_182), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_184), .B(n_353), .Y(n_396) );
OR2x2_ASAP7_75t_L g484 ( .A(n_184), .B(n_345), .Y(n_484) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g312 ( .A(n_185), .Y(n_312) );
AND2x2_ASAP7_75t_L g321 ( .A(n_185), .B(n_284), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_185), .B(n_225), .Y(n_324) );
AND2x2_ASAP7_75t_L g343 ( .A(n_185), .B(n_224), .Y(n_343) );
AND2x4_ASAP7_75t_L g362 ( .A(n_185), .B(n_285), .Y(n_362) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_189), .B(n_200), .Y(n_185) );
AO31x2_ASAP7_75t_L g533 ( .A1(n_186), .A2(n_524), .A3(n_534), .B(n_538), .Y(n_533) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_186), .A2(n_272), .A3(n_553), .B(n_556), .Y(n_552) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_188), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_SL g567 ( .A(n_188), .B(n_568), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_193), .B(n_199), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
INVx2_ASAP7_75t_L g268 ( .A(n_196), .Y(n_268) );
INVx1_ASAP7_75t_L g545 ( .A(n_196), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_197), .Y(n_547) );
INVx1_ASAP7_75t_L g524 ( .A(n_199), .Y(n_524) );
OAI21xp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_222), .B(n_263), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_203), .B(n_357), .Y(n_460) );
CKINVDCx14_ASAP7_75t_R g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_205), .B(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g293 ( .A(n_205), .Y(n_293) );
OR2x2_ASAP7_75t_L g301 ( .A(n_205), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_205), .B(n_294), .Y(n_326) );
AND2x2_ASAP7_75t_L g351 ( .A(n_205), .B(n_265), .Y(n_351) );
AND2x2_ASAP7_75t_L g369 ( .A(n_205), .B(n_299), .Y(n_369) );
INVx1_ASAP7_75t_L g408 ( .A(n_205), .Y(n_408) );
AND2x2_ASAP7_75t_L g410 ( .A(n_205), .B(n_411), .Y(n_410) );
NAND2x1p5_ASAP7_75t_SL g429 ( .A(n_205), .B(n_350), .Y(n_429) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_209), .Y(n_205) );
NOR2x1_ASAP7_75t_L g236 ( .A(n_207), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g220 ( .A(n_208), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_208), .B(n_506), .Y(n_505) );
BUFx3_ASAP7_75t_L g509 ( .A(n_208), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_208), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_208), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_SL g577 ( .A(n_208), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_216), .B(n_220), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_219), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g237 ( .A(n_221), .Y(n_237) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_221), .A2(n_257), .A3(n_260), .B(n_261), .Y(n_256) );
OAI32xp33_ASAP7_75t_L g313 ( .A1(n_222), .A2(n_305), .A3(n_314), .B1(n_316), .B2(n_318), .Y(n_313) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_238), .Y(n_222) );
INVx1_ASAP7_75t_L g353 ( .A(n_223), .Y(n_353) );
AND2x2_ASAP7_75t_L g361 ( .A(n_223), .B(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g360 ( .A(n_224), .B(n_284), .Y(n_360) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx3_ASAP7_75t_L g310 ( .A(n_225), .Y(n_310) );
AND2x2_ASAP7_75t_L g319 ( .A(n_225), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g425 ( .A(n_225), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_233), .B(n_236), .Y(n_227) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
OR2x2_ASAP7_75t_L g305 ( .A(n_238), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g427 ( .A(n_238), .Y(n_427) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_255), .Y(n_238) );
AND2x2_ASAP7_75t_L g328 ( .A(n_239), .B(n_256), .Y(n_328) );
INVx2_ASAP7_75t_L g350 ( .A(n_239), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_239), .B(n_265), .Y(n_370) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g277 ( .A(n_240), .Y(n_277) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_254), .Y(n_240) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_241), .A2(n_266), .A3(n_272), .B(n_274), .Y(n_265) );
AO31x2_ASAP7_75t_L g517 ( .A1(n_241), .A2(n_518), .A3(n_524), .B(n_525), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_246), .B(n_249), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g271 ( .A(n_247), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_SL g512 ( .A(n_253), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_255), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g359 ( .A(n_255), .Y(n_359) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
BUFx2_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
OR2x2_ASAP7_75t_L g365 ( .A(n_256), .B(n_265), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_256), .B(n_265), .Y(n_398) );
INVx2_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_276), .Y(n_263) );
OR2x2_ASAP7_75t_L g333 ( .A(n_264), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g411 ( .A(n_264), .Y(n_411) );
INVx1_ASAP7_75t_L g294 ( .A(n_265), .Y(n_294) );
INVx1_ASAP7_75t_L g302 ( .A(n_265), .Y(n_302) );
INVx1_ASAP7_75t_L g317 ( .A(n_265), .Y(n_317) );
AO31x2_ASAP7_75t_L g508 ( .A1(n_272), .A2(n_509), .A3(n_510), .B(n_514), .Y(n_508) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_SL g585 ( .A(n_273), .Y(n_585) );
OR2x2_ASAP7_75t_L g421 ( .A(n_276), .B(n_398), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_277), .B(n_293), .Y(n_334) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_277), .Y(n_336) );
OR2x2_ASAP7_75t_L g435 ( .A(n_277), .B(n_359), .Y(n_435) );
INVxp67_ASAP7_75t_L g459 ( .A(n_277), .Y(n_459) );
INVx2_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NAND2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_280), .B(n_321), .Y(n_388) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g337 ( .A(n_282), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g450 ( .A(n_283), .Y(n_450) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g479 ( .A(n_284), .B(n_312), .Y(n_479) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g405 ( .A(n_285), .B(n_312), .Y(n_405) );
AOI21x1_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_292), .B(n_328), .Y(n_442) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g306 ( .A(n_293), .Y(n_306) );
AND2x2_ASAP7_75t_L g356 ( .A(n_293), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_293), .B(n_350), .Y(n_399) );
OR2x2_ASAP7_75t_L g471 ( .A(n_293), .B(n_358), .Y(n_471) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g391 ( .A(n_297), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx2_ASAP7_75t_L g382 ( .A(n_298), .Y(n_382) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g372 ( .A(n_301), .B(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_301), .Y(n_383) );
OR2x2_ASAP7_75t_L g434 ( .A(n_301), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g489 ( .A(n_301), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B(n_313), .C(n_322), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g378 ( .A(n_306), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_306), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g451 ( .A(n_306), .B(n_328), .Y(n_451) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_309), .B(n_354), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_309), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g461 ( .A(n_309), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g404 ( .A(n_310), .Y(n_404) );
AND2x2_ASAP7_75t_L g432 ( .A(n_311), .B(n_360), .Y(n_432) );
INVx2_ASAP7_75t_L g455 ( .A(n_311), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_311), .B(n_353), .Y(n_487) );
AND2x4_ASAP7_75t_SL g441 ( .A(n_314), .B(n_319), .Y(n_441) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g394 ( .A(n_315), .B(n_320), .Y(n_394) );
OR2x2_ASAP7_75t_L g446 ( .A(n_315), .B(n_339), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_316), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_316), .B(n_328), .Y(n_482) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g430 ( .A(n_317), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g413 ( .A(n_319), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_319), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g463 ( .A(n_320), .Y(n_463) );
BUFx2_ASAP7_75t_L g331 ( .A(n_321), .Y(n_331) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g449 ( .A(n_324), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_328), .Y(n_390) );
NAND3xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_340), .C(n_355), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_332), .B1(n_335), .B2(n_337), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_337), .A2(n_363), .B1(n_444), .B2(n_447), .C1(n_449), .C2(n_451), .Y(n_443) );
AND2x2_ASAP7_75t_L g475 ( .A(n_338), .B(n_424), .Y(n_475) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g423 ( .A(n_339), .B(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_346), .B1(n_347), .B2(n_352), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_SL g419 ( .A(n_343), .Y(n_419) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
AND2x2_ASAP7_75t_L g406 ( .A(n_348), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g364 ( .A(n_349), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g358 ( .A(n_350), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g473 ( .A(n_351), .Y(n_473) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_354), .B(n_450), .Y(n_469) );
INVx1_ASAP7_75t_L g486 ( .A(n_354), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B1(n_361), .B2(n_363), .C1(n_366), .C2(n_367), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_362), .Y(n_366) );
AND2x2_ASAP7_75t_L g384 ( .A(n_362), .B(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g379 ( .A(n_365), .Y(n_379) );
OR2x2_ASAP7_75t_L g448 ( .A(n_365), .B(n_429), .Y(n_448) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B(n_377), .C(n_386), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI21xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_384), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_378), .A2(n_416), .B1(n_465), .B2(n_468), .C(n_470), .Y(n_464) );
AND2x4_ASAP7_75t_L g407 ( .A(n_379), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
AOI211x1_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_391), .C(n_395), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g456 ( .A(n_394), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_397), .B(n_445), .C(n_446), .Y(n_444) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g480 ( .A(n_398), .Y(n_480) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_452), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_409), .C(n_431), .D(n_443), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g462 ( .A(n_405), .B(n_463), .Y(n_462) );
AOI221x1_ASAP7_75t_L g431 ( .A1(n_407), .A2(n_432), .B1(n_433), .B2(n_436), .C(n_439), .Y(n_431) );
AND2x2_ASAP7_75t_L g457 ( .A(n_407), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_416), .B2(n_420), .C(n_422), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_414), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_419), .A2(n_423), .B1(n_426), .B2(n_428), .Y(n_422) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_423), .A2(n_440), .B(n_442), .Y(n_439) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g445 ( .A(n_425), .Y(n_445) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g466 ( .A(n_435), .Y(n_466) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_448), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_464), .C(n_476), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B1(n_460), .B2(n_461), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g472 ( .A(n_459), .B(n_473), .Y(n_472) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_459), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_474), .Y(n_470) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_480), .B1(n_481), .B2(n_483), .C(n_485), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g795 ( .A(n_490), .Y(n_795) );
BUFx12f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g826 ( .A(n_492), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g813 ( .A(n_493), .Y(n_813) );
NOR2x1p5_ASAP7_75t_L g493 ( .A(n_494), .B(n_705), .Y(n_493) );
NAND4xp75_ASAP7_75t_L g494 ( .A(n_495), .B(n_650), .C(n_670), .D(n_686), .Y(n_494) );
NOR2x1p5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_620), .Y(n_495) );
NAND4xp75_ASAP7_75t_L g496 ( .A(n_497), .B(n_558), .C(n_597), .D(n_606), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_527), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_507), .Y(n_498) );
AND2x4_ASAP7_75t_L g730 ( .A(n_499), .B(n_657), .Y(n_730) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
INVx2_ASAP7_75t_L g591 ( .A(n_500), .Y(n_591) );
AND2x2_ASAP7_75t_L g614 ( .A(n_500), .B(n_576), .Y(n_614) );
OR2x2_ASAP7_75t_L g669 ( .A(n_500), .B(n_508), .Y(n_669) );
AND2x2_ASAP7_75t_L g587 ( .A(n_507), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g737 ( .A(n_507), .B(n_614), .Y(n_737) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
OR2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g605 ( .A(n_508), .Y(n_605) );
AND2x2_ASAP7_75t_L g611 ( .A(n_508), .B(n_517), .Y(n_611) );
INVx1_ASAP7_75t_L g629 ( .A(n_508), .Y(n_629) );
INVx2_ASAP7_75t_L g658 ( .A(n_508), .Y(n_658) );
INVx3_ASAP7_75t_L g634 ( .A(n_516), .Y(n_634) );
INVx2_ASAP7_75t_L g639 ( .A(n_516), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_516), .B(n_590), .Y(n_644) );
AND2x2_ASAP7_75t_L g667 ( .A(n_516), .B(n_646), .Y(n_667) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_516), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_516), .B(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g656 ( .A(n_517), .Y(n_656) );
AND2x2_ASAP7_75t_L g704 ( .A(n_517), .B(n_658), .Y(n_704) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_529), .B(n_648), .Y(n_695) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g692 ( .A(n_530), .B(n_648), .Y(n_692) );
INVx1_ASAP7_75t_L g793 ( .A(n_530), .Y(n_793) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g743 ( .A(n_531), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g596 ( .A(n_532), .Y(n_596) );
OR2x2_ASAP7_75t_L g677 ( .A(n_532), .B(n_551), .Y(n_677) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g619 ( .A(n_533), .Y(n_619) );
AND2x4_ASAP7_75t_L g625 ( .A(n_533), .B(n_626), .Y(n_625) );
AOI32xp33_ASAP7_75t_L g763 ( .A1(n_540), .A2(n_666), .A3(n_764), .B1(n_766), .B2(n_767), .Y(n_763) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g712 ( .A(n_541), .B(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_550), .Y(n_541) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_542), .Y(n_560) );
OR2x2_ASAP7_75t_L g594 ( .A(n_542), .B(n_552), .Y(n_594) );
INVx1_ASAP7_75t_L g609 ( .A(n_542), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_542), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g624 ( .A(n_542), .Y(n_624) );
INVx2_ASAP7_75t_L g649 ( .A(n_542), .Y(n_649) );
AND2x2_ASAP7_75t_L g768 ( .A(n_542), .B(n_562), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_550), .B(n_601), .Y(n_688) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g561 ( .A(n_552), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g617 ( .A(n_552), .Y(n_617) );
INVx2_ASAP7_75t_L g626 ( .A(n_552), .Y(n_626) );
AND2x4_ASAP7_75t_L g648 ( .A(n_552), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_552), .Y(n_740) );
AOI22x1_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_569), .B1(n_587), .B2(n_592), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_561), .B(n_718), .C(n_719), .D(n_720), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_561), .B(n_618), .Y(n_748) );
INVx4_ASAP7_75t_SL g601 ( .A(n_562), .Y(n_601) );
BUFx2_ASAP7_75t_L g664 ( .A(n_562), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_562), .B(n_609), .Y(n_727) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g689 ( .A(n_571), .B(n_638), .Y(n_689) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g612 ( .A(n_575), .B(n_590), .Y(n_612) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_576), .B(n_591), .Y(n_636) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_586), .Y(n_576) );
OAI21x1_ASAP7_75t_L g631 ( .A1(n_577), .A2(n_578), .B(n_586), .Y(n_631) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B(n_585), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_588), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g654 ( .A(n_588), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g693 ( .A(n_589), .B(n_611), .Y(n_693) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g736 ( .A(n_591), .B(n_646), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_592), .A2(n_709), .B1(n_711), .B2(n_714), .C(n_716), .Y(n_708) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g602 ( .A(n_594), .Y(n_602) );
OR2x2_ASAP7_75t_L g702 ( .A(n_594), .B(n_641), .Y(n_702) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_603), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_598), .A2(n_724), .B1(n_728), .B2(n_731), .Y(n_723) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
AND2x4_ASAP7_75t_L g647 ( .A(n_599), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g759 ( .A(n_599), .B(n_677), .Y(n_759) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g607 ( .A(n_601), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g623 ( .A(n_601), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g682 ( .A(n_601), .B(n_619), .Y(n_682) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_601), .Y(n_699) );
INVx1_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_601), .B(n_626), .Y(n_756) );
AND2x4_ASAP7_75t_L g663 ( .A(n_602), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g661 ( .A(n_604), .Y(n_661) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_605), .B(n_646), .Y(n_645) );
NAND2x1_ASAP7_75t_L g765 ( .A(n_605), .B(n_667), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_610), .B1(n_613), .B2(n_615), .Y(n_606) );
AND2x2_ASAP7_75t_L g632 ( .A(n_607), .B(n_625), .Y(n_632) );
INVx1_ASAP7_75t_L g673 ( .A(n_607), .Y(n_673) );
AND2x2_ASAP7_75t_L g780 ( .A(n_607), .B(n_641), .Y(n_780) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g613 ( .A(n_611), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g753 ( .A(n_611), .Y(n_753) );
AND2x2_ASAP7_75t_L g770 ( .A(n_611), .B(n_630), .Y(n_770) );
AND2x2_ASAP7_75t_L g786 ( .A(n_611), .B(n_736), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_612), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g709 ( .A(n_612), .B(n_710), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_612), .A2(n_702), .B1(n_717), .B2(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g672 ( .A(n_614), .Y(n_672) );
AND2x2_ASAP7_75t_L g703 ( .A(n_614), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_614), .B(n_710), .Y(n_732) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g738 ( .A(n_618), .B(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_618), .A2(n_642), .B1(n_747), .B2(n_749), .Y(n_746) );
INVx3_ASAP7_75t_L g641 ( .A(n_619), .Y(n_641) );
AND2x2_ASAP7_75t_L g773 ( .A(n_619), .B(n_626), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_637), .Y(n_620) );
AOI32xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_627), .A3(n_630), .B1(n_632), .B2(n_633), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_624), .Y(n_719) );
INVx1_ASAP7_75t_L g744 ( .A(n_624), .Y(n_744) );
INVx3_ASAP7_75t_L g700 ( .A(n_625), .Y(n_700) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_628), .A2(n_776), .B1(n_777), .B2(n_778), .C(n_779), .Y(n_775) );
BUFx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g752 ( .A(n_630), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g788 ( .A(n_630), .B(n_749), .Y(n_788) );
BUFx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g646 ( .A(n_631), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_633), .B(n_661), .Y(n_660) );
AO22x1_ASAP7_75t_L g690 ( .A1(n_633), .A2(n_691), .B1(n_693), .B2(n_694), .Y(n_690) );
NAND2x1p5_ASAP7_75t_L g794 ( .A(n_633), .B(n_661), .Y(n_794) );
AND2x4_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g710 ( .A(n_634), .Y(n_710) );
INVx1_ASAP7_75t_L g720 ( .A(n_634), .Y(n_720) );
AND2x2_ASAP7_75t_L g640 ( .A(n_635), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_636), .Y(n_722) );
INVx1_ASAP7_75t_L g762 ( .A(n_636), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_642), .C(n_647), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2x1p5_ASAP7_75t_L g749 ( .A(n_639), .B(n_669), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_640), .B(n_699), .Y(n_776) );
AOI31xp33_ASAP7_75t_L g659 ( .A1(n_641), .A2(n_660), .A3(n_662), .B(n_665), .Y(n_659) );
INVx4_ASAP7_75t_L g718 ( .A(n_641), .Y(n_718) );
OR2x2_ASAP7_75t_L g755 ( .A(n_641), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AND2x4_ASAP7_75t_L g657 ( .A(n_646), .B(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_648), .Y(n_653) );
AND2x2_ASAP7_75t_L g684 ( .A(n_648), .B(n_682), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g650 ( .A(n_651), .B(n_659), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g777 ( .A(n_654), .Y(n_777) );
INVx1_ASAP7_75t_L g685 ( .A(n_655), .Y(n_685) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g715 ( .A(n_656), .Y(n_715) );
AND2x2_ASAP7_75t_L g714 ( .A(n_657), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI322xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .A3(n_674), .B1(n_678), .B2(n_681), .C1(n_683), .C2(n_685), .Y(n_671) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI211x1_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_690), .C(n_696), .Y(n_686) );
INVx1_ASAP7_75t_L g791 ( .A(n_687), .Y(n_791) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g745 ( .A(n_689), .Y(n_745) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OA21x2_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_701), .B(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g766 ( .A(n_700), .Y(n_766) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp33_ASAP7_75t_L g761 ( .A(n_704), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_774), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_741), .C(n_757), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_723), .C(n_733), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_710), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_714), .A2(n_770), .B(n_771), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_718), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_718), .B(n_768), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_719), .B(n_793), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_720), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_730), .A2(n_780), .B(n_781), .Y(n_779) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_737), .B(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B(n_746), .C(n_750), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_SL g760 ( .A(n_752), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_756), .Y(n_778) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_763), .C(n_769), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_768), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g789 ( .A(n_768), .Y(n_789) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g785 ( .A(n_773), .Y(n_785) );
NOR3xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_783), .C(n_790), .Y(n_774) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI21xp33_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_787), .B(n_789), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI21xp33_ASAP7_75t_R g790 ( .A1(n_791), .A2(n_792), .B(n_794), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_798), .A2(n_811), .B(n_815), .Y(n_810) );
INVxp67_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
BUFx12f_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx4_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AO21x1_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_810), .B(n_820), .Y(n_806) );
CKINVDCx11_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx3_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx4_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
BUFx10_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
endmodule