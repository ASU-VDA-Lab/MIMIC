module fake_netlist_1_7568_n_1366 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1366);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1366;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g322 ( .A(n_64), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_233), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_312), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_74), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_98), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_39), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_49), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_106), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_1), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_28), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_109), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_172), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_314), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_78), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_250), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_204), .Y(n_341) );
INVxp33_ASAP7_75t_L g342 ( .A(n_5), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_111), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_112), .Y(n_344) );
CKINVDCx14_ASAP7_75t_R g345 ( .A(n_131), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_82), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_231), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_23), .Y(n_348) );
CKINVDCx16_ASAP7_75t_R g349 ( .A(n_241), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_46), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_310), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_202), .Y(n_352) );
CKINVDCx14_ASAP7_75t_R g353 ( .A(n_113), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_277), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_299), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_47), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_22), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_189), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_169), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_83), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_155), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_196), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_88), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_89), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_35), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_2), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_313), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_236), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_207), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_66), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_176), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_285), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_53), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_55), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_301), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_263), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_218), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_173), .B(n_211), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_84), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_121), .B(n_146), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_297), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_276), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_280), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_77), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_264), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_52), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_41), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_97), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_281), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_286), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_287), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_254), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_188), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_150), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_247), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_291), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_65), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_116), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_99), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_158), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_37), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_129), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_78), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g404 ( .A(n_115), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_283), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_62), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_137), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_295), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_193), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_48), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_147), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_31), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_309), .Y(n_413) );
INVxp33_ASAP7_75t_SL g414 ( .A(n_140), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_65), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_187), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_25), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_95), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_302), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_235), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_167), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_262), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_74), .Y(n_423) );
INVxp33_ASAP7_75t_SL g424 ( .A(n_132), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_256), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_186), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_265), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_33), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_108), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_138), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_39), .Y(n_431) );
INVxp33_ASAP7_75t_L g432 ( .A(n_305), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_107), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_163), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_308), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_56), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_136), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_245), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_240), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_49), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_55), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_157), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_296), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_252), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_177), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_92), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_242), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_260), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_184), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_52), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_134), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_3), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_45), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_50), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_34), .Y(n_455) );
INVxp33_ASAP7_75t_SL g456 ( .A(n_54), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_77), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_273), .Y(n_458) );
BUFx5_ASAP7_75t_L g459 ( .A(n_237), .Y(n_459) );
BUFx10_ASAP7_75t_L g460 ( .A(n_289), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_12), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_127), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_20), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_318), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_105), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_320), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_300), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_30), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_63), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_215), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_94), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_311), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_269), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_292), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_144), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_53), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_174), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_208), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_165), .Y(n_479) );
INVxp33_ASAP7_75t_SL g480 ( .A(n_234), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_154), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_122), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_183), .Y(n_483) );
BUFx2_ASAP7_75t_SL g484 ( .A(n_274), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_319), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_206), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_68), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_15), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_275), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_342), .B(n_0), .Y(n_490) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_348), .B(n_0), .Y(n_491) );
NAND2xp33_ASAP7_75t_L g492 ( .A(n_459), .B(n_432), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_346), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_457), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_356), .B(n_1), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_342), .Y(n_498) );
INVx6_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_346), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_482), .B(n_2), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_363), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_432), .B(n_3), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_423), .B(n_4), .Y(n_504) );
BUFx12f_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_363), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_365), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_348), .B(n_4), .Y(n_508) );
AND2x6_ASAP7_75t_L g509 ( .A(n_396), .B(n_90), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_337), .B(n_5), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_386), .Y(n_511) );
OAI22x1_ASAP7_75t_L g512 ( .A1(n_386), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_512) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_324), .A2(n_93), .B(n_91), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_460), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_323), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_409), .B(n_6), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_360), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_323), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_397), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_350), .B(n_7), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_411), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_329), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_466), .B(n_8), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_323), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_350), .B(n_9), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_323), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_441), .B(n_9), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_478), .B(n_10), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_493), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_514), .B(n_335), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_508), .A2(n_327), .B1(n_328), .B2(n_322), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_515), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_498), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_493), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_515), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_515), .Y(n_539) );
BUFx3_ASAP7_75t_L g540 ( .A(n_509), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_515), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_495), .B(n_454), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_514), .B(n_354), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_515), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_517), .B(n_345), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_508), .B(n_324), .Y(n_546) );
INVx4_ASAP7_75t_L g547 ( .A(n_509), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_517), .B(n_345), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_508), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_514), .B(n_425), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_495), .B(n_461), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_493), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_508), .B(n_333), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_496), .Y(n_554) );
INVx4_ASAP7_75t_L g555 ( .A(n_509), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_496), .Y(n_556) );
NOR3xp33_ASAP7_75t_L g557 ( .A(n_490), .B(n_469), .C(n_373), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_496), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_490), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_518), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_518), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_490), .B(n_353), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
AND2x6_ASAP7_75t_L g565 ( .A(n_521), .B(n_396), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_514), .B(n_458), .Y(n_566) );
BUFx10_ASAP7_75t_L g567 ( .A(n_499), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_518), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_521), .B(n_333), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_516), .B(n_331), .C(n_374), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_521), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_503), .Y(n_573) );
INVx3_ASAP7_75t_L g574 ( .A(n_521), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_499), .B(n_470), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_518), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_503), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_518), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_526), .B(n_441), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_526), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_560), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_573), .B(n_499), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_573), .B(n_499), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_577), .B(n_499), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g585 ( .A1(n_560), .A2(n_512), .B1(n_524), .B2(n_516), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_577), .B(n_522), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_557), .A2(n_529), .B1(n_510), .B2(n_492), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_563), .B(n_505), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_557), .A2(n_529), .B1(n_510), .B2(n_522), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_563), .B(n_522), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_545), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_535), .B(n_523), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_550), .B(n_505), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_545), .B(n_510), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_547), .B(n_526), .Y(n_597) );
OR2x6_ASAP7_75t_L g598 ( .A(n_542), .B(n_505), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_547), .B(n_526), .Y(n_599) );
NOR2x1p5_ASAP7_75t_L g600 ( .A(n_542), .B(n_523), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_579), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_545), .B(n_349), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_548), .B(n_529), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_532), .B(n_524), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_549), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_579), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_579), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_579), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_536), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
OAI22xp5_ASAP7_75t_SL g611 ( .A1(n_542), .A2(n_357), .B1(n_507), .B2(n_456), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_536), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_550), .B(n_497), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_540), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_566), .B(n_497), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_565), .A2(n_528), .B1(n_509), .B2(n_512), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_532), .B(n_528), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_548), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_548), .B(n_355), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_535), .B(n_528), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_572), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_572), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_572), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_572), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_551), .Y(n_625) );
AND2x6_ASAP7_75t_SL g626 ( .A(n_543), .B(n_504), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_547), .B(n_528), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_551), .A2(n_357), .B1(n_456), .B2(n_402), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_574), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_533), .B(n_421), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g631 ( .A(n_551), .B(n_566), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_574), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_547), .B(n_462), .Y(n_633) );
CKINVDCx11_ASAP7_75t_R g634 ( .A(n_567), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_565), .A2(n_509), .B1(n_512), .B2(n_494), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_574), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_574), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_571), .B(n_504), .Y(n_639) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_533), .B(n_479), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_547), .B(n_486), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_543), .B(n_501), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_565), .A2(n_509), .B1(n_494), .B2(n_502), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_580), .Y(n_644) );
AO22x1_ASAP7_75t_L g645 ( .A1(n_565), .A2(n_424), .B1(n_480), .B2(n_414), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_565), .A2(n_509), .B1(n_500), .B2(n_506), .Y(n_646) );
NAND2xp33_ASAP7_75t_L g647 ( .A(n_565), .B(n_459), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_540), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_555), .B(n_368), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_555), .B(n_368), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_555), .B(n_375), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_580), .Y(n_652) );
INVx8_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_575), .B(n_472), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_565), .A2(n_500), .B1(n_506), .B2(n_502), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_580), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_575), .B(n_375), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_546), .B(n_414), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_553), .B(n_424), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_567), .Y(n_660) );
AO22x1_ASAP7_75t_L g661 ( .A1(n_565), .A2(n_480), .B1(n_364), .B2(n_417), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_555), .B(n_422), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_SL g663 ( .A1(n_580), .A2(n_353), .B(n_442), .C(n_404), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_580), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_565), .Y(n_665) );
NAND2xp33_ASAP7_75t_L g666 ( .A(n_571), .B(n_459), .Y(n_666) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_555), .B(n_491), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_553), .B(n_511), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_567), .B(n_364), .Y(n_669) );
BUFx3_ASAP7_75t_L g670 ( .A(n_567), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_570), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_531), .B(n_387), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_537), .B(n_422), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_537), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_613), .B(n_552), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_631), .B(n_387), .Y(n_676) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_618), .B(n_540), .Y(n_677) );
INVx3_ASAP7_75t_SL g678 ( .A(n_598), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_598), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_601), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_589), .B(n_402), .C(n_394), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_613), .B(n_552), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_660), .B(n_439), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_592), .B(n_417), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_625), .B(n_394), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_634), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_639), .B(n_413), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_597), .A2(n_556), .B(n_554), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_656), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_595), .B(n_413), .Y(n_690) );
NOR2xp67_ASAP7_75t_L g691 ( .A(n_595), .B(n_453), .Y(n_691) );
AND2x6_ASAP7_75t_L g692 ( .A(n_653), .B(n_491), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_585), .A2(n_416), .B1(n_437), .B2(n_554), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_666), .B(n_513), .C(n_556), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_597), .A2(n_559), .B(n_558), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_615), .B(n_558), .Y(n_696) );
AOI22x1_ASAP7_75t_L g697 ( .A1(n_667), .A2(n_564), .B1(n_568), .B2(n_559), .Y(n_697) );
BUFx3_ASAP7_75t_L g698 ( .A(n_598), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_615), .B(n_564), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_626), .B(n_416), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_602), .B(n_437), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_604), .B(n_568), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_669), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_596), .B(n_453), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_599), .A2(n_513), .B(n_332), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_619), .B(n_325), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_593), .B(n_436), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_609), .B(n_330), .Y(n_708) );
INVx4_ASAP7_75t_L g709 ( .A(n_653), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_642), .A2(n_463), .B(n_366), .C(n_370), .Y(n_710) );
NOR2xp67_ASAP7_75t_L g711 ( .A(n_587), .B(n_586), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_591), .B(n_384), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_596), .B(n_403), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_599), .A2(n_513), .B(n_334), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_603), .B(n_468), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_611), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_603), .B(n_379), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_620), .B(n_487), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_670), .B(n_439), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_620), .B(n_449), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_628), .B(n_401), .C(n_339), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_585), .A2(n_442), .B1(n_404), .B2(n_410), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_642), .A2(n_463), .B(n_406), .C(n_431), .Y(n_723) );
NOR2xp67_ASAP7_75t_L g724 ( .A(n_616), .B(n_489), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_600), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_612), .B(n_672), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_617), .A2(n_428), .B(n_452), .C(n_450), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_654), .B(n_489), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_661), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_606), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_627), .A2(n_513), .B(n_340), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_581), .B(n_455), .Y(n_732) );
O2A1O1Ixp33_ASAP7_75t_L g733 ( .A1(n_590), .A2(n_476), .B(n_440), .C(n_397), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_667), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_630), .B(n_511), .Y(n_735) );
BUFx12f_ASAP7_75t_L g736 ( .A(n_630), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_SL g737 ( .A1(n_654), .A2(n_380), .B(n_519), .C(n_338), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_607), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_582), .B(n_519), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_583), .B(n_440), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_588), .B(n_658), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_658), .B(n_351), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_621), .A2(n_341), .B(n_326), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_608), .Y(n_744) );
O2A1O1Ixp5_ASAP7_75t_SL g745 ( .A1(n_633), .A2(n_344), .B(n_347), .C(n_343), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_656), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_640), .A2(n_488), .B1(n_415), .B2(n_412), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_659), .B(n_465), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_584), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_665), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_671), .A2(n_488), .B(n_358), .C(n_361), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_640), .A2(n_415), .B1(n_412), .B2(n_362), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_645), .B(n_474), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_657), .B(n_484), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_655), .B(n_359), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_594), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_623), .Y(n_757) );
INVx4_ASAP7_75t_L g758 ( .A(n_653), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_616), .A2(n_369), .B1(n_372), .B2(n_367), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_665), .B(n_376), .Y(n_760) );
BUFx12f_ASAP7_75t_L g761 ( .A(n_614), .Y(n_761) );
AOI21x1_ASAP7_75t_L g762 ( .A1(n_633), .A2(n_534), .B(n_530), .Y(n_762) );
BUFx2_ASAP7_75t_L g763 ( .A(n_673), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_674), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_668), .A2(n_415), .B1(n_412), .B2(n_383), .C(n_385), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_624), .A2(n_382), .B(n_377), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_605), .Y(n_767) );
BUFx5_ASAP7_75t_L g768 ( .A(n_632), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_671), .B(n_412), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_610), .Y(n_770) );
AND2x4_ASAP7_75t_L g771 ( .A(n_636), .B(n_388), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_635), .A2(n_390), .B1(n_391), .B2(n_389), .Y(n_772) );
OA22x2_ASAP7_75t_L g773 ( .A1(n_641), .A2(n_395), .B1(n_399), .B2(n_393), .Y(n_773) );
O2A1O1Ixp33_ASAP7_75t_L g774 ( .A1(n_668), .A2(n_407), .B(n_408), .C(n_400), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_637), .A2(n_426), .B(n_418), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_SL g776 ( .A1(n_643), .A2(n_380), .B(n_534), .C(n_530), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_644), .A2(n_430), .B(n_429), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_664), .B(n_433), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_622), .A2(n_438), .B(n_434), .Y(n_779) );
OR2x2_ASAP7_75t_L g780 ( .A(n_655), .B(n_635), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_629), .A2(n_445), .B(n_444), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_652), .A2(n_447), .B1(n_448), .B2(n_446), .Y(n_782) );
BUFx3_ASAP7_75t_L g783 ( .A(n_614), .Y(n_783) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_614), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_647), .B(n_451), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_649), .B(n_467), .Y(n_786) );
NOR2x1_ASAP7_75t_SL g787 ( .A(n_650), .B(n_419), .Y(n_787) );
BUFx3_ASAP7_75t_L g788 ( .A(n_614), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_651), .A2(n_662), .B(n_648), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_638), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_646), .A2(n_473), .B1(n_475), .B2(n_471), .Y(n_791) );
INVxp67_ASAP7_75t_L g792 ( .A(n_646), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_638), .A2(n_481), .B1(n_483), .B2(n_477), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_638), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_638), .B(n_485), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_648), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_648), .B(n_419), .Y(n_797) );
INVx4_ASAP7_75t_L g798 ( .A(n_648), .Y(n_798) );
AOI21x1_ASAP7_75t_L g799 ( .A1(n_663), .A2(n_534), .B(n_530), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g800 ( .A(n_663), .B(n_352), .Y(n_800) );
INVx4_ASAP7_75t_L g801 ( .A(n_634), .Y(n_801) );
O2A1O1Ixp33_ASAP7_75t_L g802 ( .A1(n_585), .A2(n_371), .B(n_381), .C(n_352), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_630), .A2(n_371), .B1(n_392), .B2(n_381), .Y(n_803) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_660), .B(n_392), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_601), .Y(n_805) );
INVx3_ASAP7_75t_SL g806 ( .A(n_598), .Y(n_806) );
O2A1O1Ixp33_ASAP7_75t_L g807 ( .A1(n_585), .A2(n_420), .B(n_443), .C(n_435), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_598), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_597), .A2(n_435), .B(n_420), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_SL g810 ( .A1(n_642), .A2(n_539), .B(n_541), .C(n_538), .Y(n_810) );
NAND2xp33_ASAP7_75t_SL g811 ( .A(n_665), .B(n_443), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_L g812 ( .A1(n_585), .A2(n_464), .B(n_427), .C(n_378), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_601), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_625), .B(n_10), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_625), .B(n_11), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_601), .Y(n_816) );
A2O1A1Ixp33_ASAP7_75t_L g817 ( .A1(n_613), .A2(n_464), .B(n_427), .C(n_398), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_631), .B(n_11), .Y(n_818) );
INVxp67_ASAP7_75t_L g819 ( .A(n_592), .Y(n_819) );
NOR2x1_ASAP7_75t_L g820 ( .A(n_598), .B(n_336), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_631), .B(n_12), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_597), .A2(n_539), .B(n_538), .Y(n_822) );
NOR2xp33_ASAP7_75t_SL g823 ( .A(n_801), .B(n_336), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_705), .A2(n_578), .B(n_544), .Y(n_824) );
AND2x4_ASAP7_75t_L g825 ( .A(n_734), .B(n_13), .Y(n_825) );
INVx8_ASAP7_75t_L g826 ( .A(n_808), .Y(n_826) );
INVx1_ASAP7_75t_SL g827 ( .A(n_678), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_684), .B(n_13), .Y(n_828) );
O2A1O1Ixp33_ASAP7_75t_SL g829 ( .A1(n_776), .A2(n_737), .B(n_810), .C(n_817), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_747), .A2(n_405), .B1(n_398), .B2(n_518), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_711), .B(n_14), .Y(n_831) );
INVx3_ASAP7_75t_L g832 ( .A(n_801), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_L g833 ( .A1(n_710), .A2(n_544), .B(n_561), .C(n_541), .Y(n_833) );
INVxp67_ASAP7_75t_L g834 ( .A(n_685), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_747), .A2(n_405), .B1(n_527), .B2(n_525), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_698), .B(n_14), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_714), .A2(n_578), .B(n_562), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_721), .A2(n_405), .B1(n_525), .B2(n_527), .C(n_578), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_735), .B(n_15), .Y(n_839) );
A2O1A1Ixp33_ASAP7_75t_L g840 ( .A1(n_812), .A2(n_527), .B(n_525), .C(n_561), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_790), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_731), .A2(n_562), .B(n_561), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_702), .A2(n_576), .B(n_569), .Y(n_843) );
OR2x2_ASAP7_75t_L g844 ( .A(n_819), .B(n_16), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_764), .Y(n_845) );
CKINVDCx6p67_ASAP7_75t_R g846 ( .A(n_686), .Y(n_846) );
O2A1O1Ixp33_ASAP7_75t_SL g847 ( .A1(n_723), .A2(n_569), .B(n_576), .C(n_562), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_679), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_761), .Y(n_849) );
BUFx3_ASAP7_75t_L g850 ( .A(n_725), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_726), .B(n_16), .Y(n_851) );
INVx2_ASAP7_75t_SL g852 ( .A(n_820), .Y(n_852) );
NOR2xp33_ASAP7_75t_SL g853 ( .A(n_709), .B(n_525), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_694), .A2(n_527), .B(n_100), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_687), .B(n_17), .Y(n_855) );
AOI21xp33_ASAP7_75t_L g856 ( .A1(n_690), .A2(n_17), .B(n_18), .Y(n_856) );
AO31x2_ASAP7_75t_L g857 ( .A1(n_803), .A2(n_527), .A3(n_20), .B(n_18), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_756), .Y(n_858) );
BUFx8_ASAP7_75t_L g859 ( .A(n_717), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_681), .A2(n_527), .B1(n_22), .B2(n_19), .Y(n_860) );
AOI221x1_ASAP7_75t_L g861 ( .A1(n_752), .A2(n_19), .B1(n_21), .B2(n_23), .C(n_24), .Y(n_861) );
INVx8_ASAP7_75t_L g862 ( .A(n_707), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g863 ( .A1(n_802), .A2(n_25), .B(n_21), .C(n_24), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_693), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_864) );
NAND2x1_ASAP7_75t_L g865 ( .A(n_798), .B(n_96), .Y(n_865) );
OAI21xp5_ASAP7_75t_L g866 ( .A1(n_688), .A2(n_102), .B(n_101), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_701), .B(n_26), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_815), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_807), .A2(n_27), .B(n_29), .C(n_30), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_703), .B(n_29), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_708), .Y(n_871) );
INVx3_ASAP7_75t_SL g872 ( .A(n_707), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_722), .A2(n_31), .B(n_32), .C(n_33), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_675), .A2(n_104), .B(n_103), .Y(n_874) );
A2O1A1Ixp33_ASAP7_75t_L g875 ( .A1(n_733), .A2(n_32), .B(n_34), .C(n_35), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_693), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_682), .A2(n_36), .B1(n_38), .B2(n_40), .Y(n_877) );
AOI22x1_ASAP7_75t_SL g878 ( .A1(n_716), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_703), .B(n_42), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_L g880 ( .A1(n_727), .A2(n_43), .B(n_44), .C(n_45), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_696), .A2(n_114), .B(n_110), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_700), .B(n_43), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_691), .A2(n_44), .B1(n_46), .B2(n_47), .Y(n_883) );
INVx3_ASAP7_75t_SL g884 ( .A(n_708), .Y(n_884) );
O2A1O1Ixp33_ASAP7_75t_L g885 ( .A1(n_774), .A2(n_48), .B(n_50), .C(n_51), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_699), .Y(n_886) );
O2A1O1Ixp33_ASAP7_75t_L g887 ( .A1(n_751), .A2(n_51), .B(n_54), .C(n_56), .Y(n_887) );
A2O1A1Ixp33_ASAP7_75t_L g888 ( .A1(n_741), .A2(n_57), .B(n_58), .C(n_59), .Y(n_888) );
A2O1A1Ixp33_ASAP7_75t_L g889 ( .A1(n_749), .A2(n_57), .B(n_58), .C(n_59), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_676), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_890) );
O2A1O1Ixp33_ASAP7_75t_L g891 ( .A1(n_728), .A2(n_60), .B(n_61), .C(n_63), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_780), .A2(n_64), .B1(n_66), .B2(n_67), .Y(n_892) );
O2A1O1Ixp33_ASAP7_75t_L g893 ( .A1(n_704), .A2(n_67), .B(n_68), .C(n_69), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_695), .A2(n_118), .B(n_117), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_770), .Y(n_895) );
OAI21x1_ASAP7_75t_L g896 ( .A1(n_697), .A2(n_120), .B(n_119), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_732), .A2(n_69), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_680), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_814), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_899) );
A2O1A1Ixp33_ASAP7_75t_L g900 ( .A1(n_754), .A2(n_73), .B(n_75), .C(n_76), .Y(n_900) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_713), .A2(n_73), .B1(n_75), .B2(n_76), .C1(n_79), .C2(n_80), .Y(n_901) );
AO32x2_ASAP7_75t_L g902 ( .A1(n_791), .A2(n_782), .A3(n_798), .B1(n_745), .B2(n_773), .Y(n_902) );
NOR3xp33_ASAP7_75t_L g903 ( .A(n_742), .B(n_79), .C(n_80), .Y(n_903) );
A2O1A1Ixp33_ASAP7_75t_L g904 ( .A1(n_759), .A2(n_81), .B(n_82), .C(n_83), .Y(n_904) );
O2A1O1Ixp33_ASAP7_75t_L g905 ( .A1(n_715), .A2(n_81), .B(n_84), .C(n_85), .Y(n_905) );
O2A1O1Ixp33_ASAP7_75t_L g906 ( .A1(n_792), .A2(n_85), .B(n_86), .C(n_87), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_724), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_907) );
AOI222xp33_ASAP7_75t_SL g908 ( .A1(n_763), .A2(n_89), .B1(n_123), .B2(n_124), .C1(n_125), .C2(n_126), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_730), .B(n_128), .Y(n_909) );
O2A1O1Ixp33_ASAP7_75t_L g910 ( .A1(n_740), .A2(n_130), .B(n_133), .C(n_135), .Y(n_910) );
AO31x2_ASAP7_75t_L g911 ( .A1(n_809), .A2(n_139), .A3(n_141), .B(n_142), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_712), .B(n_143), .Y(n_912) );
BUFx10_ASAP7_75t_L g913 ( .A(n_771), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_718), .B(n_145), .Y(n_914) );
OAI21xp5_ASAP7_75t_L g915 ( .A1(n_789), .A2(n_148), .B(n_149), .Y(n_915) );
AOI21x1_ASAP7_75t_L g916 ( .A1(n_797), .A2(n_151), .B(n_152), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_729), .A2(n_153), .B1(n_156), .B2(n_159), .Y(n_917) );
AO21x1_ASAP7_75t_L g918 ( .A1(n_811), .A2(n_160), .B(n_161), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_706), .B(n_162), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_683), .Y(n_920) );
OR2x6_ASAP7_75t_L g921 ( .A(n_709), .B(n_164), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_720), .B(n_166), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_738), .B(n_168), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_822), .A2(n_170), .B(n_171), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_744), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_805), .Y(n_926) );
INVx5_ASAP7_75t_L g927 ( .A(n_758), .Y(n_927) );
AOI21xp5_ASAP7_75t_R g928 ( .A1(n_771), .A2(n_175), .B(n_178), .Y(n_928) );
BUFx6f_ASAP7_75t_L g929 ( .A(n_784), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_813), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_759), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_816), .Y(n_932) );
OAI21xp33_ASAP7_75t_SL g933 ( .A1(n_772), .A2(n_182), .B(n_185), .Y(n_933) );
A2O1A1Ixp33_ASAP7_75t_L g934 ( .A1(n_786), .A2(n_190), .B(n_191), .C(n_192), .Y(n_934) );
A2O1A1Ixp33_ASAP7_75t_L g935 ( .A1(n_778), .A2(n_194), .B(n_195), .C(n_197), .Y(n_935) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_748), .B(n_198), .Y(n_936) );
AO22x1_ASAP7_75t_L g937 ( .A1(n_692), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_818), .B(n_203), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_821), .B(n_205), .Y(n_939) );
AO31x2_ASAP7_75t_L g940 ( .A1(n_795), .A2(n_209), .A3(n_210), .B(n_212), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_750), .B(n_213), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_757), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_760), .A2(n_214), .B(n_216), .C(n_217), .Y(n_943) );
O2A1O1Ixp33_ASAP7_75t_L g944 ( .A1(n_755), .A2(n_219), .B(n_220), .C(n_221), .Y(n_944) );
O2A1O1Ixp33_ASAP7_75t_L g945 ( .A1(n_739), .A2(n_222), .B(n_223), .C(n_224), .Y(n_945) );
AO32x2_ASAP7_75t_L g946 ( .A1(n_772), .A2(n_225), .A3(n_226), .B1(n_227), .B2(n_228), .Y(n_946) );
A2O1A1Ixp33_ASAP7_75t_L g947 ( .A1(n_743), .A2(n_229), .B(n_230), .C(n_232), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_750), .A2(n_238), .B1(n_239), .B2(n_243), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_765), .B(n_244), .C(n_246), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_692), .B(n_248), .Y(n_950) );
OAI22x1_ASAP7_75t_L g951 ( .A1(n_793), .A2(n_249), .B1(n_251), .B2(n_253), .Y(n_951) );
OAI21x1_ASAP7_75t_L g952 ( .A1(n_769), .A2(n_255), .B(n_257), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_746), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g954 ( .A(n_753), .B(n_258), .C(n_261), .Y(n_954) );
AO31x2_ASAP7_75t_L g955 ( .A1(n_787), .A2(n_266), .A3(n_267), .B(n_268), .Y(n_955) );
AOI221xp5_ASAP7_75t_SL g956 ( .A1(n_766), .A2(n_270), .B1(n_271), .B2(n_272), .C(n_279), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_758), .B(n_321), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_719), .B(n_282), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_767), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_775), .B(n_284), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_804), .A2(n_288), .B1(n_290), .B2(n_293), .Y(n_961) );
AO32x2_ASAP7_75t_L g962 ( .A1(n_793), .A2(n_294), .A3(n_298), .B1(n_304), .B2(n_306), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_689), .B(n_317), .Y(n_963) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_784), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_777), .B(n_307), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_767), .B(n_316), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_785), .A2(n_796), .B(n_779), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_677), .B(n_781), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_783), .Y(n_969) );
AO32x2_ASAP7_75t_L g970 ( .A1(n_768), .A2(n_747), .A3(n_803), .B1(n_752), .B2(n_791), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_768), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_768), .B(n_788), .Y(n_972) );
BUFx3_ASAP7_75t_L g973 ( .A(n_768), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_768), .Y(n_974) );
O2A1O1Ixp33_ASAP7_75t_L g975 ( .A1(n_794), .A2(n_737), .B(n_666), .C(n_723), .Y(n_975) );
NAND2xp33_ASAP7_75t_L g976 ( .A(n_675), .B(n_653), .Y(n_976) );
AOI21xp5_ASAP7_75t_L g977 ( .A1(n_705), .A2(n_599), .B(n_597), .Y(n_977) );
OAI21x1_ASAP7_75t_L g978 ( .A1(n_799), .A2(n_762), .B(n_697), .Y(n_978) );
O2A1O1Ixp33_ASAP7_75t_SL g979 ( .A1(n_776), .A2(n_737), .B(n_810), .C(n_817), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_942), .Y(n_980) );
AND2x6_ASAP7_75t_SL g981 ( .A(n_921), .B(n_846), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_886), .B(n_871), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_926), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_930), .B(n_932), .Y(n_984) );
AND2x4_ASAP7_75t_SL g985 ( .A(n_921), .B(n_913), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g986 ( .A1(n_829), .A2(n_979), .B(n_854), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_845), .B(n_851), .Y(n_987) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_841), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_884), .B(n_825), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_977), .A2(n_837), .B(n_824), .Y(n_990) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_876), .A2(n_864), .B1(n_834), .B2(n_823), .Y(n_991) );
OAI22x1_ASAP7_75t_L g992 ( .A1(n_825), .A2(n_836), .B1(n_890), .B2(n_855), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_851), .Y(n_993) );
INVx2_ASAP7_75t_SL g994 ( .A(n_849), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_868), .B(n_828), .Y(n_995) );
NOR2x1_ASAP7_75t_R g996 ( .A(n_927), .B(n_836), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g997 ( .A(n_872), .B(n_862), .Y(n_997) );
INVx2_ASAP7_75t_SL g998 ( .A(n_826), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_898), .B(n_925), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_859), .A2(n_867), .B1(n_903), .B2(n_862), .Y(n_1000) );
AOI21xp5_ASAP7_75t_L g1001 ( .A1(n_842), .A2(n_967), .B(n_939), .Y(n_1001) );
INVx5_ASAP7_75t_L g1002 ( .A(n_927), .Y(n_1002) );
OA21x2_ASAP7_75t_L g1003 ( .A1(n_956), .A2(n_896), .B(n_952), .Y(n_1003) );
OA21x2_ASAP7_75t_L g1004 ( .A1(n_915), .A2(n_866), .B(n_861), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_826), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_844), .Y(n_1006) );
INVxp67_ASAP7_75t_L g1007 ( .A(n_859), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_870), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_850), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_839), .B(n_913), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_882), .A2(n_856), .B1(n_860), .B2(n_901), .Y(n_1011) );
AO31x2_ASAP7_75t_L g1012 ( .A1(n_918), .A2(n_951), .A3(n_869), .B(n_863), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_827), .B(n_848), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_879), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_953), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_858), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_895), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_847), .A2(n_843), .B(n_975), .Y(n_1018) );
OAI222xp33_ASAP7_75t_L g1019 ( .A1(n_878), .A2(n_892), .B1(n_883), .B2(n_907), .C1(n_877), .C2(n_830), .Y(n_1019) );
AOI21xp5_ASAP7_75t_L g1020 ( .A1(n_976), .A2(n_923), .B(n_909), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_920), .B(n_832), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_927), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_914), .A2(n_912), .B1(n_897), .B2(n_831), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_957), .B(n_973), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_857), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_857), .Y(n_1026) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_938), .A2(n_853), .B(n_833), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_928), .A2(n_957), .B1(n_835), .B2(n_873), .Y(n_1028) );
AO21x2_ASAP7_75t_L g1029 ( .A1(n_916), .A2(n_941), .B(n_954), .Y(n_1029) );
INVx4_ASAP7_75t_SL g1030 ( .A(n_955), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_880), .Y(n_1031) );
INVx4_ASAP7_75t_L g1032 ( .A(n_929), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_887), .B(n_885), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_959), .Y(n_1034) );
OR2x6_ASAP7_75t_L g1035 ( .A(n_937), .B(n_906), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_919), .B(n_922), .Y(n_1036) );
OA21x2_ASAP7_75t_L g1037 ( .A1(n_924), .A2(n_894), .B(n_881), .Y(n_1037) );
OA21x2_ASAP7_75t_L g1038 ( .A1(n_874), .A2(n_935), .B(n_943), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_893), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_969), .B(n_899), .Y(n_1040) );
AOI21xp5_ASAP7_75t_L g1041 ( .A1(n_960), .A2(n_965), .B(n_972), .Y(n_1041) );
A2O1A1Ixp33_ASAP7_75t_L g1042 ( .A1(n_905), .A2(n_891), .B(n_933), .C(n_936), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_904), .B(n_875), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_900), .B(n_852), .Y(n_1044) );
OAI21x1_ASAP7_75t_L g1045 ( .A1(n_865), .A2(n_974), .B(n_971), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_968), .A2(n_958), .B1(n_838), .B2(n_931), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_911), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_889), .Y(n_1048) );
OA21x2_ASAP7_75t_L g1049 ( .A1(n_947), .A2(n_934), .B(n_949), .Y(n_1049) );
BUFx4f_ASAP7_75t_L g1050 ( .A(n_929), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_888), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_970), .B(n_946), .Y(n_1052) );
AO31x2_ASAP7_75t_L g1053 ( .A1(n_948), .A2(n_966), .A3(n_963), .B(n_950), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_964), .B(n_961), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_964), .B(n_917), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_940), .B(n_911), .Y(n_1056) );
BUFx8_ASAP7_75t_SL g1057 ( .A(n_908), .Y(n_1057) );
NAND3xp33_ASAP7_75t_L g1058 ( .A(n_945), .B(n_910), .C(n_944), .Y(n_1058) );
INVx4_ASAP7_75t_SL g1059 ( .A(n_955), .Y(n_1059) );
OA21x2_ASAP7_75t_L g1060 ( .A1(n_962), .A2(n_978), .B(n_956), .Y(n_1060) );
INVx4_ASAP7_75t_SL g1061 ( .A(n_962), .Y(n_1061) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_902), .A2(n_628), .B1(n_721), .B2(n_834), .C(n_589), .Y(n_1062) );
OAI21xp5_ASAP7_75t_L g1063 ( .A1(n_902), .A2(n_711), .B(n_977), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1064 ( .A1(n_902), .A2(n_829), .B(n_979), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_825), .A2(n_747), .B1(n_736), .B2(n_630), .Y(n_1065) );
BUFx8_ASAP7_75t_L g1066 ( .A(n_825), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_884), .B(n_631), .Y(n_1067) );
BUFx10_ASAP7_75t_L g1068 ( .A(n_825), .Y(n_1068) );
A2O1A1Ixp33_ASAP7_75t_L g1069 ( .A1(n_855), .A2(n_812), .B(n_802), .C(n_807), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_834), .A2(n_747), .B1(n_721), .B2(n_640), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_884), .B(n_625), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_841), .Y(n_1072) );
A2O1A1Ixp33_ASAP7_75t_L g1073 ( .A1(n_855), .A2(n_812), .B(n_802), .C(n_807), .Y(n_1073) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_829), .A2(n_979), .B(n_810), .Y(n_1074) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_886), .B(n_927), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_942), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1077 ( .A1(n_829), .A2(n_979), .B(n_810), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_886), .B(n_613), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_884), .B(n_631), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_942), .Y(n_1080) );
NAND2xp5_ASAP7_75t_SL g1081 ( .A(n_823), .B(n_808), .Y(n_1081) );
INVxp67_ASAP7_75t_L g1082 ( .A(n_825), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_898), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_834), .A2(n_747), .B1(n_721), .B2(n_640), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_942), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_886), .B(n_613), .Y(n_1086) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_834), .A2(n_690), .B1(n_687), .B2(n_611), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_834), .A2(n_690), .B1(n_687), .B2(n_611), .Y(n_1088) );
AO31x2_ASAP7_75t_L g1089 ( .A1(n_918), .A2(n_854), .A3(n_840), .B(n_817), .Y(n_1089) );
AO21x2_ASAP7_75t_L g1090 ( .A1(n_978), .A2(n_854), .B(n_800), .Y(n_1090) );
INVxp67_ASAP7_75t_L g1091 ( .A(n_825), .Y(n_1091) );
OR2x2_ASAP7_75t_L g1092 ( .A(n_884), .B(n_625), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_884), .B(n_631), .Y(n_1093) );
AOI21xp5_ASAP7_75t_L g1094 ( .A1(n_829), .A2(n_979), .B(n_810), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_942), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_884), .B(n_625), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_849), .Y(n_1097) );
OR2x6_ASAP7_75t_L g1098 ( .A(n_921), .B(n_801), .Y(n_1098) );
INVx3_ASAP7_75t_SL g1099 ( .A(n_846), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_942), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_849), .Y(n_1101) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_834), .A2(n_690), .B1(n_687), .B2(n_611), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_884), .B(n_631), .Y(n_1103) );
OAI211xp5_ASAP7_75t_L g1104 ( .A1(n_901), .A2(n_693), .B(n_589), .C(n_876), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_942), .Y(n_1105) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_841), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_898), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_876), .A2(n_693), .B1(n_806), .B2(n_678), .Y(n_1108) );
OR2x6_ASAP7_75t_L g1109 ( .A(n_921), .B(n_801), .Y(n_1109) );
OAI222xp33_ASAP7_75t_L g1110 ( .A1(n_878), .A2(n_693), .B1(n_921), .B2(n_876), .C1(n_722), .C2(n_864), .Y(n_1110) );
A2O1A1Ixp33_ASAP7_75t_L g1111 ( .A1(n_855), .A2(n_812), .B(n_802), .C(n_807), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_942), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_996), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_999), .B(n_1083), .Y(n_1114) );
AOI21xp5_ASAP7_75t_SL g1115 ( .A1(n_1028), .A2(n_1024), .B(n_992), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1107), .B(n_983), .Y(n_1116) );
NOR2x1_ASAP7_75t_L g1117 ( .A(n_1098), .B(n_1109), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_983), .B(n_1076), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1080), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1080), .B(n_1085), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1121 ( .A(n_1002), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1085), .B(n_1095), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_1100), .B(n_1105), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1100), .B(n_1105), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1112), .B(n_1016), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1112), .B(n_1017), .Y(n_1126) );
AND2x4_ASAP7_75t_L g1127 ( .A(n_1032), .B(n_1075), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1025), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1026), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_984), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1015), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_987), .B(n_993), .Y(n_1132) );
OR2x6_ASAP7_75t_L g1133 ( .A(n_1098), .B(n_1109), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1134 ( .A(n_1002), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_982), .Y(n_1135) );
BUFx3_ASAP7_75t_L g1136 ( .A(n_1002), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1060), .Y(n_1137) );
AO21x2_ASAP7_75t_L g1138 ( .A1(n_1063), .A2(n_1001), .B(n_990), .Y(n_1138) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_1075), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1061), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1065), .B(n_1051), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_1066), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1061), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1052), .Y(n_1144) );
OAI21xp5_ASAP7_75t_L g1145 ( .A1(n_1069), .A2(n_1111), .B(n_1073), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_1050), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_995), .Y(n_1147) );
BUFx6f_ASAP7_75t_L g1148 ( .A(n_1050), .Y(n_1148) );
BUFx3_ASAP7_75t_L g1149 ( .A(n_1022), .Y(n_1149) );
AO21x2_ASAP7_75t_L g1150 ( .A1(n_1074), .A2(n_1077), .B(n_1094), .Y(n_1150) );
INVx3_ASAP7_75t_L g1151 ( .A(n_1032), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_1070), .A2(n_1084), .B1(n_1011), .B2(n_1082), .Y(n_1152) );
BUFx3_ASAP7_75t_L g1153 ( .A(n_1066), .Y(n_1153) );
AOI322xp5_ASAP7_75t_L g1154 ( .A1(n_1108), .A2(n_1087), .A3(n_1088), .B1(n_1102), .B2(n_1000), .C1(n_1007), .C2(n_1091), .Y(n_1154) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_989), .Y(n_1155) );
OAI222xp33_ASAP7_75t_L g1156 ( .A1(n_1035), .A2(n_1062), .B1(n_991), .B2(n_1044), .C1(n_1033), .C2(n_1057), .Y(n_1156) );
INVx2_ASAP7_75t_SL g1157 ( .A(n_985), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_1036), .A2(n_1023), .B1(n_1035), .B2(n_1031), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1006), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1034), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g1161 ( .A(n_1042), .B(n_1039), .C(n_1048), .Y(n_1161) );
OR2x6_ASAP7_75t_L g1162 ( .A(n_1081), .B(n_1027), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1008), .B(n_1014), .Y(n_1163) );
AOI21x1_ASAP7_75t_L g1164 ( .A1(n_986), .A2(n_1003), .B(n_1018), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1078), .Y(n_1165) );
BUFx3_ASAP7_75t_L g1166 ( .A(n_1099), .Y(n_1166) );
INVx3_ASAP7_75t_L g1167 ( .A(n_1068), .Y(n_1167) );
AOI33xp33_ASAP7_75t_L g1168 ( .A1(n_1067), .A2(n_1079), .A3(n_1103), .B1(n_1093), .B2(n_994), .B3(n_1097), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1086), .B(n_1068), .Y(n_1169) );
INVxp67_ASAP7_75t_L g1170 ( .A(n_1071), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1171 ( .A(n_1013), .Y(n_1171) );
AO21x2_ASAP7_75t_L g1172 ( .A1(n_1041), .A2(n_1090), .B(n_1029), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1043), .B(n_1012), .Y(n_1173) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1045), .B(n_1059), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1104), .B(n_1106), .Y(n_1175) );
BUFx3_ASAP7_75t_L g1176 ( .A(n_998), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_988), .B(n_1092), .Y(n_1177) );
AO21x2_ASAP7_75t_L g1178 ( .A1(n_1058), .A2(n_1020), .B(n_1055), .Y(n_1178) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1030), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1012), .B(n_1040), .Y(n_1180) );
OAI31xp33_ASAP7_75t_L g1181 ( .A1(n_1110), .A2(n_1019), .A3(n_1010), .B(n_1096), .Y(n_1181) );
OAI21xp5_ASAP7_75t_L g1182 ( .A1(n_1046), .A2(n_1054), .B(n_1004), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_1005), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1072), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_997), .B(n_1021), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1012), .B(n_1101), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1053), .B(n_1038), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1188 ( .A(n_981), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1009), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1089), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1053), .B(n_1038), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1049), .B(n_1037), .Y(n_1192) );
BUFx3_ASAP7_75t_L g1193 ( .A(n_1002), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_980), .Y(n_1194) );
AO21x2_ASAP7_75t_L g1195 ( .A1(n_1056), .A2(n_1064), .B(n_1063), .Y(n_1195) );
OA21x2_ASAP7_75t_L g1196 ( .A1(n_1056), .A2(n_1064), .B(n_1047), .Y(n_1196) );
OR2x6_ASAP7_75t_L g1197 ( .A(n_1098), .B(n_1109), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_980), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1078), .B(n_693), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1144), .B(n_1186), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1128), .Y(n_1201) );
NOR2xp33_ASAP7_75t_SL g1202 ( .A(n_1117), .B(n_1156), .Y(n_1202) );
AO21x2_ASAP7_75t_L g1203 ( .A1(n_1164), .A2(n_1182), .B(n_1145), .Y(n_1203) );
INVx1_ASAP7_75t_SL g1204 ( .A(n_1139), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1144), .B(n_1173), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1128), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1186), .B(n_1180), .Y(n_1207) );
INVx5_ASAP7_75t_SL g1208 ( .A(n_1133), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1129), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1173), .B(n_1180), .Y(n_1210) );
AND2x4_ASAP7_75t_L g1211 ( .A(n_1179), .B(n_1140), .Y(n_1211) );
INVx3_ASAP7_75t_L g1212 ( .A(n_1174), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1120), .B(n_1122), .Y(n_1213) );
BUFx3_ASAP7_75t_L g1214 ( .A(n_1127), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1120), .B(n_1122), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1194), .B(n_1198), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1137), .Y(n_1217) );
AOI221xp5_ASAP7_75t_SL g1218 ( .A1(n_1152), .A2(n_1158), .B1(n_1175), .B2(n_1141), .C(n_1170), .Y(n_1218) );
AOI21xp33_ASAP7_75t_L g1219 ( .A1(n_1161), .A2(n_1181), .B(n_1178), .Y(n_1219) );
AND2x4_ASAP7_75t_L g1220 ( .A(n_1179), .B(n_1140), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_1141), .A2(n_1199), .B1(n_1165), .B2(n_1197), .Y(n_1221) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_1174), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1125), .B(n_1126), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1187), .B(n_1191), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1187), .B(n_1191), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1118), .B(n_1123), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_1133), .A2(n_1197), .B1(n_1169), .B2(n_1188), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1190), .B(n_1143), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1126), .B(n_1119), .Y(n_1229) );
BUFx2_ASAP7_75t_L g1230 ( .A(n_1162), .Y(n_1230) );
BUFx3_ASAP7_75t_L g1231 ( .A(n_1136), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1118), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1123), .B(n_1124), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1124), .Y(n_1234) );
BUFx2_ASAP7_75t_L g1235 ( .A(n_1162), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1163), .B(n_1130), .Y(n_1236) );
INVx2_ASAP7_75t_SL g1237 ( .A(n_1136), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1163), .B(n_1131), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1116), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1116), .B(n_1160), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1171), .B(n_1114), .Y(n_1241) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_1162), .Y(n_1242) );
NOR2xp33_ASAP7_75t_L g1243 ( .A(n_1236), .B(n_1185), .Y(n_1243) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1217), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1210), .B(n_1192), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1205), .B(n_1168), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1207), .B(n_1195), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1205), .B(n_1135), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1236), .B(n_1189), .Y(n_1249) );
BUFx3_ASAP7_75t_L g1250 ( .A(n_1231), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1207), .B(n_1195), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1224), .B(n_1196), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1225), .B(n_1138), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1225), .B(n_1138), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1200), .B(n_1184), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_1222), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1232), .B(n_1147), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1213), .B(n_1178), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_1241), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1232), .B(n_1159), .Y(n_1260) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_1204), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1213), .B(n_1178), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1234), .B(n_1154), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1234), .B(n_1239), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1200), .B(n_1177), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1239), .B(n_1115), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1228), .B(n_1150), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1201), .Y(n_1268) );
BUFx3_ASAP7_75t_L g1269 ( .A(n_1231), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1215), .B(n_1172), .Y(n_1270) );
AOI22xp33_ASAP7_75t_SL g1271 ( .A1(n_1202), .A2(n_1197), .B1(n_1133), .B2(n_1113), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1215), .B(n_1172), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1201), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1206), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1240), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1209), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1226), .B(n_1197), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1245), .B(n_1203), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1245), .B(n_1203), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1268), .Y(n_1280) );
AOI21x1_ASAP7_75t_SL g1281 ( .A1(n_1263), .A2(n_1220), .B(n_1211), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1245), .B(n_1203), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1268), .Y(n_1283) );
OR2x6_ASAP7_75t_L g1284 ( .A(n_1256), .B(n_1222), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1253), .B(n_1203), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1275), .B(n_1223), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1253), .B(n_1223), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1254), .B(n_1212), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1289 ( .A(n_1250), .Y(n_1289) );
AND2x4_ASAP7_75t_L g1290 ( .A(n_1267), .B(n_1212), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1273), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1244), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1247), .B(n_1251), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1254), .B(n_1212), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1274), .Y(n_1295) );
OR2x6_ASAP7_75t_L g1296 ( .A(n_1256), .B(n_1115), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_1261), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1298 ( .A(n_1259), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1276), .Y(n_1299) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1251), .B(n_1233), .Y(n_1300) );
INVx1_ASAP7_75t_SL g1301 ( .A(n_1250), .Y(n_1301) );
NOR3xp33_ASAP7_75t_L g1302 ( .A(n_1271), .B(n_1219), .C(n_1218), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1258), .B(n_1216), .Y(n_1303) );
BUFx2_ASAP7_75t_L g1304 ( .A(n_1269), .Y(n_1304) );
NOR2xp33_ASAP7_75t_L g1305 ( .A(n_1243), .B(n_1188), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1258), .B(n_1216), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1298), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1287), .B(n_1262), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1287), .B(n_1262), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1278), .B(n_1252), .Y(n_1310) );
NAND3xp33_ASAP7_75t_L g1311 ( .A(n_1302), .B(n_1218), .C(n_1271), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1297), .B(n_1270), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1300), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g1314 ( .A1(n_1284), .A2(n_1227), .B1(n_1133), .B2(n_1221), .Y(n_1314) );
A2O1A1Ixp33_ASAP7_75t_L g1315 ( .A1(n_1305), .A2(n_1202), .B(n_1227), .C(n_1221), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1280), .Y(n_1316) );
OAI22xp33_ASAP7_75t_L g1317 ( .A1(n_1296), .A2(n_1246), .B1(n_1277), .B2(n_1266), .Y(n_1317) );
NOR2xp67_ASAP7_75t_SL g1318 ( .A(n_1304), .B(n_1153), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1280), .Y(n_1319) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1304), .A2(n_1142), .B(n_1183), .Y(n_1320) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1286), .B(n_1249), .Y(n_1321) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1292), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1293), .B(n_1252), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1283), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1278), .B(n_1252), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1283), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1291), .Y(n_1327) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_1296), .A2(n_1277), .B1(n_1257), .B2(n_1255), .C(n_1266), .Y(n_1328) );
OR2x6_ASAP7_75t_L g1329 ( .A(n_1320), .B(n_1153), .Y(n_1329) );
O2A1O1Ixp33_ASAP7_75t_L g1330 ( .A1(n_1311), .A2(n_1166), .B(n_1183), .C(n_1155), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_1314), .A2(n_1290), .B1(n_1282), .B2(n_1279), .Y(n_1331) );
AOI22xp5_ASAP7_75t_L g1332 ( .A1(n_1318), .A2(n_1270), .B1(n_1272), .B2(n_1248), .Y(n_1332) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1322), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1323), .B(n_1303), .Y(n_1334) );
NAND2xp5_ASAP7_75t_SL g1335 ( .A(n_1315), .B(n_1289), .Y(n_1335) );
NAND2x1p5_ASAP7_75t_L g1336 ( .A(n_1307), .B(n_1193), .Y(n_1336) );
NOR2x1_ASAP7_75t_L g1337 ( .A(n_1317), .B(n_1269), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1313), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1316), .Y(n_1339) );
AOI221xp5_ASAP7_75t_L g1340 ( .A1(n_1317), .A2(n_1306), .B1(n_1285), .B2(n_1294), .C(n_1288), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1319), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1339), .Y(n_1342) );
AOI22xp5_ASAP7_75t_L g1343 ( .A1(n_1335), .A2(n_1328), .B1(n_1321), .B2(n_1312), .Y(n_1343) );
AOI221xp5_ASAP7_75t_L g1344 ( .A1(n_1340), .A2(n_1321), .B1(n_1310), .B2(n_1325), .C(n_1308), .Y(n_1344) );
OAI21xp5_ASAP7_75t_SL g1345 ( .A1(n_1337), .A2(n_1301), .B(n_1157), .Y(n_1345) );
OAI21xp33_ASAP7_75t_L g1346 ( .A1(n_1331), .A2(n_1325), .B(n_1309), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1341), .Y(n_1347) );
A2O1A1Ixp33_ASAP7_75t_L g1348 ( .A1(n_1330), .A2(n_1289), .B(n_1269), .C(n_1157), .Y(n_1348) );
AOI21xp33_ASAP7_75t_L g1349 ( .A1(n_1329), .A2(n_1134), .B(n_1121), .Y(n_1349) );
NAND3xp33_ASAP7_75t_SL g1350 ( .A(n_1345), .B(n_1336), .C(n_1332), .Y(n_1350) );
A2O1A1Ixp33_ASAP7_75t_L g1351 ( .A1(n_1346), .A2(n_1338), .B(n_1334), .C(n_1121), .Y(n_1351) );
AOI221xp5_ASAP7_75t_L g1352 ( .A1(n_1344), .A2(n_1327), .B1(n_1326), .B2(n_1324), .C(n_1333), .Y(n_1352) );
OAI211xp5_ASAP7_75t_SL g1353 ( .A1(n_1343), .A2(n_1265), .B(n_1257), .C(n_1238), .Y(n_1353) );
AOI221x1_ASAP7_75t_L g1354 ( .A1(n_1348), .A2(n_1151), .B1(n_1291), .B2(n_1299), .C(n_1295), .Y(n_1354) );
O2A1O1Ixp33_ASAP7_75t_L g1355 ( .A1(n_1349), .A2(n_1176), .B(n_1167), .C(n_1237), .Y(n_1355) );
OAI211xp5_ASAP7_75t_SL g1356 ( .A1(n_1351), .A2(n_1347), .B(n_1342), .C(n_1167), .Y(n_1356) );
OAI211xp5_ASAP7_75t_SL g1357 ( .A1(n_1352), .A2(n_1167), .B(n_1265), .C(n_1238), .Y(n_1357) );
AOI22xp5_ASAP7_75t_L g1358 ( .A1(n_1350), .A2(n_1290), .B1(n_1270), .B2(n_1272), .Y(n_1358) );
NAND4xp25_ASAP7_75t_L g1359 ( .A(n_1358), .B(n_1354), .C(n_1355), .D(n_1353), .Y(n_1359) );
OR5x1_ASAP7_75t_L g1360 ( .A(n_1359), .B(n_1356), .C(n_1357), .D(n_1208), .E(n_1281), .Y(n_1360) );
OAI22xp5_ASAP7_75t_SL g1361 ( .A1(n_1360), .A2(n_1149), .B1(n_1146), .B2(n_1237), .Y(n_1361) );
NOR2x2_ASAP7_75t_L g1362 ( .A(n_1361), .B(n_1162), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_1362), .A2(n_1208), .B1(n_1260), .B2(n_1264), .Y(n_1363) );
AOI21xp5_ASAP7_75t_L g1364 ( .A1(n_1363), .A2(n_1148), .B(n_1132), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_1364), .A2(n_1208), .B1(n_1148), .B2(n_1214), .Y(n_1365) );
AOI221xp5_ASAP7_75t_SL g1366 ( .A1(n_1365), .A2(n_1242), .B1(n_1235), .B2(n_1230), .C(n_1229), .Y(n_1366) );
endmodule