module fake_jpeg_31857_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_57),
.B(n_59),
.C(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_61),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_17),
.B1(n_38),
.B2(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_51),
.B1(n_48),
.B2(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_7),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_51),
.B1(n_47),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_62),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_45),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_8),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_85),
.B(n_22),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_6),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_84),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_41),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_23),
.B(n_34),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_24),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_98),
.C(n_86),
.Y(n_103)
);

AOI221xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_96),
.B1(n_90),
.B2(n_31),
.C(n_33),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_21),
.C(n_25),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_109),
.Y(n_111)
);

XNOR2x1_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_109),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_103),
.C(n_102),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_113),
.B1(n_112),
.B2(n_111),
.Y(n_118)
);

OAI321xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_106),
.A3(n_104),
.B1(n_39),
.B2(n_28),
.C(n_26),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_100),
.Y(n_120)
);


endmodule