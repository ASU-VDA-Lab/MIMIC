module fake_jpeg_18016_n_355 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_355);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_30),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_54),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_55),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_1),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_28),
.B1(n_36),
.B2(n_22),
.Y(n_98)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx9p33_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_87),
.Y(n_101)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_84),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_50),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_31),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_38),
.C(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_51),
.B(n_35),
.Y(n_87)
);

CKINVDCx6p67_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_104),
.Y(n_131)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_109),
.B1(n_32),
.B2(n_23),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_25),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_105),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_31),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_32),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_25),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_31),
.B1(n_23),
.B2(n_29),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_116),
.Y(n_125)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_63),
.B1(n_77),
.B2(n_68),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_126),
.B1(n_139),
.B2(n_96),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_58),
.B(n_67),
.C(n_35),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_113),
.B(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_59),
.B1(n_73),
.B2(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_137),
.Y(n_165)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_25),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_37),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_102),
.Y(n_146)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_29),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_157),
.B1(n_158),
.B2(n_146),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_101),
.B1(n_97),
.B2(n_94),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_97),
.B1(n_65),
.B2(n_80),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_119),
.A2(n_65),
.B1(n_78),
.B2(n_76),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_173),
.B1(n_169),
.B2(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_78),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_170),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_128),
.B1(n_125),
.B2(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_127),
.B1(n_147),
.B2(n_120),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_116),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_29),
.B(n_32),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_44),
.C(n_112),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_152),
.C(n_173),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_72),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_89),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_190),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_175),
.B(n_181),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_178),
.C(n_192),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_123),
.C(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_179),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_182),
.B(n_176),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_130),
.B1(n_121),
.B2(n_120),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_121),
.B1(n_148),
.B2(n_149),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_110),
.B1(n_67),
.B2(n_89),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_157),
.B1(n_173),
.B2(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_134),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_130),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_191),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_164),
.C(n_158),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_154),
.Y(n_220)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_209),
.B1(n_129),
.B2(n_141),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_173),
.B1(n_163),
.B2(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_200),
.A2(n_205),
.B1(n_213),
.B2(n_162),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_170),
.B1(n_161),
.B2(n_169),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_209),
.A2(n_195),
.B(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

AO22x2_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_161),
.B1(n_169),
.B2(n_72),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_156),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_218),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_193),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_129),
.B1(n_150),
.B2(n_162),
.Y(n_240)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_162),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_138),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_177),
.C(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_182),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_225),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_228),
.C(n_233),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_224),
.A2(n_241),
.B(n_207),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_202),
.B1(n_198),
.B2(n_210),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_178),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_187),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_200),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_199),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_176),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_203),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_219),
.B1(n_197),
.B2(n_208),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_244),
.B1(n_204),
.B2(n_218),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_208),
.B1(n_217),
.B2(n_138),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_92),
.B1(n_27),
.B2(n_33),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_201),
.B(n_118),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_112),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_258),
.Y(n_275)
);

NOR2x1_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_213),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_250),
.B(n_265),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_254),
.B(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_199),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_263),
.B1(n_268),
.B2(n_2),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_227),
.B(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_244),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_207),
.B1(n_212),
.B2(n_211),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_215),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_223),
.CI(n_238),
.CON(n_266),
.SN(n_266)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_236),
.CI(n_224),
.CON(n_271),
.SN(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_79),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_228),
.C(n_238),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_272),
.C(n_278),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_242),
.C(n_229),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_284),
.C(n_288),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_217),
.B1(n_105),
.B2(n_136),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_268),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_285),
.B1(n_35),
.B2(n_27),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_136),
.C(n_79),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_255),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_136),
.C(n_37),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_37),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_30),
.C(n_38),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_249),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_303),
.C(n_304),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_248),
.B(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_253),
.B(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_258),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_271),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_284),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_264),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_6),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_279),
.C(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_315),
.C(n_318),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_288),
.C(n_281),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_304),
.C(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_282),
.C(n_38),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_291),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_320),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_289),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_323),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_307),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_319),
.C(n_324),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_307),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_24),
.B(n_20),
.Y(n_337)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_39),
.B1(n_33),
.B2(n_27),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_309),
.A2(n_282),
.B(n_39),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_24),
.B(n_20),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_335),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_333),
.A2(n_337),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_7),
.B(n_8),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_8),
.B(n_9),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_338),
.A2(n_11),
.B(n_12),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_38),
.C(n_9),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_326),
.B(n_322),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_340),
.A2(n_342),
.B(n_345),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_341),
.Y(n_346)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_325),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_11),
.C2(n_17),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_344),
.A3(n_338),
.B1(n_339),
.B2(n_336),
.C1(n_331),
.C2(n_18),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_349),
.A2(n_350),
.B(n_347),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_15),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_15),
.B(n_16),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_352),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_16),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_354),
.B(n_17),
.Y(n_355)
);


endmodule