module fake_jpeg_15461_n_215 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_57),
.B1(n_62),
.B2(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_52),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_25),
.B(n_28),
.C(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_15),
.B1(n_27),
.B2(n_23),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_42),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_41),
.B1(n_39),
.B2(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_27),
.B1(n_20),
.B2(n_18),
.Y(n_62)
);

AO22x2_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_32),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_65),
.B1(n_63),
.B2(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_39),
.B1(n_33),
.B2(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_72),
.B1(n_63),
.B2(n_65),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_73),
.B1(n_54),
.B2(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_32),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_63),
.C(n_32),
.Y(n_85)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_30),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_73),
.C(n_78),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_98),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_59),
.B1(n_48),
.B2(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_30),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_48),
.B1(n_50),
.B2(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_85),
.C(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_64),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_88),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_120),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_118),
.B(n_57),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_64),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_81),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_128),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_108),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_57),
.B(n_50),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_121),
.B1(n_109),
.B2(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_94),
.B1(n_98),
.B2(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_70),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_94),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_84),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.C(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_113),
.B1(n_116),
.B2(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_151),
.B1(n_158),
.B2(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_134),
.B1(n_131),
.B2(n_142),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_126),
.B1(n_129),
.B2(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_118),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_104),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_159),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_110),
.B1(n_120),
.B2(n_72),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_50),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_163),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_72),
.C(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_169),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_124),
.B1(n_100),
.B2(n_51),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_155),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_153),
.B(n_148),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_168),
.B(n_162),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_156),
.B(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_172),
.B1(n_167),
.B2(n_169),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_51),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_185),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_91),
.B1(n_14),
.B2(n_10),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_172),
.C(n_167),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_192),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_47),
.C(n_32),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_178),
.A3(n_177),
.B1(n_184),
.B2(n_176),
.C1(n_52),
.C2(n_56),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_201),
.C(n_19),
.Y(n_204)
);

OAI321xp33_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_10),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_6),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_1),
.B(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_194),
.B1(n_17),
.B2(n_8),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_204),
.Y(n_208)
);

AOI31xp33_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_206),
.B(n_7),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_9),
.B(n_34),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_34),
.C(n_8),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_202),
.A2(n_197),
.B(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.C(n_9),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_208),
.B1(n_9),
.B2(n_34),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_211),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);


endmodule