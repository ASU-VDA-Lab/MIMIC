module real_jpeg_4608_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_0),
.Y(n_195)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_0),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_0),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_0),
.Y(n_370)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_1),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_1),
.Y(n_412)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_1),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_2),
.A2(n_48),
.B1(n_128),
.B2(n_253),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_2),
.A2(n_48),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_2),
.A2(n_48),
.B1(n_246),
.B2(n_443),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_3),
.A2(n_247),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_3),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_3),
.A2(n_296),
.B1(n_304),
.B2(n_325),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_3),
.A2(n_137),
.B1(n_304),
.B2(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_3),
.A2(n_304),
.B1(n_411),
.B2(n_463),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_92),
.B1(n_93),
.B2(n_98),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_4),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_98),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_98),
.B1(n_197),
.B2(n_203),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_6),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_6),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_6),
.A2(n_92),
.B1(n_213),
.B2(n_277),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_6),
.A2(n_213),
.B1(n_296),
.B2(n_299),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_6),
.A2(n_213),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_7),
.Y(n_511)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_8),
.Y(n_284)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_10),
.A2(n_269),
.B1(n_271),
.B2(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_10),
.B(n_284),
.C(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_10),
.B(n_114),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_10),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_10),
.B(n_90),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_10),
.B(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_12),
.Y(n_514)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_14),
.A2(n_135),
.B1(n_137),
.B2(n_140),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_14),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_140),
.B1(n_166),
.B2(n_170),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_14),
.A2(n_140),
.B1(n_236),
.B2(n_240),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_15),
.A2(n_58),
.B1(n_157),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_15),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_15),
.A2(n_256),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_15),
.A2(n_92),
.B1(n_248),
.B2(n_256),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_15),
.A2(n_253),
.B1(n_256),
.B2(n_440),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_16),
.A2(n_52),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_16),
.A2(n_59),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_16),
.A2(n_59),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_16),
.A2(n_59),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_18),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_18),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_18),
.A2(n_127),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_18),
.A2(n_94),
.B1(n_127),
.B2(n_208),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_18),
.A2(n_127),
.B1(n_198),
.B2(n_427),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_509),
.B(n_512),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_220),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_219),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_159),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_24),
.B(n_159),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_141),
.B2(n_142),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_60),
.C(n_99),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_27),
.A2(n_143),
.B1(n_144),
.B2(n_158),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_27),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_27),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_46),
.B1(n_54),
.B2(n_56),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_28),
.A2(n_54),
.B1(n_56),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_28),
.A2(n_255),
.B(n_257),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_28),
.A2(n_54),
.B1(n_255),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_29),
.B(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_29),
.A2(n_434),
.B(n_436),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_31),
.Y(n_414)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_32),
.Y(n_157)
);

INVx8_ASAP7_75t_L g435 ( 
.A(n_32),
.Y(n_435)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_38),
.Y(n_416)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_41),
.Y(n_132)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_41),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_41),
.Y(n_357)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_43),
.Y(n_149)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_47),
.B(n_55),
.Y(n_210)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_54),
.B(n_274),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_54),
.A2(n_211),
.B(n_462),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_55),
.B(n_212),
.Y(n_257)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_60),
.A2(n_61),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_61),
.B1(n_99),
.B2(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_89),
.B(n_91),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_62),
.A2(n_268),
.B(n_275),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_62),
.A2(n_89),
.B1(n_303),
.B2(n_348),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_62),
.A2(n_275),
.B(n_348),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_62),
.A2(n_89),
.B1(n_442),
.B2(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_63),
.A2(n_90),
.B1(n_165),
.B2(n_174),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_63),
.A2(n_90),
.B1(n_165),
.B2(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_63),
.A2(n_90),
.B1(n_207),
.B2(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_63),
.B(n_276),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_76),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g246 ( 
.A(n_65),
.Y(n_246)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_67),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_75),
.Y(n_374)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_76),
.A2(n_303),
.B(n_308),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_82),
.Y(n_369)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_82),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_84),
.Y(n_327)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_89),
.A2(n_308),
.B(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_90),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g377 ( 
.A(n_95),
.B(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_97),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_97),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_97),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_97),
.Y(n_444)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_122),
.B1(n_133),
.B2(n_134),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_133),
.B1(n_134),
.B2(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_101),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_101),
.A2(n_133),
.B1(n_178),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_101),
.A2(n_133),
.B1(n_389),
.B2(n_439),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_109),
.B2(n_112),
.Y(n_102)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_103),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_105),
.Y(n_360)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_108),
.Y(n_352)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_108),
.Y(n_410)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_114)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_111),
.Y(n_376)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_123),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

AOI22x1_ASAP7_75t_L g465 ( 
.A1(n_114),
.A2(n_176),
.B1(n_392),
.B2(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_131),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_133),
.B(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_133),
.A2(n_389),
.B(n_391),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_135),
.B(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_138),
.Y(n_361)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_149),
.Y(n_253)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_184),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_160),
.B(n_163),
.CI(n_184),
.CON(n_222),
.SN(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_175),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_176),
.A2(n_351),
.B(n_358),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_176),
.B(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_176),
.A2(n_358),
.B(n_482),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B(n_209),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_206),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_209),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_186),
.A2(n_206),
.B1(n_228),
.B2(n_453),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_193),
.B(n_196),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_196),
.B1(n_235),
.B2(n_242),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_187),
.A2(n_288),
.B(n_293),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_187),
.A2(n_274),
.B(n_293),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_187),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_422)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_188),
.B(n_295),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_188),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_188),
.A2(n_365),
.B1(n_396),
.B2(n_399),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_188),
.A2(n_399),
.B1(n_426),
.B2(n_459),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_189),
.Y(n_329)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_190),
.Y(n_400)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_191),
.Y(n_299)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_202),
.Y(n_298)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_206),
.Y(n_453)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_218),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_258),
.B(n_508),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_222),
.B(n_223),
.Y(n_508)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_222),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.C(n_232),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_229),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_232),
.B(n_468),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_251),
.C(n_254),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_233),
.B(n_451),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_234),
.B(n_244),
.Y(n_476)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_235),
.Y(n_459)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_239),
.Y(n_367)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_242),
.Y(n_337)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_245),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_251),
.B(n_254),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_252),
.Y(n_466)
);

AOI32xp33_ASAP7_75t_L g371 ( 
.A1(n_253),
.A2(n_354),
.A3(n_372),
.B1(n_375),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_257),
.Y(n_436)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI311xp33_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_447),
.A3(n_484),
.B1(n_502),
.C1(n_503),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_403),
.B(n_446),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_380),
.B(n_402),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_342),
.B(n_379),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_311),
.B(n_341),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_286),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_286),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_278),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_267),
.A2(n_278),
.B1(n_279),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_SL g351 ( 
.A1(n_274),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_274),
.B(n_418),
.Y(n_417)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_274),
.A2(n_417),
.B(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_300),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_301),
.C(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_291),
.Y(n_398)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_298),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_309),
.B2(n_310),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_333),
.B(n_340),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_322),
.B(n_332),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_321),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_331),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_331),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_328),
.B(n_330),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_330),
.A2(n_364),
.B(n_370),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_338),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_344),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_362),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_349),
.C(n_362),
.Y(n_381)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx6_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_371),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx5_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_381),
.B(n_382),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_387),
.B2(n_401),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_386),
.C(n_401),
.Y(n_404)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_393),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_394),
.C(n_395),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_404),
.B(n_405),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_431),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_406)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_421),
.B2(n_422),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_409),
.B(n_421),
.Y(n_480)
);

OAI32xp33_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.A3(n_413),
.B1(n_415),
.B2(n_417),
.Y(n_409)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_428),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_428),
.B(n_429),
.C(n_431),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_437),
.B2(n_445),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_432),
.B(n_438),
.C(n_441),
.Y(n_493)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_437),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_441),
.Y(n_437)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_470),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_448),
.A2(n_470),
.B(n_504),
.C(n_507),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_467),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_449),
.B(n_467),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_454),
.Y(n_449)
);

FAx1_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_452),
.CI(n_454),
.CON(n_483),
.SN(n_483)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_460),
.C(n_465),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_458),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_458),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_460),
.A2(n_461),
.B1(n_465),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_483),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_471),
.B(n_483),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_476),
.C(n_477),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_472),
.A2(n_473),
.B1(n_476),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.C(n_481),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_478),
.A2(n_479),
.B1(n_481),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_481),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_483),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_497),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_505),
.B(n_506),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_494),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_494),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_491),
.C(n_493),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_500),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_492),
.B1(n_493),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_493),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_499),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_510),
.Y(n_513)
);

INVx13_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);


endmodule