module fake_jpeg_18165_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_8),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_66),
.Y(n_93)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_75),
.B1(n_65),
.B2(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_92),
.B1(n_59),
.B2(n_64),
.Y(n_102)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_105),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_53),
.B1(n_64),
.B2(n_62),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_102),
.B1(n_107),
.B2(n_61),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_103),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_71),
.C(n_61),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_69),
.B1(n_56),
.B2(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_114),
.B1(n_122),
.B2(n_123),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_49),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_4),
.B(n_5),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_84),
.B1(n_76),
.B2(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_51),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_119),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_0),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_51),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_70),
.C(n_68),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_1),
.C(n_2),
.Y(n_132)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_57),
.B1(n_55),
.B2(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_73),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_50),
.B1(n_17),
.B2(n_24),
.Y(n_125)
);

NAND2x1_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_50),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_135),
.B(n_136),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_7),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_110),
.B(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_142),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_120),
.C(n_31),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_144),
.C(n_139),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_153),
.B(n_149),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_146),
.C(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_148),
.B1(n_146),
.B2(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_34),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_32),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_37),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_29),
.B(n_11),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_40),
.B(n_12),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_41),
.C(n_13),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_25),
.A3(n_26),
.B1(n_46),
.B2(n_124),
.C(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_131),
.Y(n_165)
);


endmodule