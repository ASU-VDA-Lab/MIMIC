module fake_netlist_1_7849_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_1), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
CKINVDCx16_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
NAND2x1_ASAP7_75t_L g18 ( .A(n_15), .B(n_0), .Y(n_18) );
OAI22xp33_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_14), .B1(n_13), .B2(n_17), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_11), .A2(n_6), .B(n_7), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_12), .B(n_1), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
NAND2xp33_ASAP7_75t_R g25 ( .A(n_20), .B(n_3), .Y(n_25) );
BUFx12f_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_18), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVxp67_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_24), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
OAI33xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_18), .A3(n_26), .B1(n_22), .B2(n_4), .B3(n_5), .Y(n_32) );
NAND4xp25_ASAP7_75t_L g33 ( .A(n_31), .B(n_30), .C(n_28), .D(n_26), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVx2_ASAP7_75t_SL g35 ( .A(n_34), .Y(n_35) );
XNOR2xp5_ASAP7_75t_L g36 ( .A(n_33), .B(n_26), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_12), .B1(n_21), .B2(n_3), .Y(n_37) );
OAI211xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_5), .B(n_12), .C(n_33), .Y(n_38) );
AOI22xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_12), .B1(n_35), .B2(n_37), .Y(n_39) );
endmodule