module fake_jpeg_20531_n_31 (n_3, n_2, n_1, n_0, n_4, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_SL g5 ( 
.A(n_1),
.B(n_4),
.Y(n_5)
);

BUFx5_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_3),
.B(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_4),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_12),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_14),
.B1(n_5),
.B2(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_6),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_15),
.A2(n_16),
.B(n_18),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_9),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_5),
.B(n_12),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_15),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_25),
.C(n_20),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_15),
.B1(n_10),
.B2(n_9),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AO221x1_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_2),
.B1(n_10),
.B2(n_14),
.C(n_23),
.Y(n_31)
);


endmodule