module fake_jpeg_13288_n_68 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_14),
.B1(n_9),
.B2(n_12),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_22),
.B1(n_26),
.B2(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

NAND2x1_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_33),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_14),
.B1(n_12),
.B2(n_19),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_18),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_41),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_42),
.B(n_35),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_25),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_30),
.C(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_39),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_15),
.C(n_19),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_50),
.B1(n_46),
.B2(n_34),
.Y(n_58)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_60),
.B(n_36),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_47),
.C(n_49),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_61),
.C(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_63),
.B(n_13),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_54),
.C(n_15),
.Y(n_63)
);

AOI21x1_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_37),
.B(n_23),
.Y(n_66)
);

OAI31xp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_66),
.A3(n_6),
.B(n_2),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_1),
.C(n_3),
.Y(n_68)
);


endmodule