module fake_jpeg_716_n_529 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_529);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_529;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_434;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_49),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_51),
.B(n_57),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_95),
.Y(n_106)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_53),
.Y(n_163)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_63),
.B(n_64),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_70),
.B(n_74),
.Y(n_130)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_71),
.Y(n_164)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_17),
.B(n_6),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_92),
.Y(n_112)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_6),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_6),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_37),
.B(n_5),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_23),
.Y(n_117)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

BUFx16f_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_58),
.B(n_93),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_103),
.B(n_40),
.C(n_99),
.Y(n_195)
);

INVx2_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_104),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_117),
.B(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_23),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_19),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_127),
.B(n_128),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_19),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_47),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_55),
.B(n_39),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_144),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_82),
.B(n_47),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_45),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_31),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_46),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_71),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_69),
.A2(n_31),
.B1(n_39),
.B2(n_45),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_40),
.B1(n_48),
.B2(n_32),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_50),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_48),
.B1(n_40),
.B2(n_42),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_167),
.B(n_195),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_168),
.B(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_59),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_169),
.B(n_170),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_96),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_90),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_172),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_67),
.B1(n_94),
.B2(n_87),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_174),
.A2(n_198),
.B1(n_164),
.B2(n_155),
.Y(n_229)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_178),
.A2(n_190),
.B1(n_211),
.B2(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_86),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_117),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_181),
.B(n_188),
.Y(n_233)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_86),
.Y(n_188)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_38),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_192),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_106),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_53),
.B1(n_152),
.B2(n_108),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_210),
.Y(n_247)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_106),
.A2(n_32),
.B1(n_25),
.B2(n_42),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_107),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_136),
.A2(n_32),
.B1(n_25),
.B2(n_42),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_48),
.B1(n_25),
.B2(n_41),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_194),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_116),
.C(n_145),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_172),
.C(n_166),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_174),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_189),
.B1(n_212),
.B2(n_178),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_177),
.A2(n_104),
.B(n_154),
.C(n_41),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_246),
.B(n_232),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_173),
.A2(n_151),
.B1(n_118),
.B2(n_125),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_210),
.B1(n_139),
.B2(n_124),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_137),
.B1(n_88),
.B2(n_68),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_171),
.B1(n_199),
.B2(n_185),
.Y(n_253)
);

OAI22x1_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_129),
.B1(n_110),
.B2(n_131),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_198),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_230),
.C(n_187),
.Y(n_292)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_254),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_227),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_196),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_263),
.Y(n_304)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_257),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_206),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_259),
.B(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

OR2x2_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_175),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_274),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_222),
.A2(n_196),
.B1(n_173),
.B2(n_172),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_239),
.B1(n_249),
.B2(n_224),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_222),
.A2(n_198),
.B1(n_137),
.B2(n_125),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_268),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_222),
.A2(n_184),
.B(n_180),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_267),
.A2(n_241),
.B(n_250),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_182),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_235),
.B(n_175),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_272),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_203),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

OR2x2_ASAP7_75t_SL g274 ( 
.A(n_233),
.B(n_219),
.Y(n_274)
);

BUFx16f_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_189),
.Y(n_313)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_280),
.Y(n_288)
);

BUFx4f_ASAP7_75t_SL g281 ( 
.A(n_248),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_236),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_229),
.B1(n_243),
.B2(n_215),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_306),
.B1(n_265),
.B2(n_253),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_305),
.C(n_273),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_267),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_269),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_219),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_309),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_307),
.B(n_258),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_254),
.C(n_261),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_198),
.B1(n_124),
.B2(n_139),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_241),
.B(n_250),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_308),
.A2(n_252),
.B1(n_281),
.B2(n_262),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_249),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_189),
.B(n_248),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_275),
.B(n_260),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_238),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_256),
.B1(n_259),
.B2(n_270),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_315),
.A2(n_334),
.B1(n_301),
.B2(n_288),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_284),
.B(n_274),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_316),
.B(n_340),
.C(n_333),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_263),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_336),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_341),
.B1(n_345),
.B2(n_289),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_275),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_SL g350 ( 
.A(n_319),
.B(n_338),
.C(n_299),
.Y(n_350)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_310),
.B(n_307),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_322),
.B(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_323),
.Y(n_361)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_339),
.C(n_286),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_255),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_313),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_310),
.B(n_307),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_289),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_278),
.Y(n_333)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_301),
.A2(n_260),
.B1(n_277),
.B2(n_264),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_238),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_281),
.Y(n_337)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_R g338 ( 
.A1(n_304),
.A2(n_257),
.B1(n_281),
.B2(n_244),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_234),
.C(n_150),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_262),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_343),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_295),
.B(n_234),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_217),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_286),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_290),
.A2(n_224),
.B1(n_220),
.B2(n_257),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_284),
.B(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_292),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_355),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_352),
.C(n_363),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_282),
.C(n_302),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_356),
.B(n_357),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_288),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_327),
.A2(n_298),
.B(n_287),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_360),
.A2(n_367),
.B(n_319),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_331),
.B1(n_342),
.B2(n_343),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_297),
.C(n_309),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_318),
.A2(n_290),
.B1(n_287),
.B2(n_306),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_364),
.A2(n_220),
.B1(n_204),
.B2(n_197),
.Y(n_405)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_306),
.Y(n_368)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_293),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_371),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_314),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_375),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_314),
.B(n_283),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_283),
.B(n_308),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_326),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_361),
.A2(n_334),
.B1(n_315),
.B2(n_366),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_380),
.A2(n_381),
.B1(n_391),
.B2(n_394),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_340),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_363),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_390),
.A2(n_405),
.B1(n_379),
.B2(n_359),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_368),
.A2(n_345),
.B1(n_321),
.B2(n_326),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_402),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_335),
.B1(n_332),
.B2(n_330),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_320),
.Y(n_395)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_395),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_291),
.Y(n_396)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_396),
.Y(n_415)
);

BUFx12_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_365),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_403),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_209),
.C(n_236),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_407),
.C(n_360),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_355),
.B(n_201),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_400),
.B(n_409),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_214),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_358),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_214),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_393),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_358),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_376),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_142),
.C(n_183),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_408),
.B(n_372),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_356),
.B(n_221),
.Y(n_409)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_434),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_428),
.B1(n_397),
.B2(n_190),
.Y(n_449)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_422),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_383),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_420),
.Y(n_456)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_421),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_385),
.B(n_357),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_401),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_424),
.Y(n_444)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_379),
.C(n_367),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_425),
.B(n_426),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_364),
.C(n_354),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_359),
.C(n_377),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_430),
.B(n_431),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_377),
.C(n_347),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_433),
.B(n_415),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_402),
.C(n_404),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_438),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_407),
.C(n_392),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_409),
.C(n_400),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_446),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_429),
.A2(n_387),
.B(n_390),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_391),
.C(n_387),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_448),
.Y(n_470)
);

OAI322xp33_ASAP7_75t_L g448 ( 
.A1(n_427),
.A2(n_397),
.A3(n_347),
.B1(n_221),
.B2(n_217),
.C1(n_176),
.C2(n_202),
.Y(n_448)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_138),
.C(n_121),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_452),
.C(n_455),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_105),
.C(n_148),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_414),
.Y(n_453)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_193),
.C(n_77),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_413),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_458),
.B(n_462),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_436),
.A2(n_411),
.B(n_422),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_461),
.B(n_465),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_432),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_416),
.C(n_56),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_453),
.A2(n_416),
.B(n_27),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_466),
.B(n_8),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_444),
.A2(n_155),
.B1(n_61),
.B2(n_158),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_467),
.A2(n_468),
.B1(n_472),
.B2(n_43),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_445),
.A2(n_158),
.B1(n_129),
.B2(n_134),
.Y(n_468)
);

FAx1_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_163),
.CI(n_134),
.CON(n_472),
.SN(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_134),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_452),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_438),
.A2(n_27),
.B(n_21),
.Y(n_474)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_440),
.A2(n_27),
.B1(n_21),
.B2(n_158),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_475),
.A2(n_474),
.B1(n_472),
.B2(n_466),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_460),
.B(n_442),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_477),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_456),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_457),
.B(n_451),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_482),
.Y(n_497)
);

OAI22x1_ASAP7_75t_L g479 ( 
.A1(n_471),
.A2(n_470),
.B1(n_472),
.B2(n_469),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_483),
.B1(n_489),
.B2(n_492),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_481),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_441),
.C(n_455),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_463),
.A2(n_454),
.B1(n_450),
.B2(n_21),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_160),
.C(n_43),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_485),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_43),
.C(n_20),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_475),
.B(n_11),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_486),
.B(n_468),
.Y(n_496)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_487),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_20),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_18),
.C(n_8),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_501),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_480),
.A2(n_459),
.B(n_467),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_498),
.A2(n_503),
.B(n_505),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_459),
.B(n_20),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_500),
.A2(n_2),
.B(n_3),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_18),
.C(n_5),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_502),
.B(n_0),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_14),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_479),
.A2(n_481),
.B(n_484),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g506 ( 
.A1(n_494),
.A2(n_487),
.A3(n_490),
.B1(n_485),
.B2(n_3),
.C1(n_4),
.C2(n_11),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_507),
.Y(n_519)
);

FAx1_ASAP7_75t_SL g507 ( 
.A(n_499),
.B(n_4),
.CI(n_13),
.CON(n_507),
.SN(n_507)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_508),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_509),
.A2(n_511),
.B(n_503),
.Y(n_516)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_2),
.B(n_4),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_2),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_512),
.B(n_514),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_4),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_516),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_513),
.A2(n_493),
.B(n_12),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_520),
.B(n_12),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_510),
.A2(n_493),
.B(n_507),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_506),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_521),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_515),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g526 ( 
.A1(n_524),
.A2(n_1),
.A3(n_13),
.B1(n_14),
.B2(n_518),
.C1(n_522),
.C2(n_525),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_14),
.B(n_1),
.Y(n_527)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_527),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_528),
.Y(n_529)
);


endmodule