module fake_jpeg_15892_n_288 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_29),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_23),
.B1(n_22),
.B2(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_36),
.B1(n_22),
.B2(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_66),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_23),
.B1(n_36),
.B2(n_22),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_15),
.B1(n_21),
.B2(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_15),
.B1(n_21),
.B2(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_39),
.Y(n_78)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_43),
.B1(n_44),
.B2(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_76),
.B1(n_63),
.B2(n_73),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_21),
.B1(n_24),
.B2(n_28),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_86),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_45),
.C(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_96),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_45),
.C(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_95),
.Y(n_104)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_18),
.B(n_29),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_39),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_45),
.C(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_108),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_109),
.B1(n_99),
.B2(n_79),
.Y(n_134)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_74),
.B1(n_59),
.B2(n_71),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_67),
.B(n_26),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_129),
.B(n_20),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_38),
.B1(n_39),
.B2(n_62),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_117),
.Y(n_138)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_119),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_18),
.C(n_28),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_88),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_57),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_81),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_32),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_90),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_20),
.B(n_32),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_130),
.A2(n_142),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_145),
.B1(n_147),
.B2(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_135),
.B(n_17),
.Y(n_178)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_86),
.C(n_97),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_132),
.C(n_151),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_92),
.C(n_94),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_98),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_96),
.B1(n_63),
.B2(n_76),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_92),
.B1(n_99),
.B2(n_79),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_111),
.B(n_112),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_34),
.B1(n_71),
.B2(n_59),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_26),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_34),
.B1(n_74),
.B2(n_30),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_34),
.B1(n_38),
.B2(n_25),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_157),
.B1(n_159),
.B2(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_106),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_25),
.B1(n_10),
.B2(n_13),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_138),
.B(n_133),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_186),
.B(n_133),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_113),
.B1(n_112),
.B2(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_173),
.C(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_178),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_146),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_156),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_116),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_128),
.C(n_48),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_181),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_188),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_105),
.B1(n_128),
.B2(n_2),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_69),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_167),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_195),
.C(n_201),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_171),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_140),
.C(n_154),
.Y(n_195)
);

OAI22x1_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_130),
.B1(n_153),
.B2(n_159),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_208),
.B1(n_176),
.B2(n_172),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_130),
.B(n_158),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_199),
.B(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_128),
.Y(n_201)
);

XOR2x2_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_17),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_69),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_175),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_0),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_165),
.B1(n_169),
.B2(n_180),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_206),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_193),
.C(n_201),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_219),
.C(n_224),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_177),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_174),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_199),
.C(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_200),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_165),
.C(n_180),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_222),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_169),
.B1(n_163),
.B2(n_184),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_227),
.B1(n_208),
.B2(n_192),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_161),
.C(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_163),
.B1(n_10),
.B2(n_11),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_226),
.A2(n_205),
.B1(n_191),
.B2(n_203),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_38),
.B1(n_9),
.B2(n_7),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_204),
.B(n_198),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_213),
.B1(n_212),
.B2(n_9),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_220),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_192),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_211),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_38),
.B1(n_50),
.B2(n_7),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_48),
.C(n_26),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_26),
.C(n_17),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_8),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_0),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_232),
.C(n_240),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_216),
.B(n_219),
.C(n_221),
.D(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_252),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_253),
.B(n_10),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_230),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_262),
.B(n_251),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_230),
.B(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_6),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_256),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_50),
.C(n_2),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_253),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_263),
.B(n_260),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_268),
.B(n_270),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_5),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_6),
.B(n_12),
.Y(n_268)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_6),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_7),
.B(n_12),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_4),
.B(n_11),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_277),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_13),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_279),
.B1(n_274),
.B2(n_12),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_1),
.B(n_2),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_1),
.B(n_3),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_1),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_3),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_287),
.Y(n_288)
);


endmodule