module fake_netlist_6_3410_n_1033 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1033);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1033;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_953;
wire n_448;
wire n_844;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_970;
wire n_849;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_1001;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g224 ( 
.A(n_49),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_165),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_149),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_107),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_114),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_201),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_81),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_109),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_113),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_112),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_31),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_181),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_177),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_128),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_3),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_27),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_108),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_31),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_211),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_192),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_53),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_58),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_189),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_14),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_56),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_39),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_12),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_171),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_134),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_191),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_220),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_219),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_188),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_16),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_45),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_141),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_44),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_48),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_222),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_102),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_218),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_144),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_69),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_71),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_90),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_94),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_133),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_6),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_203),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_3),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_169),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_98),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_46),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_21),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_156),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_62),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_153),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_18),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_67),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_166),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_93),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_215),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_150),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_70),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_172),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_30),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_99),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_106),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_163),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_66),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_184),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_221),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_225),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_300),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_266),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_241),
.B(n_0),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_241),
.B(n_0),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_236),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_1),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_243),
.B(n_2),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_266),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_275),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_245),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_303),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_257),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_226),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_270),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_275),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_259),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_227),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_251),
.B(n_2),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_224),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_251),
.B(n_4),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_308),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_235),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_239),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_268),
.B(n_5),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_5),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_295),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_230),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_240),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_244),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_230),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_231),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_228),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_250),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_252),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_258),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_246),
.B(n_6),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_231),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_329),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_334),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_318),
.B(n_287),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_322),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_278),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_246),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_256),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_286),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_256),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_329),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_360),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_277),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_277),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_294),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_337),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_358),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_248),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_361),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_361),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_261),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_325),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_R g412 ( 
.A(n_325),
.B(n_232),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_347),
.A2(n_291),
.B(n_297),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_R g415 ( 
.A(n_330),
.B(n_232),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_330),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_341),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_338),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_319),
.B(n_291),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_350),
.B(n_307),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_357),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_337),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_331),
.B(n_316),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_343),
.B(n_234),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_425),
.B(n_282),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_402),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_356),
.C(n_355),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_427),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_426),
.A2(n_368),
.B1(n_324),
.B2(n_321),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_382),
.B(n_379),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_401),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_281),
.B1(n_315),
.B2(n_326),
.Y(n_442)
);

BUFx4f_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_344),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_392),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_413),
.A2(n_327),
.B1(n_346),
.B2(n_282),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_425),
.B(n_305),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_401),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_425),
.B(n_305),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_425),
.B(n_305),
.Y(n_455)
);

INVx8_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_395),
.Y(n_457)
);

CKINVDCx8_ASAP7_75t_R g458 ( 
.A(n_427),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_386),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_305),
.B1(n_294),
.B2(n_233),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_233),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_317),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_237),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_317),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_381),
.B(n_238),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_242),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_375),
.B(n_247),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_414),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_348),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_381),
.B(n_249),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_253),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_377),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_406),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_374),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_394),
.B(n_260),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_417),
.B(n_262),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_417),
.B(n_263),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_377),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_402),
.B(n_264),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_402),
.B(n_265),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_377),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_269),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_271),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_419),
.B(n_272),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_396),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_430),
.B(n_274),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_411),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_276),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_413),
.A2(n_294),
.B1(n_279),
.B2(n_301),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_400),
.B(n_280),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_404),
.B(n_284),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_439),
.A2(n_410),
.B1(n_423),
.B2(n_416),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_503),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_495),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_503),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_L g513 ( 
.A(n_451),
.B(n_410),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_507),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_457),
.B(n_376),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_450),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_416),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_495),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_463),
.B(n_423),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_451),
.A2(n_378),
.B(n_404),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_465),
.B(n_407),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_462),
.B(n_407),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_408),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_453),
.B(n_408),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_461),
.A2(n_348),
.B1(n_352),
.B2(n_296),
.Y(n_530)
);

AND2x6_ASAP7_75t_SL g531 ( 
.A(n_472),
.B(n_320),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_507),
.A2(n_320),
.B1(n_328),
.B2(n_352),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_463),
.A2(n_412),
.B1(n_415),
.B2(n_314),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_505),
.B(n_289),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_464),
.B(n_398),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_471),
.B(n_292),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_461),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_502),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_471),
.B(n_397),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_474),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_483),
.B(n_373),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_504),
.B(n_398),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_505),
.B(n_434),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_299),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_460),
.B(n_304),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_442),
.A2(n_478),
.B1(n_480),
.B2(n_479),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_470),
.B(n_306),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_443),
.A2(n_311),
.B(n_309),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_482),
.B(n_40),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_L g552 ( 
.A(n_475),
.B(n_312),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_456),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_449),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_486),
.B(n_313),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_485),
.B(n_328),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_L g558 ( 
.A(n_435),
.B(n_428),
.C(n_388),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_438),
.B(n_41),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_489),
.B(n_373),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_488),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_469),
.A2(n_428),
.B(n_403),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_468),
.A2(n_403),
.B1(n_388),
.B2(n_9),
.Y(n_564)
);

AND2x6_ASAP7_75t_SL g565 ( 
.A(n_458),
.B(n_7),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_498),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_492),
.B(n_500),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_456),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_438),
.B(n_42),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_477),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_499),
.B(n_47),
.Y(n_571)
);

O2A1O1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_468),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_473),
.B(n_10),
.Y(n_573)
);

AND2x6_ASAP7_75t_SL g574 ( 
.A(n_502),
.B(n_483),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_506),
.B(n_50),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_487),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_473),
.B(n_10),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_484),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_506),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_456),
.B(n_11),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_490),
.B(n_51),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_443),
.B(n_52),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_477),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_497),
.B(n_13),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_491),
.B(n_496),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_432),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_433),
.B(n_54),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_432),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_540),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_568),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_516),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_509),
.B(n_497),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_538),
.B(n_433),
.Y(n_594)
);

O2A1O1Ixp5_ASAP7_75t_L g595 ( 
.A1(n_545),
.A2(n_455),
.B(n_452),
.C(n_454),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_586),
.A2(n_493),
.B(n_444),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_536),
.A2(n_493),
.B(n_444),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_578),
.B(n_526),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_521),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_554),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_508),
.B(n_454),
.C(n_452),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_515),
.A2(n_501),
.B(n_494),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_545),
.A2(n_455),
.B(n_501),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_554),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_513),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_523),
.A2(n_514),
.B1(n_549),
.B2(n_528),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_543),
.A2(n_494),
.B(n_459),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_527),
.A2(n_494),
.B1(n_459),
.B2(n_437),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_512),
.B(n_437),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_525),
.A2(n_459),
.B(n_437),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_549),
.B(n_517),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_530),
.B(n_15),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_534),
.A2(n_119),
.B1(n_216),
.B2(n_212),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_117),
.B(n_210),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_567),
.A2(n_116),
.B(n_209),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_567),
.A2(n_115),
.B(n_208),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_537),
.B(n_17),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_559),
.A2(n_569),
.B1(n_587),
.B2(n_589),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_529),
.B(n_17),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_535),
.A2(n_118),
.B(n_207),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_537),
.B(n_552),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_580),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_524),
.B(n_18),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_529),
.A2(n_111),
.B1(n_206),
.B2(n_204),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_556),
.A2(n_582),
.B(n_581),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_535),
.A2(n_575),
.B(n_548),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_581),
.A2(n_110),
.B(n_202),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_541),
.Y(n_631)
);

OA22x2_ASAP7_75t_L g632 ( 
.A1(n_563),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_510),
.Y(n_633)
);

OAI21xp33_ASAP7_75t_L g634 ( 
.A1(n_573),
.A2(n_19),
.B(n_22),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_573),
.B(n_23),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_544),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_584),
.A2(n_120),
.B(n_200),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_577),
.B(n_23),
.C(n_24),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_551),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_577),
.B(n_25),
.C(n_26),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_584),
.A2(n_121),
.B(n_199),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_544),
.B(n_25),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_583),
.A2(n_122),
.B(n_198),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_531),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_511),
.B(n_26),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_583),
.A2(n_105),
.B(n_196),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_585),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_518),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_562),
.A2(n_123),
.B(n_195),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_557),
.B(n_28),
.C(n_29),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_518),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_592),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g653 ( 
.A1(n_606),
.A2(n_564),
.B(n_557),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_611),
.B(n_561),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_594),
.A2(n_628),
.B(n_619),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_595),
.A2(n_585),
.B(n_566),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_599),
.Y(n_657)
);

OAI22x1_ASAP7_75t_L g658 ( 
.A1(n_612),
.A2(n_621),
.B1(n_644),
.B2(n_561),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_598),
.B(n_522),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_590),
.Y(n_660)
);

OAI21xp33_ASAP7_75t_SL g661 ( 
.A1(n_635),
.A2(n_539),
.B(n_547),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_593),
.B(n_542),
.Y(n_662)
);

OA21x2_ASAP7_75t_L g663 ( 
.A1(n_603),
.A2(n_562),
.B(n_566),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_633),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_623),
.B(n_551),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_596),
.A2(n_588),
.B(n_546),
.Y(n_666)
);

OA21x2_ASAP7_75t_L g667 ( 
.A1(n_610),
.A2(n_576),
.B(n_533),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_627),
.A2(n_533),
.B(n_560),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_618),
.A2(n_572),
.B(n_579),
.C(n_547),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_602),
.A2(n_597),
.B(n_607),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_624),
.B(n_617),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_642),
.Y(n_672)
);

AOI21x1_ASAP7_75t_L g673 ( 
.A1(n_648),
.A2(n_555),
.B(n_571),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_629),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_620),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_629),
.B(n_639),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_629),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_639),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_645),
.B(n_532),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_553),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_622),
.A2(n_571),
.B(n_550),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_643),
.A2(n_579),
.B(n_558),
.Y(n_682)
);

AOI21xp33_ASAP7_75t_L g683 ( 
.A1(n_634),
.A2(n_574),
.B(n_32),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_631),
.B(n_30),
.Y(n_684)
);

AOI21x1_ASAP7_75t_L g685 ( 
.A1(n_651),
.A2(n_126),
.B(n_223),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_625),
.Y(n_686)
);

AOI221xp5_ASAP7_75t_L g687 ( 
.A1(n_647),
.A2(n_565),
.B1(n_33),
.B2(n_34),
.C(n_35),
.Y(n_687)
);

OAI21xp33_ASAP7_75t_L g688 ( 
.A1(n_650),
.A2(n_32),
.B(n_33),
.Y(n_688)
);

OAI21x1_ASAP7_75t_SL g689 ( 
.A1(n_646),
.A2(n_605),
.B(n_616),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_601),
.A2(n_124),
.B(n_190),
.Y(n_690)
);

INVx6_ASAP7_75t_L g691 ( 
.A(n_600),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_609),
.A2(n_608),
.B(n_624),
.Y(n_692)
);

AO31x2_ASAP7_75t_L g693 ( 
.A1(n_613),
.A2(n_34),
.A3(n_35),
.B(n_36),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_638),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_636),
.B(n_55),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_615),
.A2(n_129),
.B(n_187),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_640),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_698)
);

BUFx4_ASAP7_75t_SL g699 ( 
.A(n_591),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_600),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_649),
.A2(n_57),
.B(n_59),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_614),
.A2(n_60),
.B(n_61),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_630),
.A2(n_63),
.B(n_64),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_636),
.B(n_65),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_641),
.A2(n_68),
.B(n_72),
.C(n_73),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_626),
.A2(n_74),
.B(n_75),
.Y(n_706)
);

AOI21xp33_ASAP7_75t_L g707 ( 
.A1(n_600),
.A2(n_76),
.B(n_78),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_706),
.A2(n_637),
.B(n_604),
.C(n_82),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_655),
.A2(n_604),
.B(n_80),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_704),
.B(n_79),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_654),
.B(n_83),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_653),
.B(n_662),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_686),
.B(n_84),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_679),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_652),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_687),
.B(n_88),
.C(n_89),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_699),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_671),
.B(n_91),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_665),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_675),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_694),
.B(n_97),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_672),
.B(n_100),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_688),
.A2(n_103),
.B1(n_104),
.B2(n_127),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_659),
.B(n_130),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_687),
.B(n_131),
.C(n_135),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_700),
.B(n_136),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_657),
.B(n_137),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_655),
.A2(n_138),
.B(n_139),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_SL g731 ( 
.A(n_690),
.B(n_140),
.C(n_142),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_660),
.B(n_143),
.Y(n_732)
);

CKINVDCx11_ASAP7_75t_R g733 ( 
.A(n_699),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_669),
.A2(n_146),
.B(n_148),
.C(n_152),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_695),
.A2(n_154),
.B(n_155),
.C(n_157),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_658),
.B(n_158),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_691),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_691),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_691),
.B(n_159),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_683),
.B(n_160),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_674),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_700),
.B(n_162),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_674),
.B(n_194),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_677),
.B(n_164),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_677),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_678),
.B(n_167),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_SL g747 ( 
.A1(n_698),
.A2(n_170),
.B(n_173),
.C(n_174),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_SL g748 ( 
.A1(n_697),
.A2(n_175),
.B(n_176),
.C(n_178),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_678),
.B(n_179),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_676),
.B(n_186),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_680),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_682),
.A2(n_661),
.B(n_689),
.C(n_656),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_682),
.B(n_180),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_681),
.A2(n_182),
.B(n_183),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_663),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_681),
.A2(n_185),
.B(n_666),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_668),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_663),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_692),
.B(n_696),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_758),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_737),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_712),
.B(n_693),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_743),
.B(n_692),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_716),
.A2(n_707),
.B1(n_702),
.B2(n_703),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_715),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_739),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_720),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_724),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_730),
.A2(n_666),
.B1(n_673),
.B2(n_670),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_723),
.A2(n_670),
.B1(n_705),
.B2(n_667),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_757),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_745),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_751),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_741),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_756),
.A2(n_752),
.B(n_759),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_741),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_739),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_718),
.B(n_667),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_721),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_718),
.B(n_693),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_711),
.B(n_693),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_738),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_733),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_743),
.B(n_701),
.Y(n_784)
);

BUFx8_ASAP7_75t_SL g785 ( 
.A(n_717),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_749),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_710),
.A2(n_726),
.B1(n_731),
.B2(n_740),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_756),
.A2(n_685),
.B(n_705),
.Y(n_788)
);

BUFx12f_ASAP7_75t_L g789 ( 
.A(n_739),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_744),
.Y(n_790)
);

CKINVDCx11_ASAP7_75t_R g791 ( 
.A(n_727),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_752),
.A2(n_708),
.B(n_709),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_746),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_731),
.A2(n_723),
.B1(n_736),
.B2(n_753),
.Y(n_794)
);

AO21x1_ASAP7_75t_L g795 ( 
.A1(n_734),
.A2(n_735),
.B(n_729),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_750),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_755),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_750),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_732),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_755),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_713),
.A2(n_722),
.B1(n_728),
.B2(n_725),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_714),
.A2(n_719),
.B1(n_729),
.B2(n_754),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_742),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_754),
.B(n_734),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_747),
.Y(n_806)
);

AO21x1_ASAP7_75t_L g807 ( 
.A1(n_735),
.A2(n_635),
.B(n_712),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_748),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_712),
.A2(n_612),
.B1(n_687),
.B2(n_650),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_718),
.B(n_629),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_724),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_712),
.A2(n_612),
.B1(n_687),
.B2(n_650),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_758),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_715),
.Y(n_814)
);

AOI21x1_ASAP7_75t_L g815 ( 
.A1(n_709),
.A2(n_681),
.B(n_756),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_758),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_756),
.A2(n_665),
.B(n_681),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_760),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_760),
.B(n_813),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_813),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_816),
.Y(n_821)
);

AO21x2_ASAP7_75t_L g822 ( 
.A1(n_792),
.A2(n_775),
.B(n_817),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_816),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_771),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_762),
.B(n_801),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_797),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_801),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_815),
.A2(n_788),
.B(n_769),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_781),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_766),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_773),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_778),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_765),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_780),
.B(n_805),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_789),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_763),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_767),
.Y(n_837)
);

AO21x2_ASAP7_75t_L g838 ( 
.A1(n_795),
.A2(n_770),
.B(n_788),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_814),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_778),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_763),
.B(n_786),
.Y(n_841)
);

AO21x1_ASAP7_75t_SL g842 ( 
.A1(n_787),
.A2(n_794),
.B(n_803),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_763),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_805),
.B(n_777),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_784),
.B(n_766),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_779),
.B(n_772),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_784),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_794),
.B(n_784),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_774),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_776),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_768),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_806),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_764),
.A2(n_803),
.B(n_808),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_789),
.Y(n_854)
);

BUFx8_ASAP7_75t_SL g855 ( 
.A(n_785),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_806),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_806),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_796),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_807),
.Y(n_860)
);

CKINVDCx14_ASAP7_75t_R g861 ( 
.A(n_783),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_825),
.B(n_811),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_824),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_825),
.B(n_848),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_824),
.Y(n_865)
);

BUFx2_ASAP7_75t_SL g866 ( 
.A(n_835),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_825),
.B(n_848),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_829),
.B(n_793),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_818),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_848),
.B(n_790),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_829),
.B(n_800),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_841),
.B(n_800),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_819),
.B(n_809),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_841),
.B(n_804),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_820),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_841),
.B(n_804),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_832),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_847),
.B(n_799),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_821),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_847),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_821),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_819),
.B(n_812),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_826),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_834),
.B(n_766),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_834),
.B(n_777),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_832),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_847),
.B(n_799),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_843),
.B(n_777),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_823),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_819),
.B(n_809),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_860),
.Y(n_891)
);

OAI22xp33_ASAP7_75t_L g892 ( 
.A1(n_860),
.A2(n_812),
.B1(n_798),
.B2(n_802),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_836),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_862),
.B(n_851),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_864),
.B(n_843),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_862),
.B(n_851),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_870),
.B(n_831),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_870),
.B(n_831),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_871),
.B(n_846),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_892),
.A2(n_842),
.B1(n_836),
.B2(n_845),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_864),
.B(n_843),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_867),
.B(n_832),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_892),
.B(n_834),
.C(n_859),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_867),
.B(n_840),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_871),
.B(n_846),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_874),
.B(n_876),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_SL g907 ( 
.A1(n_873),
.A2(n_861),
.B(n_845),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_874),
.B(n_846),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_876),
.B(n_837),
.Y(n_909)
);

OA211x2_ASAP7_75t_L g910 ( 
.A1(n_873),
.A2(n_764),
.B(n_842),
.C(n_835),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_880),
.B(n_840),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_880),
.B(n_836),
.Y(n_912)
);

OAI221xp5_ASAP7_75t_L g913 ( 
.A1(n_882),
.A2(n_854),
.B1(n_835),
.B2(n_890),
.C(n_885),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_SL g914 ( 
.A1(n_891),
.A2(n_858),
.B(n_857),
.Y(n_914)
);

OAI21xp33_ASAP7_75t_L g915 ( 
.A1(n_882),
.A2(n_853),
.B(n_859),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_880),
.B(n_836),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_890),
.A2(n_853),
.B(n_859),
.Y(n_917)
);

INVxp67_ASAP7_75t_SL g918 ( 
.A(n_911),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_897),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_895),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_902),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_898),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_894),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_902),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_895),
.B(n_893),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_896),
.B(n_872),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_909),
.B(n_872),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_901),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_901),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_899),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_912),
.B(n_893),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_905),
.B(n_887),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_906),
.B(n_887),
.Y(n_933)
);

NAND2x1_ASAP7_75t_L g934 ( 
.A(n_931),
.B(n_904),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_920),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_920),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_928),
.B(n_893),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_931),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_923),
.B(n_913),
.C(n_903),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_932),
.B(n_908),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_919),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_926),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_931),
.B(n_928),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_935),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_935),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_941),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_939),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_942),
.B(n_930),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_936),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_934),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_936),
.Y(n_951)
);

OAI22xp33_ASAP7_75t_SL g952 ( 
.A1(n_937),
.A2(n_930),
.B1(n_922),
.B2(n_918),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_950),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_945),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_946),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_945),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_947),
.B(n_855),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_957),
.B(n_947),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_956),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_955),
.A2(n_907),
.B1(n_938),
.B2(n_948),
.Y(n_960)
);

AOI322xp5_ASAP7_75t_L g961 ( 
.A1(n_957),
.A2(n_900),
.A3(n_915),
.B1(n_917),
.B2(n_949),
.C1(n_951),
.C2(n_944),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_959),
.B(n_953),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_958),
.B(n_954),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_960),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_961),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_959),
.Y(n_966)
);

AOI21xp33_ASAP7_75t_SL g967 ( 
.A1(n_965),
.A2(n_952),
.B(n_761),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_966),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_963),
.B(n_956),
.C(n_782),
.Y(n_969)
);

OAI221xp5_ASAP7_75t_L g970 ( 
.A1(n_964),
.A2(n_854),
.B1(n_866),
.B2(n_940),
.C(n_914),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_SL g971 ( 
.A1(n_962),
.A2(n_933),
.B(n_921),
.Y(n_971)
);

NAND4xp25_ASAP7_75t_SL g972 ( 
.A(n_965),
.B(n_783),
.C(n_785),
.D(n_904),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_965),
.A2(n_853),
.B(n_943),
.Y(n_973)
);

OAI211xp5_ASAP7_75t_SL g974 ( 
.A1(n_965),
.A2(n_791),
.B(n_927),
.C(n_884),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_SL g975 ( 
.A1(n_963),
.A2(n_854),
.B(n_782),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_968),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_969),
.B(n_791),
.C(n_839),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_973),
.Y(n_978)
);

NAND5xp2_ASAP7_75t_L g979 ( 
.A(n_970),
.B(n_810),
.C(n_910),
.D(n_833),
.E(n_837),
.Y(n_979)
);

AND2x2_ASAP7_75t_SL g980 ( 
.A(n_972),
.B(n_943),
.Y(n_980)
);

NAND5xp2_ASAP7_75t_L g981 ( 
.A(n_975),
.B(n_810),
.C(n_910),
.D(n_839),
.E(n_833),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_925),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_925),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_976),
.B(n_974),
.C(n_830),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_L g985 ( 
.A(n_977),
.B(n_830),
.C(n_868),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_978),
.B(n_929),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_977),
.B(n_830),
.Y(n_987)
);

NOR4xp25_ASAP7_75t_L g988 ( 
.A(n_983),
.B(n_868),
.C(n_858),
.D(n_857),
.Y(n_988)
);

AOI322xp5_ASAP7_75t_L g989 ( 
.A1(n_980),
.A2(n_891),
.A3(n_924),
.B1(n_911),
.B2(n_912),
.C1(n_916),
.C2(n_878),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_852),
.C(n_884),
.Y(n_990)
);

NAND3x1_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_866),
.C(n_852),
.Y(n_991)
);

OAI211xp5_ASAP7_75t_L g992 ( 
.A1(n_979),
.A2(n_830),
.B(n_856),
.C(n_885),
.Y(n_992)
);

AOI322xp5_ASAP7_75t_L g993 ( 
.A1(n_976),
.A2(n_924),
.A3(n_916),
.B1(n_878),
.B2(n_888),
.C1(n_883),
.C2(n_845),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_987),
.B(n_830),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_986),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_990),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_984),
.Y(n_998)
);

OAI22x1_ASAP7_75t_L g999 ( 
.A1(n_985),
.A2(n_989),
.B1(n_992),
.B2(n_988),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_993),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_987),
.A2(n_822),
.B1(n_838),
.B2(n_844),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_986),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_991),
.Y(n_1003)
);

AOI211xp5_ASAP7_75t_L g1004 ( 
.A1(n_998),
.A2(n_856),
.B(n_845),
.C(n_849),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_995),
.Y(n_1005)
);

NAND4xp25_ASAP7_75t_L g1006 ( 
.A(n_1000),
.B(n_996),
.C(n_1003),
.D(n_997),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_1002),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_L g1008 ( 
.A(n_994),
.B(n_893),
.C(n_849),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_1001),
.B(n_845),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1001),
.B(n_865),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_996),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_1006),
.B(n_865),
.Y(n_1013)
);

XNOR2x1_ASAP7_75t_L g1014 ( 
.A(n_1010),
.B(n_844),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1007),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_1012),
.B(n_888),
.Y(n_1016)
);

AO22x2_ASAP7_75t_L g1017 ( 
.A1(n_1015),
.A2(n_1008),
.B1(n_1005),
.B2(n_1011),
.Y(n_1017)
);

XOR2xp5_ASAP7_75t_L g1018 ( 
.A(n_1014),
.B(n_1004),
.Y(n_1018)
);

XOR2xp5_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_1009),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_1016),
.A2(n_856),
.B1(n_844),
.B2(n_850),
.Y(n_1020)
);

AOI221xp5_ASAP7_75t_SL g1021 ( 
.A1(n_1019),
.A2(n_850),
.B1(n_849),
.B2(n_877),
.C(n_886),
.Y(n_1021)
);

XNOR2xp5_ASAP7_75t_L g1022 ( 
.A(n_1018),
.B(n_844),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1022),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1021),
.A2(n_1017),
.B1(n_1020),
.B2(n_844),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

AOI211xp5_ASAP7_75t_L g1026 ( 
.A1(n_1024),
.A2(n_850),
.B(n_889),
.C(n_879),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1025),
.B(n_822),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1026),
.A2(n_822),
.B(n_844),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_1027),
.A2(n_828),
.B(n_827),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

AOI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_1030),
.A2(n_889),
.B1(n_869),
.B2(n_875),
.C(n_863),
.Y(n_1031)
);

OAI221xp5_ASAP7_75t_R g1032 ( 
.A1(n_1031),
.A2(n_1029),
.B1(n_886),
.B2(n_877),
.C(n_883),
.Y(n_1032)
);

AOI211xp5_ASAP7_75t_L g1033 ( 
.A1(n_1032),
.A2(n_881),
.B(n_863),
.C(n_879),
.Y(n_1033)
);


endmodule