module fake_jpeg_2118_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_77),
.Y(n_86)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_1),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_81),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_1),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_63),
.B1(n_55),
.B2(n_70),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_95),
.B1(n_64),
.B2(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_74),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_72),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_78),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_55),
.B1(n_70),
.B2(n_72),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_76),
.B1(n_64),
.B2(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_63),
.B1(n_53),
.B2(n_68),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_99),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_109),
.B1(n_73),
.B2(n_60),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_59),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_104),
.B1(n_97),
.B2(n_110),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_127),
.B1(n_4),
.B2(n_5),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_85),
.B(n_83),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_134),
.B(n_73),
.C(n_60),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_83),
.C(n_93),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_28),
.C(n_47),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_51),
.B1(n_61),
.B2(n_58),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_52),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_73),
.B(n_60),
.C(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_107),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_144),
.B(n_149),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_2),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_3),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_151),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_52),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.C(n_147),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_27),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_24),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_150),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_10),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_10),
.B(n_13),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_154),
.B(n_125),
.Y(n_160)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_13),
.CON(n_154),
.SN(n_154)
);

CKINVDCx12_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_34),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_32),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_132),
.B(n_128),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_166),
.B(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_169),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_49),
.B(n_33),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_46),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_178),
.C(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_16),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_35),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_167),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_175),
.B1(n_179),
.B2(n_153),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_184),
.C(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_148),
.C(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_172),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_166),
.B(n_163),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_168),
.C(n_163),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_160),
.B(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_144),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_193),
.B(n_29),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_170),
.C(n_37),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_187),
.C(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_181),
.C(n_182),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_39),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_199),
.B1(n_194),
.B2(n_19),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_205),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.C(n_208),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_207),
.A2(n_21),
.B(n_43),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_40),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_41),
.A3(n_44),
.B1(n_19),
.B2(n_20),
.C1(n_17),
.C2(n_18),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_18),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_20),
.Y(n_215)
);


endmodule