module real_aes_3046_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_1037, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_1038, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_1037;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_1038;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_571;
wire n_1034;
wire n_694;
wire n_491;
wire n_923;
wire n_549;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_973;
wire n_960;
wire n_455;
wire n_671;
wire n_725;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_936;
wire n_610;
wire n_581;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_649;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_691;
wire n_765;
wire n_481;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_831;
wire n_487;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_0), .A2(n_366), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_1), .A2(n_81), .B1(n_464), .B2(n_468), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_2), .A2(n_272), .B1(n_708), .B2(n_884), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_3), .A2(n_103), .B1(n_429), .B2(n_433), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_4), .A2(n_369), .B1(n_429), .B2(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_5), .A2(n_176), .B1(n_703), .B2(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_6), .A2(n_275), .B1(n_571), .B2(n_574), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_7), .A2(n_344), .B1(n_454), .B2(n_510), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_8), .A2(n_37), .B1(n_446), .B2(n_760), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_9), .A2(n_27), .B1(n_424), .B2(n_552), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_10), .A2(n_345), .B1(n_450), .B2(n_453), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_11), .A2(n_85), .B1(n_913), .B2(n_914), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_12), .A2(n_67), .B1(n_504), .B2(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_13), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_14), .A2(n_378), .B1(n_491), .B2(n_625), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_15), .A2(n_211), .B1(n_416), .B2(n_423), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_16), .A2(n_150), .B1(n_444), .B2(n_542), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_17), .A2(n_184), .B1(n_453), .B2(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_18), .A2(n_124), .B1(n_499), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_19), .A2(n_238), .B1(n_495), .B2(n_496), .Y(n_584) );
AO222x2_ASAP7_75t_L g580 ( .A1(n_20), .A2(n_201), .B1(n_253), .B2(n_488), .C1(n_491), .C2(n_492), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_21), .A2(n_155), .B1(n_440), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_22), .A2(n_23), .B1(n_565), .B2(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_24), .A2(n_363), .B1(n_507), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_25), .A2(n_127), .B1(n_506), .B2(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_26), .A2(n_186), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_28), .A2(n_35), .B1(n_689), .B2(n_691), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_29), .A2(n_245), .B1(n_571), .B2(n_572), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_30), .A2(n_178), .B1(n_535), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_31), .A2(n_126), .B1(n_528), .B2(n_886), .Y(n_885) );
AO22x1_ASAP7_75t_L g685 ( .A1(n_32), .A2(n_233), .B1(n_686), .B2(n_687), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_33), .A2(n_128), .B1(n_527), .B2(n_528), .Y(n_526) );
INVx1_ASAP7_75t_SL g404 ( .A(n_34), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g986 ( .A(n_34), .B(n_43), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_36), .A2(n_227), .B1(n_706), .B2(n_917), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_38), .A2(n_329), .B1(n_765), .B2(n_814), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_39), .A2(n_194), .B1(n_498), .B2(n_499), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_40), .A2(n_78), .B1(n_495), .B2(n_496), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_41), .B(n_538), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_42), .B(n_488), .Y(n_562) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_43), .A2(n_352), .B1(n_403), .B2(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_44), .B(n_488), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_45), .A2(n_308), .B1(n_819), .B2(n_881), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_46), .A2(n_84), .B1(n_780), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_47), .A2(n_361), .B1(n_643), .B2(n_687), .Y(n_1007) );
INVx1_ASAP7_75t_L g405 ( .A(n_48), .Y(n_405) );
AO22x1_ASAP7_75t_L g1014 ( .A1(n_49), .A2(n_165), .B1(n_699), .B2(n_778), .Y(n_1014) );
XNOR2xp5_ASAP7_75t_L g931 ( .A(n_50), .B(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_51), .A2(n_95), .B1(n_514), .B2(n_576), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_52), .A2(n_331), .B1(n_640), .B2(n_694), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_53), .A2(n_310), .B1(n_706), .B2(n_917), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_54), .A2(n_188), .B1(n_468), .B2(n_851), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_55), .A2(n_360), .B1(n_824), .B2(n_900), .Y(n_967) );
AO22x1_ASAP7_75t_L g688 ( .A1(n_56), .A2(n_375), .B1(n_689), .B2(n_691), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_57), .A2(n_893), .B1(n_906), .B2(n_907), .Y(n_892) );
INVx1_ASAP7_75t_L g906 ( .A(n_57), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_58), .A2(n_236), .B1(n_504), .B2(n_569), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_59), .A2(n_174), .B1(n_495), .B2(n_623), .Y(n_622) );
AO22x2_ASAP7_75t_L g413 ( .A1(n_60), .A2(n_181), .B1(n_403), .B2(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_61), .A2(n_370), .B1(n_434), .B2(n_801), .Y(n_800) );
AO22x1_ASAP7_75t_L g816 ( .A1(n_62), .A2(n_288), .B1(n_817), .B2(n_819), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_63), .A2(n_349), .B1(n_460), .B2(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_64), .A2(n_246), .B1(n_780), .B2(n_881), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_65), .A2(n_134), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_66), .A2(n_154), .B1(n_849), .B2(n_973), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_68), .A2(n_219), .B1(n_450), .B2(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_69), .A2(n_145), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_70), .A2(n_333), .B1(n_491), .B2(n_492), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_71), .A2(n_217), .B1(n_430), .B2(n_548), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_72), .A2(n_392), .B1(n_393), .B2(n_480), .Y(n_391) );
INVx1_ASAP7_75t_L g480 ( .A(n_72), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_73), .A2(n_89), .B1(n_190), .B2(n_488), .C1(n_498), .C2(n_583), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_74), .A2(n_285), .B1(n_513), .B2(n_514), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_75), .A2(n_256), .B1(n_534), .B2(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_76), .A2(n_192), .B1(n_513), .B2(n_574), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_77), .A2(n_101), .B1(n_464), .B2(n_468), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_79), .A2(n_379), .B1(n_498), .B2(n_583), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_80), .A2(n_359), .B1(n_498), .B2(n_583), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_82), .A2(n_1018), .B1(n_1019), .B2(n_1032), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g1018 ( .A(n_82), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_83), .A2(n_229), .B1(n_857), .B2(n_858), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_86), .B(n_397), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_87), .A2(n_137), .B1(n_503), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_88), .A2(n_199), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_90), .A2(n_116), .B1(n_504), .B2(n_569), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_91), .A2(n_205), .B1(n_514), .B2(n_576), .Y(n_575) );
OA22x2_ASAP7_75t_L g616 ( .A1(n_92), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_92), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_93), .A2(n_99), .B1(n_574), .B2(n_576), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_94), .A2(n_299), .B1(n_513), .B2(n_574), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_96), .A2(n_297), .B1(n_429), .B2(n_433), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_97), .A2(n_132), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_98), .A2(n_355), .B1(n_504), .B2(n_569), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_100), .A2(n_315), .B1(n_823), .B2(n_824), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_102), .A2(n_225), .B1(n_513), .B2(n_514), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_104), .A2(n_241), .B1(n_703), .B2(n_826), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_105), .A2(n_193), .B1(n_552), .B2(n_814), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_106), .A2(n_374), .B1(n_513), .B2(n_514), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_107), .A2(n_258), .B1(n_643), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_108), .A2(n_339), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_109), .A2(n_257), .B1(n_705), .B2(n_727), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_110), .A2(n_141), .B1(n_416), .B2(n_554), .Y(n_854) );
XNOR2xp5_ASAP7_75t_L g577 ( .A(n_111), .B(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_112), .A2(n_356), .B1(n_479), .B2(n_513), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_113), .A2(n_209), .B1(n_491), .B2(n_492), .Y(n_668) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_114), .A2(n_290), .B1(n_403), .B2(n_411), .Y(n_410) );
AOI222xp33_ASAP7_75t_SL g902 ( .A1(n_115), .A2(n_276), .B1(n_348), .B2(n_543), .C1(n_606), .C2(n_834), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_117), .A2(n_226), .B1(n_454), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_118), .A2(n_142), .B1(n_691), .B2(n_888), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g936 ( .A(n_119), .Y(n_936) );
XOR2x2_ASAP7_75t_L g792 ( .A(n_120), .B(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_121), .A2(n_291), .B1(n_730), .B2(n_734), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_122), .A2(n_372), .B1(n_729), .B2(n_730), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_123), .A2(n_332), .B1(n_530), .B2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_125), .A2(n_138), .B1(n_761), .B2(n_834), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_129), .A2(n_166), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_130), .A2(n_202), .B1(n_464), .B2(n_468), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_131), .A2(n_204), .B1(n_641), .B2(n_863), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_133), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_135), .A2(n_278), .B1(n_506), .B2(n_652), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_136), .A2(n_170), .B1(n_496), .B2(n_552), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_139), .A2(n_175), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_140), .A2(n_309), .B1(n_572), .B2(n_592), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_143), .A2(n_235), .B1(n_765), .B2(n_814), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_144), .A2(n_342), .B1(n_504), .B2(n_569), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_146), .A2(n_265), .B1(n_440), .B2(n_444), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_147), .A2(n_168), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g887 ( .A1(n_148), .A2(n_172), .B1(n_221), .B2(n_397), .C1(n_691), .C2(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_149), .A2(n_305), .B1(n_572), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_151), .A2(n_314), .B1(n_641), .B2(n_1029), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_152), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_153), .A2(n_210), .B1(n_886), .B2(n_1011), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_156), .A2(n_343), .B1(n_504), .B2(n_569), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_157), .A2(n_270), .B1(n_491), .B2(n_625), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_158), .B(n_637), .Y(n_636) );
AO21x2_ASAP7_75t_L g756 ( .A1(n_159), .A2(n_757), .B(n_781), .Y(n_756) );
INVx1_ASAP7_75t_L g783 ( .A(n_159), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_160), .A2(n_248), .B1(n_534), .B2(n_535), .Y(n_533) );
AO22x2_ASAP7_75t_L g742 ( .A1(n_161), .A2(n_743), .B1(n_754), .B2(n_755), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_161), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_162), .A2(n_325), .B1(n_464), .B2(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_163), .B(n_831), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_164), .A2(n_239), .B1(n_479), .B2(n_655), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_167), .A2(n_182), .B1(n_464), .B2(n_468), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_169), .A2(n_371), .B1(n_702), .B2(n_828), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_171), .A2(n_346), .B1(n_550), .B2(n_554), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_173), .A2(n_307), .B1(n_491), .B2(n_492), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_177), .A2(n_279), .B1(n_565), .B2(n_583), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_179), .A2(n_196), .B1(n_417), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_180), .A2(n_282), .B1(n_450), .B2(n_775), .Y(n_904) );
INVx1_ASAP7_75t_L g985 ( .A(n_181), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_183), .A2(n_286), .B1(n_423), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_185), .A2(n_334), .B1(n_530), .B2(n_532), .Y(n_529) );
AO222x2_ASAP7_75t_SL g759 ( .A1(n_187), .A2(n_283), .B1(n_341), .B2(n_606), .C1(n_760), .C2(n_761), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_189), .A2(n_302), .B1(n_571), .B2(n_572), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_191), .A2(n_380), .B1(n_513), .B2(n_514), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_195), .A2(n_254), .B1(n_506), .B2(n_514), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_197), .A2(n_249), .B1(n_495), .B2(n_496), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_198), .A2(n_323), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_200), .A2(n_295), .B1(n_886), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_203), .A2(n_287), .B1(n_545), .B2(n_547), .Y(n_964) );
XNOR2x2_ASAP7_75t_L g682 ( .A(n_206), .B(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_207), .A2(n_289), .B1(n_511), .B2(n_826), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_208), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_212), .B(n_691), .Y(n_937) );
NAND2xp5_ASAP7_75t_SL g965 ( .A(n_213), .B(n_538), .Y(n_965) );
AOI222xp33_ASAP7_75t_L g997 ( .A1(n_214), .A2(n_998), .B1(n_1015), .B2(n_1017), .C1(n_1033), .C2(n_1034), .Y(n_997) );
INVx1_ASAP7_75t_L g1001 ( .A(n_214), .Y(n_1001) );
XNOR2x1_ASAP7_75t_L g909 ( .A(n_215), .B(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g995 ( .A(n_216), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_218), .A2(n_311), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_220), .A2(n_301), .B1(n_761), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_222), .A2(n_381), .B1(n_510), .B2(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_223), .A2(n_873), .B1(n_889), .B2(n_890), .Y(n_872) );
INVx1_ASAP7_75t_L g890 ( .A(n_223), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_224), .B(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_228), .A2(n_337), .B1(n_444), .B2(n_863), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_230), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_231), .A2(n_243), .B1(n_545), .B2(n_547), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_232), .A2(n_336), .B1(n_504), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_234), .A2(n_340), .B1(n_652), .B2(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_237), .B(n_696), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_240), .A2(n_293), .B1(n_640), .B2(n_641), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_242), .A2(n_318), .B1(n_547), .B2(n_925), .Y(n_924) );
XNOR2x1_ASAP7_75t_L g559 ( .A(n_244), .B(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_247), .A2(n_317), .B1(n_554), .B2(n_643), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g945 ( .A(n_250), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_251), .A2(n_319), .B1(n_574), .B2(n_576), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_252), .A2(n_373), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_255), .A2(n_300), .B1(n_846), .B2(n_847), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_259), .Y(n_770) );
XOR2x2_ASAP7_75t_L g959 ( .A(n_260), .B(n_960), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_261), .A2(n_376), .B1(n_430), .B2(n_548), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_262), .A2(n_367), .B1(n_651), .B2(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_263), .A2(n_365), .B1(n_775), .B2(n_849), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g935 ( .A(n_264), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_266), .A2(n_335), .B1(n_457), .B2(n_460), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g948 ( .A1(n_267), .A2(n_354), .B1(n_528), .B2(n_884), .Y(n_948) );
XNOR2x1_ASAP7_75t_L g633 ( .A(n_268), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g515 ( .A(n_269), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_271), .A2(n_277), .B1(n_513), .B2(n_514), .Y(n_795) );
INVx1_ASAP7_75t_SL g996 ( .A(n_273), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_274), .A2(n_296), .B1(n_473), .B2(n_477), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_280), .A2(n_322), .B1(n_572), .B2(n_592), .Y(n_676) );
OA22x2_ASAP7_75t_L g594 ( .A1(n_281), .A2(n_595), .B1(n_596), .B2(n_610), .Y(n_594) );
INVx1_ASAP7_75t_L g610 ( .A(n_281), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_284), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_290), .B(n_984), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_292), .A2(n_347), .B1(n_686), .B2(n_923), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_294), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_298), .B(n_397), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_303), .A2(n_321), .B1(n_545), .B2(n_547), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_304), .A2(n_328), .B1(n_457), .B2(n_572), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_306), .A2(n_338), .B1(n_546), .B2(n_691), .Y(n_719) );
INVx3_ASAP7_75t_L g403 ( .A(n_312), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_313), .A2(n_327), .B1(n_534), .B2(n_778), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_316), .Y(n_773) );
OA22x2_ASAP7_75t_L g520 ( .A1(n_320), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_320), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_324), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_326), .B(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_330), .B(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_350), .A2(n_357), .B1(n_495), .B2(n_623), .Y(n_671) );
INVx1_ASAP7_75t_L g680 ( .A(n_351), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_353), .B(n_696), .Y(n_805) );
INVx1_ASAP7_75t_L g980 ( .A(n_358), .Y(n_980) );
NAND2xp5_ASAP7_75t_SL g994 ( .A(n_358), .B(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g981 ( .A(n_362), .Y(n_981) );
AND2x2_ASAP7_75t_R g1033 ( .A(n_362), .B(n_980), .Y(n_1033) );
INVx1_ASAP7_75t_L g815 ( .A(n_364), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_364), .A2(n_809), .B1(n_836), .B2(n_1037), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_364), .A2(n_821), .B1(n_829), .B2(n_1038), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_364), .B(n_816), .Y(n_838) );
INVxp67_ASAP7_75t_L g993 ( .A(n_368), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_377), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_975), .B(n_987), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_658), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI21xp33_ASAP7_75t_SL g975 ( .A1(n_385), .A2(n_976), .B(n_977), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_631), .B1(n_656), .B2(n_657), .Y(n_385) );
XOR2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_517), .Y(n_386) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_387), .B(n_517), .Y(n_656) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22x1_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_481), .B2(n_516), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_448), .Y(n_393) );
NAND4xp25_ASAP7_75t_SL g394 ( .A(n_395), .B(n_415), .C(n_428), .D(n_439), .Y(n_394) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx3_ASAP7_75t_SL g540 ( .A(n_398), .Y(n_540) );
INVx3_ASAP7_75t_L g606 ( .A(n_398), .Y(n_606) );
INVx4_ASAP7_75t_SL g637 ( .A(n_398), .Y(n_637) );
INVx4_ASAP7_75t_SL g696 ( .A(n_398), .Y(n_696) );
BUFx2_ASAP7_75t_L g832 ( .A(n_398), .Y(n_832) );
INVx6_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_408), .Y(n_399) );
AND2x4_ASAP7_75t_L g425 ( .A(n_400), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g446 ( .A(n_400), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g488 ( .A(n_400), .B(n_408), .Y(n_488) );
AND2x2_ASAP7_75t_L g496 ( .A(n_400), .B(n_426), .Y(n_496) );
AND2x2_ASAP7_75t_L g499 ( .A(n_400), .B(n_447), .Y(n_499) );
AND2x2_ASAP7_75t_L g583 ( .A(n_400), .B(n_447), .Y(n_583) );
AND2x2_ASAP7_75t_L g623 ( .A(n_400), .B(n_426), .Y(n_623) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_406), .Y(n_400) );
AND2x2_ASAP7_75t_L g421 ( .A(n_401), .B(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
INVx2_ASAP7_75t_L g443 ( .A(n_401), .Y(n_443) );
OAI22x1_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_403), .Y(n_407) );
INVx2_ASAP7_75t_L g411 ( .A(n_403), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_403), .Y(n_414) );
INVx2_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
AND2x2_ASAP7_75t_L g442 ( .A(n_406), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g471 ( .A(n_406), .Y(n_471) );
AND2x4_ASAP7_75t_L g452 ( .A(n_408), .B(n_421), .Y(n_452) );
AND2x4_ASAP7_75t_L g459 ( .A(n_408), .B(n_455), .Y(n_459) );
AND2x2_ASAP7_75t_L g476 ( .A(n_408), .B(n_442), .Y(n_476) );
AND2x6_ASAP7_75t_L g513 ( .A(n_408), .B(n_442), .Y(n_513) );
AND2x2_ASAP7_75t_L g571 ( .A(n_408), .B(n_421), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_408), .B(n_455), .Y(n_576) );
AND2x2_ASAP7_75t_L g592 ( .A(n_408), .B(n_421), .Y(n_592) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g420 ( .A(n_410), .Y(n_420) );
AND2x4_ASAP7_75t_L g432 ( .A(n_410), .B(n_412), .Y(n_432) );
AND2x2_ASAP7_75t_L g437 ( .A(n_410), .B(n_413), .Y(n_437) );
INVxp67_ASAP7_75t_L g447 ( .A(n_412), .Y(n_447) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g419 ( .A(n_413), .B(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g553 ( .A(n_418), .Y(n_553) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_418), .Y(n_643) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
AND2x4_ASAP7_75t_L g462 ( .A(n_419), .B(n_455), .Y(n_462) );
AND2x2_ASAP7_75t_L g467 ( .A(n_419), .B(n_442), .Y(n_467) );
AND2x4_ASAP7_75t_L g495 ( .A(n_419), .B(n_421), .Y(n_495) );
AND2x6_ASAP7_75t_L g514 ( .A(n_419), .B(n_455), .Y(n_514) );
AND2x2_ASAP7_75t_L g569 ( .A(n_419), .B(n_442), .Y(n_569) );
AND2x2_ASAP7_75t_SL g588 ( .A(n_419), .B(n_442), .Y(n_588) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_420), .Y(n_427) );
AND2x2_ASAP7_75t_L g431 ( .A(n_421), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g491 ( .A(n_421), .B(n_432), .Y(n_491) );
AND2x4_ASAP7_75t_L g455 ( .A(n_422), .B(n_443), .Y(n_455) );
BUFx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g556 ( .A(n_425), .Y(n_556) );
INVx1_ASAP7_75t_L g645 ( .A(n_425), .Y(n_645) );
BUFx3_ASAP7_75t_L g723 ( .A(n_425), .Y(n_723) );
BUFx4f_ASAP7_75t_L g923 ( .A(n_425), .Y(n_923) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g546 ( .A(n_431), .Y(n_546) );
INVx2_ASAP7_75t_L g690 ( .A(n_431), .Y(n_690) );
BUFx5_ASAP7_75t_L g888 ( .A(n_431), .Y(n_888) );
AND2x4_ASAP7_75t_L g441 ( .A(n_432), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g479 ( .A(n_432), .B(n_455), .Y(n_479) );
AND2x2_ASAP7_75t_L g498 ( .A(n_432), .B(n_442), .Y(n_498) );
AND2x2_ASAP7_75t_L g565 ( .A(n_432), .B(n_442), .Y(n_565) );
AND2x2_ASAP7_75t_L g574 ( .A(n_432), .B(n_455), .Y(n_574) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g548 ( .A(n_435), .Y(n_548) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx12f_ASAP7_75t_L g691 ( .A(n_436), .Y(n_691) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x4_ASAP7_75t_L g454 ( .A(n_437), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g470 ( .A(n_437), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_437), .B(n_438), .Y(n_492) );
AND2x4_ASAP7_75t_L g504 ( .A(n_437), .B(n_471), .Y(n_504) );
AND2x4_ASAP7_75t_L g572 ( .A(n_437), .B(n_455), .Y(n_572) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_437), .B(n_438), .Y(n_625) );
BUFx4f_ASAP7_75t_SL g542 ( .A(n_440), .Y(n_542) );
BUFx2_ASAP7_75t_L g760 ( .A(n_440), .Y(n_760) );
BUFx2_ASAP7_75t_L g834 ( .A(n_440), .Y(n_834) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g640 ( .A(n_441), .Y(n_640) );
BUFx3_ASAP7_75t_L g863 ( .A(n_441), .Y(n_863) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_441), .Y(n_1029) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g543 ( .A(n_445), .Y(n_543) );
INVx2_ASAP7_75t_SL g641 ( .A(n_445), .Y(n_641) );
INVx2_ASAP7_75t_L g694 ( .A(n_445), .Y(n_694) );
INVx2_ASAP7_75t_L g761 ( .A(n_445), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_445), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_942) );
INVx6_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_456), .C(n_463), .D(n_472), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g527 ( .A(n_451), .Y(n_527) );
INVx3_ASAP7_75t_L g826 ( .A(n_451), .Y(n_826) );
INVx1_ASAP7_75t_SL g849 ( .A(n_451), .Y(n_849) );
INVx2_ASAP7_75t_L g884 ( .A(n_451), .Y(n_884) );
INVx6_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
BUFx3_ASAP7_75t_L g649 ( .A(n_452), .Y(n_649) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
BUFx2_ASAP7_75t_SL g528 ( .A(n_454), .Y(n_528) );
INVx2_ASAP7_75t_L g709 ( .A(n_454), .Y(n_709) );
BUFx2_ASAP7_75t_SL g973 ( .A(n_454), .Y(n_973) );
INVx2_ASAP7_75t_L g531 ( .A(n_457), .Y(n_531) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_457), .Y(n_913) );
INVx4_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_SL g506 ( .A(n_458), .Y(n_506) );
INVx3_ASAP7_75t_L g655 ( .A(n_458), .Y(n_655) );
INVx2_ASAP7_75t_SL g702 ( .A(n_458), .Y(n_702) );
INVx2_ASAP7_75t_L g734 ( .A(n_458), .Y(n_734) );
INVx2_ASAP7_75t_SL g886 ( .A(n_458), .Y(n_886) );
INVx8_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g535 ( .A(n_461), .Y(n_535) );
INVx2_ASAP7_75t_L g700 ( .A(n_461), .Y(n_700) );
INVx2_ASAP7_75t_L g730 ( .A(n_461), .Y(n_730) );
INVx2_ASAP7_75t_SL g778 ( .A(n_461), .Y(n_778) );
INVx2_ASAP7_75t_L g824 ( .A(n_461), .Y(n_824) );
INVx2_ASAP7_75t_SL g847 ( .A(n_461), .Y(n_847) );
INVx1_ASAP7_75t_SL g952 ( .A(n_461), .Y(n_952) );
INVx8_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g705 ( .A(n_466), .Y(n_705) );
INVx2_ASAP7_75t_L g818 ( .A(n_466), .Y(n_818) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g503 ( .A(n_467), .Y(n_503) );
BUFx6f_ASAP7_75t_L g881 ( .A(n_467), .Y(n_881) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g706 ( .A(n_469), .Y(n_706) );
INVx2_ASAP7_75t_L g727 ( .A(n_469), .Y(n_727) );
INVx2_ASAP7_75t_L g780 ( .A(n_469), .Y(n_780) );
INVx5_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g602 ( .A(n_470), .Y(n_602) );
BUFx3_ASAP7_75t_L g819 ( .A(n_470), .Y(n_819) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g534 ( .A(n_475), .Y(n_534) );
INVx3_ASAP7_75t_L g651 ( .A(n_475), .Y(n_651) );
INVx2_ASAP7_75t_L g699 ( .A(n_475), .Y(n_699) );
INVx2_ASAP7_75t_SL g879 ( .A(n_475), .Y(n_879) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g729 ( .A(n_476), .Y(n_729) );
BUFx2_ASAP7_75t_L g823 ( .A(n_476), .Y(n_823) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g955 ( .A(n_478), .Y(n_955) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_479), .Y(n_507) );
INVx2_ASAP7_75t_L g653 ( .A(n_479), .Y(n_653) );
BUFx3_ASAP7_75t_L g703 ( .A(n_479), .Y(n_703) );
INVx1_ASAP7_75t_SL g516 ( .A(n_481), .Y(n_516) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
XOR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_515), .Y(n_483) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_500), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_489), .B(n_490), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_508), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
BUFx2_ASAP7_75t_L g851 ( .A(n_503), .Y(n_851) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_507), .Y(n_532) );
INVx2_ASAP7_75t_L g971 ( .A(n_507), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_512), .Y(n_508) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_511), .Y(n_775) );
XOR2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_614), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B1(n_557), .B2(n_613), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .C(n_529), .D(n_533), .Y(n_524) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND4xp25_ASAP7_75t_SL g536 ( .A(n_537), .B(n_541), .C(n_544), .D(n_549), .Y(n_536) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI21xp33_ASAP7_75t_SL g717 ( .A1(n_539), .A2(n_718), .B(n_719), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_539), .A2(n_926), .B1(n_935), .B2(n_936), .C(n_937), .Y(n_934) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g944 ( .A(n_542), .Y(n_944) );
BUFx6f_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g926 ( .A(n_546), .Y(n_926) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g686 ( .A(n_553), .Y(n_686) );
INVx1_ASAP7_75t_L g766 ( .A(n_553), .Y(n_766) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_555), .A2(n_939), .B1(n_940), .B2(n_941), .Y(n_938) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g687 ( .A(n_556), .Y(n_687) );
INVx1_ASAP7_75t_L g613 ( .A(n_557), .Y(n_613) );
OA22x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_594), .B1(n_611), .B2(n_612), .Y(n_557) );
INVx1_ASAP7_75t_L g612 ( .A(n_558), .Y(n_612) );
XOR2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_577), .Y(n_558) );
INVx1_ASAP7_75t_L g841 ( .A(n_559), .Y(n_841) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_559), .Y(n_866) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .Y(n_560) );
NAND4xp25_ASAP7_75t_SL g561 ( .A(n_562), .B(n_563), .C(n_564), .D(n_566), .Y(n_561) );
NAND4xp25_ASAP7_75t_SL g567 ( .A(n_568), .B(n_570), .C(n_573), .D(n_575), .Y(n_567) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_585), .Y(n_578) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_590), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g611 ( .A(n_594), .Y(n_611) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_597), .B(n_604), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .C(n_603), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .C(n_608), .D(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_626), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .C(n_624), .Y(n_620) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .C(n_629), .D(n_630), .Y(n_626) );
INVx2_ASAP7_75t_L g657 ( .A(n_631), .Y(n_657) );
BUFx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_646), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .C(n_639), .D(n_642), .Y(n_635) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .C(n_650), .D(n_654), .Y(n_646) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g828 ( .A(n_653), .Y(n_828) );
INVx1_ASAP7_75t_L g914 ( .A(n_653), .Y(n_914) );
INVx1_ASAP7_75t_L g976 ( .A(n_658), .Y(n_976) );
XNOR2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_786), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_739), .B1(n_784), .B2(n_785), .Y(n_660) );
INVx1_ASAP7_75t_SL g784 ( .A(n_661), .Y(n_784) );
AOI22x1_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_711), .B1(n_736), .B2(n_737), .Y(n_661) );
BUFx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g736 ( .A(n_663), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_681), .B1(n_682), .B2(n_710), .Y(n_663) );
INVx3_ASAP7_75t_SL g710 ( .A(n_664), .Y(n_710) );
XOR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_680), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_673), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_697), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .C(n_692), .Y(n_684) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g801 ( .A(n_690), .Y(n_801) );
INVx2_ASAP7_75t_L g857 ( .A(n_690), .Y(n_857) );
BUFx3_ASAP7_75t_L g811 ( .A(n_691), .Y(n_811) );
INVx2_ASAP7_75t_L g859 ( .A(n_691), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_693), .B(n_695), .Y(n_692) );
AND4x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .C(n_704), .D(n_707), .Y(n_697) );
BUFx2_ASAP7_75t_L g772 ( .A(n_703), .Y(n_772) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_709), .Y(n_1011) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g738 ( .A(n_714), .Y(n_738) );
XNOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_735), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_724), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
BUFx6f_ASAP7_75t_SL g814 ( .A(n_723), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_731), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
BUFx3_ASAP7_75t_L g846 ( .A(n_729), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g769 ( .A(n_734), .Y(n_769) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVxp33_ASAP7_75t_L g785 ( .A(n_740), .Y(n_785) );
XNOR2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_756), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g755 ( .A(n_743), .Y(n_755) );
NOR2xp67_ASAP7_75t_L g743 ( .A(n_744), .B(n_749), .Y(n_743) );
NAND4xp25_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .C(n_747), .D(n_748), .Y(n_744) );
NAND4xp25_ASAP7_75t_SL g749 ( .A(n_750), .B(n_751), .C(n_752), .D(n_753), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_767), .C(n_776), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .Y(n_758) );
NOR4xp25_ASAP7_75t_L g781 ( .A(n_759), .B(n_762), .C(n_768), .D(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g940 ( .A(n_765), .Y(n_940) );
BUFx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
OAI221xp5_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_770), .B1(n_771), .B2(n_773), .C(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g782 ( .A(n_776), .B(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_927), .B2(n_974), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
XOR2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_868), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_839), .B2(n_867), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
XNOR2x1_ASAP7_75t_L g791 ( .A(n_792), .B(n_806), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_792), .A2(n_931), .B1(n_956), .B2(n_957), .Y(n_930) );
INVx2_ASAP7_75t_L g956 ( .A(n_792), .Y(n_956) );
NOR3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_799), .C(n_803), .Y(n_793) );
NAND4xp25_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .C(n_797), .D(n_798), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
NAND4xp75_ASAP7_75t_L g806 ( .A(n_807), .B(n_835), .C(n_837), .D(n_838), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_820), .Y(n_807) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .C(n_816), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g812 ( .A(n_813), .B(n_815), .Y(n_812) );
INVx1_ASAP7_75t_L g836 ( .A(n_813), .Y(n_836) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
BUFx6f_ASAP7_75t_L g917 ( .A(n_818), .Y(n_917) );
NOR2xp67_ASAP7_75t_L g820 ( .A(n_821), .B(n_829), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .C(n_827), .Y(n_821) );
INVx2_ASAP7_75t_L g901 ( .A(n_823), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
INVx2_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g867 ( .A(n_839), .Y(n_867) );
OAI21xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_842), .B(n_865), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_SL g865 ( .A(n_842), .B(n_866), .Y(n_865) );
XOR2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_864), .Y(n_842) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_844), .B(n_853), .Y(n_843) );
NAND4xp25_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .C(n_850), .D(n_852), .Y(n_844) );
NAND4xp25_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .C(n_856), .D(n_860), .Y(n_853) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
XNOR2xp5_ASAP7_75t_L g868 ( .A(n_869), .B(n_891), .Y(n_868) );
INVx1_ASAP7_75t_SL g869 ( .A(n_870), .Y(n_869) );
BUFx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g889 ( .A(n_873), .Y(n_889) );
NAND4xp75_ASAP7_75t_L g873 ( .A(n_874), .B(n_877), .C(n_882), .D(n_887), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_885), .Y(n_882) );
XNOR2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_908), .Y(n_891) );
INVx2_ASAP7_75t_L g907 ( .A(n_893), .Y(n_907) );
NAND4xp75_ASAP7_75t_L g893 ( .A(n_894), .B(n_897), .C(n_902), .D(n_903), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_895), .B(n_896), .Y(n_894) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
AND2x2_ASAP7_75t_SL g903 ( .A(n_904), .B(n_905), .Y(n_903) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
NOR2x1_ASAP7_75t_L g910 ( .A(n_911), .B(n_919), .Y(n_910) );
NAND4xp25_ASAP7_75t_L g911 ( .A(n_912), .B(n_915), .C(n_916), .D(n_918), .Y(n_911) );
NAND4xp25_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .C(n_922), .D(n_924), .Y(n_919) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_928), .Y(n_974) );
OA22x2_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_958), .B2(n_959), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g957 ( .A(n_931), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_946), .Y(n_932) );
NOR3xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_938), .C(n_942), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_950), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_953), .Y(n_950) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx4_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NOR2x1_ASAP7_75t_L g960 ( .A(n_961), .B(n_966), .Y(n_960) );
NAND4xp25_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .C(n_964), .D(n_965), .Y(n_961) );
NAND4xp25_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .C(n_969), .D(n_972), .Y(n_966) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx4_ASAP7_75t_R g977 ( .A(n_978), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_982), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_979), .B(n_983), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g991 ( .A(n_981), .Y(n_991) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_986), .Y(n_984) );
OAI21xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_996), .B(n_997), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_989), .Y(n_988) );
AND2x4_ASAP7_75t_SL g989 ( .A(n_990), .B(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_991), .B(n_992), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
XNOR2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .Y(n_1000) );
NAND2xp5_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1008), .Y(n_1002) );
AND4x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1005), .C(n_1006), .D(n_1007), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1014), .Y(n_1008) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1012), .C(n_1013), .Y(n_1009) );
CKINVDCx6p67_ASAP7_75t_R g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1019), .Y(n_1032) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
NOR2xp67_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1026), .Y(n_1020) );
NAND4xp25_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1023), .C(n_1024), .D(n_1025), .Y(n_1021) );
NAND4xp25_ASAP7_75t_SL g1026 ( .A(n_1027), .B(n_1028), .C(n_1030), .D(n_1031), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_1035), .Y(n_1034) );
endmodule