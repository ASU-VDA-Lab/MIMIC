module fake_jpeg_11665_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_80),
.Y(n_132)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_69),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_81),
.B(n_82),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_23),
.B(n_15),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_15),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_59),
.Y(n_152)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_90),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_13),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_95),
.B(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_40),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_99),
.Y(n_137)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_40),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_45),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_113),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_112),
.Y(n_146)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_31),
.B(n_11),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_31),
.B(n_10),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_39),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_50),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_121),
.B1(n_30),
.B2(n_52),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_124),
.Y(n_155)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_61),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_141),
.A2(n_162),
.B1(n_21),
.B2(n_125),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_144),
.B(n_186),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_71),
.B(n_25),
.C(n_53),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_145),
.B(n_181),
.C(n_55),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_91),
.A2(n_30),
.B1(n_60),
.B2(n_58),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_149),
.A2(n_185),
.B1(n_192),
.B2(n_83),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_152),
.B(n_153),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_108),
.A2(n_57),
.B1(n_46),
.B2(n_21),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_156),
.A2(n_105),
.B1(n_102),
.B2(n_101),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_66),
.A2(n_41),
.B1(n_49),
.B2(n_56),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_157),
.A2(n_76),
.B1(n_73),
.B2(n_98),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_39),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_160),
.B(n_163),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_74),
.A2(n_30),
.B1(n_59),
.B2(n_29),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_34),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_179),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_79),
.A2(n_43),
.B(n_37),
.C(n_35),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_169),
.A2(n_55),
.B(n_38),
.C(n_112),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_68),
.B(n_34),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_172),
.B(n_176),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_67),
.A2(n_56),
.B1(n_49),
.B2(n_41),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_175),
.A2(n_193),
.B1(n_110),
.B2(n_103),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_68),
.B(n_43),
.Y(n_176)
);

AND2x4_ASAP7_75t_SL g179 ( 
.A(n_85),
.B(n_60),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_46),
.C(n_35),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_87),
.A2(n_60),
.B1(n_55),
.B2(n_38),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_75),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_28),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_187),
.B(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_194),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_104),
.A2(n_55),
.B1(n_38),
.B2(n_21),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_70),
.A2(n_52),
.B1(n_33),
.B2(n_29),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_100),
.B(n_33),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_64),
.B(n_51),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_198),
.B(n_209),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_93),
.B(n_51),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_94),
.B(n_47),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_210),
.B(n_217),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_132),
.B(n_47),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_211),
.B(n_221),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_212),
.Y(n_302)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_173),
.B(n_37),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_215),
.B(n_223),
.Y(n_288)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_216),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_243),
.B1(n_164),
.B2(n_189),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_222),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_146),
.Y(n_223)
);

OR2x4_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_72),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_224),
.A2(n_6),
.B(n_7),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_225),
.A2(n_231),
.B1(n_251),
.B2(n_254),
.Y(n_298)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_227),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_130),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_228),
.B(n_245),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_162),
.A2(n_63),
.B1(n_141),
.B2(n_143),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_229),
.Y(n_324)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_230),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_149),
.A2(n_89),
.B1(n_118),
.B2(n_117),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_236),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_133),
.Y(n_291)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_138),
.A2(n_38),
.B1(n_55),
.B2(n_167),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_240),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_0),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_252),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_156),
.A2(n_84),
.B1(n_114),
.B2(n_109),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_147),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_246),
.B(n_259),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_247),
.A2(n_148),
.B(n_190),
.Y(n_297)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_249),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_138),
.A2(n_124),
.B1(n_112),
.B2(n_90),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_250),
.A2(n_283),
.B1(n_154),
.B2(n_139),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_168),
.B(n_2),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_256),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_185),
.A2(n_124),
.B1(n_122),
.B2(n_116),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_257),
.A2(n_265),
.B1(n_269),
.B2(n_6),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_145),
.B(n_201),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_272),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_135),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_134),
.Y(n_260)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_142),
.Y(n_261)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_165),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_263),
.Y(n_316)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_192),
.A2(n_113),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

BUFx16f_ASAP7_75t_L g266 ( 
.A(n_134),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_266),
.B(n_268),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_275),
.Y(n_319)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_191),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_155),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_273),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_140),
.B(n_3),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_271),
.B(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_203),
.B(n_3),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_158),
.B(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_276),
.B(n_279),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_282),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_159),
.B(n_4),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_131),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_191),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_195),
.B1(n_171),
.B2(n_197),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_161),
.B(n_5),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_150),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_180),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_6),
.Y(n_333)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_285),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_221),
.A2(n_165),
.B(n_133),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_286),
.A2(n_261),
.B(n_263),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_223),
.A2(n_195),
.B1(n_197),
.B2(n_170),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_287),
.A2(n_296),
.B1(n_301),
.B2(n_332),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_267),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_293),
.A2(n_299),
.B1(n_338),
.B2(n_347),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_297),
.B(n_315),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_148),
.B1(n_170),
.B2(n_171),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_235),
.A2(n_164),
.B1(n_189),
.B2(n_183),
.Y(n_301)
);

AOI32xp33_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_154),
.A3(n_131),
.B1(n_180),
.B2(n_190),
.Y(n_312)
);

A2O1A1O1Ixp25_ASAP7_75t_L g376 ( 
.A1(n_312),
.A2(n_297),
.B(n_343),
.C(n_257),
.D(n_324),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g313 ( 
.A1(n_235),
.A2(n_139),
.A3(n_204),
.B1(n_207),
.B2(n_178),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_327),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_237),
.B(n_151),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_323),
.C(n_328),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_237),
.B(n_151),
.C(n_183),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_211),
.B(n_178),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_207),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_274),
.A2(n_242),
.B1(n_220),
.B2(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_215),
.B(n_6),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_345),
.C(n_245),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_210),
.B(n_7),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_342),
.B(n_228),
.Y(n_353)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_224),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_SL g388 ( 
.A1(n_344),
.A2(n_246),
.B(n_285),
.C(n_212),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_241),
.B(n_8),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_254),
.A2(n_8),
.B1(n_9),
.B2(n_225),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_220),
.A2(n_8),
.B1(n_276),
.B2(n_259),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_269),
.B1(n_231),
.B2(n_265),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_322),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_349),
.B(n_350),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_252),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_353),
.B(n_355),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_217),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_364),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_357),
.B(n_360),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_310),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_361),
.B(n_370),
.Y(n_417)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_318),
.Y(n_362)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_302),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_376),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_219),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_365),
.B(n_384),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_291),
.B(n_270),
.C(n_262),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_367),
.C(n_381),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_314),
.B(n_239),
.C(n_216),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_368),
.Y(n_426)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_308),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_325),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_371),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_288),
.B(n_219),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_372),
.B(n_380),
.Y(n_414)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_329),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_377),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_385),
.B1(n_390),
.B2(n_293),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_302),
.B(n_213),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_323),
.B(n_222),
.C(n_256),
.Y(n_381)
);

OAI32xp33_ASAP7_75t_L g382 ( 
.A1(n_290),
.A2(n_213),
.A3(n_248),
.B1(n_275),
.B2(n_264),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_382),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_289),
.B(n_233),
.C(n_214),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_396),
.C(n_320),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_319),
.B(n_253),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_332),
.A2(n_226),
.B1(n_236),
.B2(n_238),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_290),
.B(n_248),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_386),
.B(n_389),
.Y(n_432)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

AO21x2_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_344),
.B(n_346),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_304),
.B(n_328),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_324),
.A2(n_255),
.B1(n_249),
.B2(n_284),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_315),
.A2(n_279),
.B(n_272),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_393),
.B(n_286),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_234),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_392),
.B(n_397),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_212),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_304),
.B(n_230),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_337),
.Y(n_424)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_268),
.C(n_280),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_399),
.A2(n_401),
.B1(n_407),
.B2(n_413),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_359),
.A2(n_338),
.B1(n_298),
.B2(n_292),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_359),
.A2(n_378),
.B1(n_354),
.B2(n_298),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_379),
.A2(n_292),
.B1(n_287),
.B2(n_343),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_408),
.A2(n_440),
.B1(n_355),
.B2(n_351),
.Y(n_450)
);

AO22x2_ASAP7_75t_L g466 ( 
.A1(n_411),
.A2(n_421),
.B1(n_388),
.B2(n_309),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_357),
.A2(n_347),
.B1(n_335),
.B2(n_313),
.Y(n_413)
);

OAI22x1_ASAP7_75t_L g415 ( 
.A1(n_393),
.A2(n_327),
.B1(n_344),
.B2(n_321),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_415),
.A2(n_266),
.B(n_273),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_295),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_431),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_358),
.B(n_321),
.C(n_330),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_431),
.C(n_435),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_309),
.Y(n_457)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_352),
.A2(n_344),
.B1(n_346),
.B2(n_321),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_430),
.A2(n_437),
.B1(n_375),
.B2(n_363),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_365),
.B(n_337),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_379),
.A2(n_305),
.B1(n_303),
.B2(n_339),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_390),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_358),
.B(n_334),
.C(n_330),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_360),
.A2(n_244),
.B1(n_283),
.B2(n_305),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_366),
.B(n_334),
.C(n_294),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_383),
.C(n_396),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_352),
.B1(n_376),
.B2(n_384),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_387),
.Y(n_442)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_395),
.Y(n_444)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_410),
.Y(n_445)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_445),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_421),
.A2(n_393),
.B1(n_397),
.B2(n_351),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_446),
.A2(n_452),
.B1(n_441),
.B2(n_400),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_447),
.B(n_427),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_350),
.Y(n_449)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_449),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_450),
.A2(n_438),
.B1(n_430),
.B2(n_408),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_451),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_440),
.A2(n_381),
.B1(n_367),
.B2(n_389),
.Y(n_452)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_394),
.B1(n_374),
.B2(n_371),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_454),
.A2(n_467),
.B1(n_474),
.B2(n_451),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_434),
.B(n_386),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g485 ( 
.A(n_455),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g456 ( 
.A1(n_436),
.A2(n_382),
.A3(n_349),
.B1(n_353),
.B2(n_394),
.C1(n_385),
.C2(n_391),
.Y(n_456)
);

AOI21xp33_ASAP7_75t_L g491 ( 
.A1(n_456),
.A2(n_459),
.B(n_461),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_457),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_402),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_458),
.B(n_469),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_411),
.A2(n_388),
.B(n_398),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_404),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_462),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_438),
.A2(n_388),
.B(n_373),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_377),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_361),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_465),
.C(n_470),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_421),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_403),
.A2(n_388),
.B1(n_339),
.B2(n_244),
.Y(n_467)
);

AOI322xp5_ASAP7_75t_L g468 ( 
.A1(n_436),
.A2(n_331),
.A3(n_283),
.B1(n_294),
.B2(n_295),
.C1(n_311),
.C2(n_280),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_SL g487 ( 
.A(n_468),
.B(n_471),
.C(n_439),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_416),
.B(n_317),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_432),
.B(n_311),
.CI(n_317),
.CON(n_471),
.SN(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_232),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_475),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_331),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_473),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_403),
.A2(n_306),
.B1(n_277),
.B2(n_260),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_432),
.B(n_306),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_417),
.B(n_420),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_476),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_403),
.A2(n_266),
.B(n_273),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_477),
.A2(n_478),
.B(n_419),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_420),
.B(n_435),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_424),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_415),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_481),
.B(n_494),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_484),
.A2(n_498),
.B1(n_474),
.B2(n_477),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_487),
.B(n_513),
.Y(n_531)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_490),
.B(n_504),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_423),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_496),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_462),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_508),
.C(n_513),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_438),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_442),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_455),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_443),
.A2(n_454),
.B1(n_453),
.B2(n_467),
.Y(n_500)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_502),
.A2(n_506),
.B(n_512),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_447),
.B(n_421),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_450),
.A2(n_421),
.B1(n_400),
.B2(n_405),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_464),
.B(n_422),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_443),
.A2(n_422),
.B1(n_405),
.B2(n_425),
.Y(n_511)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_511),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_452),
.B(n_425),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_515),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_491),
.A2(n_459),
.B(n_461),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_516),
.A2(n_521),
.B(n_480),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_517),
.A2(n_519),
.B1(n_526),
.B2(n_535),
.Y(n_564)
);

OA22x2_ASAP7_75t_L g518 ( 
.A1(n_502),
.A2(n_466),
.B1(n_446),
.B2(n_478),
.Y(n_518)
);

A2O1A1Ixp33_ASAP7_75t_SL g554 ( 
.A1(n_518),
.A2(n_521),
.B(n_516),
.C(n_514),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_449),
.B1(n_460),
.B2(n_444),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_512),
.A2(n_466),
.B(n_475),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_466),
.Y(n_522)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_472),
.C(n_470),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_530),
.C(n_523),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_499),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_525),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_484),
.A2(n_471),
.B1(n_466),
.B2(n_465),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_471),
.B(n_448),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_528),
.A2(n_532),
.B(n_538),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_493),
.B(n_463),
.C(n_448),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_531),
.B(n_541),
.Y(n_547)
);

CKINVDCx14_ASAP7_75t_R g532 ( 
.A(n_499),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_498),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_488),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_507),
.A2(n_418),
.B1(n_429),
.B2(n_426),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_497),
.B(n_505),
.Y(n_536)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_536),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_483),
.A2(n_409),
.B(n_419),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_539),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_509),
.B(n_418),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_540),
.B(n_482),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_503),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_507),
.A2(n_409),
.B1(n_426),
.B2(n_428),
.Y(n_543)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_543),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_508),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_561),
.Y(n_585)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_546),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_520),
.A2(n_485),
.B1(n_482),
.B2(n_505),
.Y(n_550)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_550),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_520),
.A2(n_501),
.B1(n_486),
.B2(n_489),
.Y(n_551)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_551),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_533),
.A2(n_501),
.B1(n_489),
.B2(n_494),
.Y(n_552)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_553),
.B(n_565),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_560),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_495),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_558),
.B(n_559),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_496),
.Y(n_559)
);

XNOR2x1_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_504),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_527),
.A2(n_500),
.B1(n_487),
.B2(n_511),
.Y(n_562)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_562),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_492),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_538),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_540),
.B(n_480),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_566),
.A2(n_528),
.B(n_514),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_527),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_567),
.B(n_536),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_563),
.B(n_523),
.C(n_531),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_570),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_490),
.C(n_526),
.Y(n_570)
);

NOR2x1_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_542),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_548),
.B(n_566),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_564),
.A2(n_522),
.B1(n_542),
.B2(n_515),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_574),
.A2(n_551),
.B1(n_552),
.B2(n_548),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_529),
.C(n_534),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_576),
.B(n_577),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_547),
.B(n_519),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_578),
.A2(n_583),
.B(n_545),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_534),
.C(n_517),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_579),
.B(n_580),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_568),
.B(n_539),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_545),
.A2(n_532),
.B(n_525),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_556),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_586),
.B(n_549),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_590),
.B(n_592),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_564),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_593),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_559),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_575),
.B(n_562),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_595),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_579),
.B(n_557),
.C(n_554),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_596),
.B(n_604),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_597),
.A2(n_582),
.B1(n_588),
.B2(n_578),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_557),
.C(n_554),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_598),
.B(n_603),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_602),
.A2(n_605),
.B(n_535),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_589),
.A2(n_573),
.B1(n_587),
.B2(n_582),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_567),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_576),
.B(n_555),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_606),
.B(n_607),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_575),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_595),
.B(n_586),
.C(n_581),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_611),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_610),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_581),
.C(n_569),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_596),
.A2(n_574),
.B1(n_588),
.B2(n_555),
.Y(n_612)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_612),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_599),
.A2(n_572),
.B(n_570),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_613),
.B(n_614),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_600),
.B(n_554),
.C(n_585),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_620),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_594),
.B(n_543),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_602),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_622),
.A2(n_627),
.B(n_616),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_608),
.B(n_598),
.C(n_604),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_628),
.Y(n_632)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_611),
.B(n_604),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_617),
.B(n_597),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_619),
.B(n_592),
.C(n_605),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_630),
.B(n_616),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_625),
.A2(n_615),
.B1(n_609),
.B2(n_612),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_633),
.B(n_635),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_634),
.A2(n_637),
.B(n_518),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_623),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_636),
.B(n_638),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_630),
.A2(n_618),
.B(n_621),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_610),
.Y(n_638)
);

AOI321xp33_ASAP7_75t_L g639 ( 
.A1(n_632),
.A2(n_624),
.A3(n_622),
.B1(n_621),
.B2(n_629),
.C(n_626),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_639),
.A2(n_518),
.B1(n_561),
.B2(n_273),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_641),
.Y(n_644)
);

OAI321xp33_ASAP7_75t_L g645 ( 
.A1(n_643),
.A2(n_518),
.A3(n_640),
.B1(n_642),
.B2(n_644),
.C(n_594),
.Y(n_645)
);

BUFx24_ASAP7_75t_SL g646 ( 
.A(n_645),
.Y(n_646)
);

BUFx24_ASAP7_75t_SL g647 ( 
.A(n_646),
.Y(n_647)
);


endmodule