module fake_jpeg_23685_n_327 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_42),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_20),
.B1(n_24),
.B2(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_0),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_34),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_76),
.B1(n_85),
.B2(n_38),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_35),
.B(n_34),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_53),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_25),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_20),
.B1(n_35),
.B2(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_20),
.B1(n_37),
.B2(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_47),
.B1(n_35),
.B2(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_26),
.B(n_31),
.C(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_67),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_18),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_75),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_31),
.B1(n_25),
.B2(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_99),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_37),
.B1(n_33),
.B2(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_103),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_107),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_61),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_38),
.B1(n_30),
.B2(n_19),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_113),
.B1(n_94),
.B2(n_123),
.Y(n_148)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_111),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_53),
.A2(n_30),
.B1(n_19),
.B2(n_2),
.Y(n_113)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_122),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_48),
.B1(n_30),
.B2(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_54),
.B1(n_72),
.B2(n_87),
.Y(n_144)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_52),
.B1(n_86),
.B2(n_69),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_121),
.B1(n_94),
.B2(n_100),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_58),
.C(n_65),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_126),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_127),
.B(n_133),
.Y(n_184)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_135),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_66),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_4),
.B(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_0),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_1),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_148),
.B1(n_154),
.B2(n_104),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_54),
.A3(n_59),
.B1(n_80),
.B2(n_83),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_94),
.A2(n_72),
.B1(n_84),
.B2(n_3),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_1),
.B(n_2),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_4),
.B(n_7),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_182),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_161),
.B(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_106),
.B1(n_115),
.B2(n_88),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_144),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_90),
.B1(n_98),
.B2(n_103),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_64),
.B1(n_71),
.B2(n_8),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_168),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_64),
.B(n_102),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_166),
.B(n_188),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_112),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_191),
.B(n_133),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_131),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_173),
.A2(n_179),
.B1(n_152),
.B2(n_150),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_11),
.B(n_12),
.Y(n_221)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_155),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_112),
.B1(n_109),
.B2(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_9),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_9),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_125),
.A2(n_122),
.B(n_10),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_184),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_203),
.B1(n_207),
.B2(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_200),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_215),
.B1(n_203),
.B2(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_178),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_199),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_151),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_124),
.C(n_130),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_159),
.C(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_157),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_140),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_10),
.C(n_11),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_190),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_221),
.B(n_174),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_231),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_232),
.C(n_244),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_173),
.B1(n_170),
.B2(n_168),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_236),
.B1(n_205),
.B2(n_213),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_215),
.B1(n_198),
.B2(n_213),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_171),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_160),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_177),
.B1(n_160),
.B2(n_137),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_196),
.B1(n_197),
.B2(n_211),
.Y(n_264)
);

NAND4xp25_ASAP7_75t_SL g237 ( 
.A(n_195),
.B(n_127),
.C(n_185),
.D(n_129),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_192),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_196),
.Y(n_248)
);

NAND2x1_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_161),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_221),
.B(n_217),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_11),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_246),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_225),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_253),
.B(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_219),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_209),
.B1(n_212),
.B2(n_194),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_217),
.B1(n_193),
.B2(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.C(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_192),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_263),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_241),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_222),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_253),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_224),
.C(n_232),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_277),
.C(n_251),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_244),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_281),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_238),
.C(n_228),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_264),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_211),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_295),
.B(n_288),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_257),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_293),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_248),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_267),
.A2(n_247),
.B1(n_256),
.B2(n_255),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_286),
.B1(n_284),
.B2(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_276),
.C(n_266),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_265),
.C(n_238),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_295),
.C(n_207),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_270),
.B(n_228),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_235),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_278),
.B1(n_282),
.B2(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_235),
.C(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

AO221x1_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_280),
.B1(n_242),
.B2(n_275),
.C(n_272),
.Y(n_298)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_15),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_284),
.A2(n_269),
.B1(n_275),
.B2(n_245),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_304),
.B(n_15),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_14),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_289),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_14),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_12),
.C(n_13),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_310),
.B(n_313),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_13),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_296),
.B1(n_17),
.B2(n_16),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_301),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_317),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_299),
.B(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_312),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_296),
.B(n_303),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.C(n_316),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_319),
.A2(n_309),
.B(n_312),
.C(n_313),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_323),
.B(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_16),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_16),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_17),
.Y(n_327)
);


endmodule