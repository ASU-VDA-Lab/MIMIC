module fake_jpeg_29694_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_62),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_0),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_52),
.B1(n_43),
.B2(n_55),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_74),
.B1(n_51),
.B2(n_52),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_19),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_52),
.B1(n_54),
.B2(n_42),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_41),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_90),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_3),
.CI(n_4),
.CON(n_90),
.SN(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_3),
.B(n_4),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_5),
.B(n_6),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_14),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_106),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_39),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_21),
.B(n_23),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_30),
.B(n_31),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_25),
.B(n_27),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_117),
.B1(n_120),
.B2(n_97),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_103),
.C(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

AO221x1_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_96),
.B1(n_111),
.B2(n_112),
.C(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_103),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_124),
.B(n_118),
.C(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_124),
.Y(n_132)
);


endmodule