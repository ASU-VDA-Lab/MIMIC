module fake_jpeg_18699_n_273 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_33),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_32),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_19),
.B1(n_14),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_58),
.B1(n_37),
.B2(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_15),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_19),
.B1(n_31),
.B2(n_14),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_42),
.B1(n_37),
.B2(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_53),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_19),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_33),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_19),
.B1(n_14),
.B2(n_11),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_51),
.B1(n_57),
.B2(n_55),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_34),
.C(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_70),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_54),
.B1(n_51),
.B2(n_49),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_41),
.C(n_28),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_53),
.C(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_54),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_62),
.B1(n_83),
.B2(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_63),
.B(n_72),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_98),
.B(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_59),
.B(n_70),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_66),
.C(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_47),
.B1(n_56),
.B2(n_37),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_65),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_110),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_71),
.B(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_68),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_71),
.C(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_114),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_91),
.C(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_91),
.B1(n_67),
.B2(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_128),
.B1(n_47),
.B2(n_56),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_141),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_58),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_18),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_76),
.B1(n_78),
.B2(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_136),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_112),
.B1(n_98),
.B2(n_48),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_41),
.B(n_23),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_23),
.B(n_22),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_100),
.B1(n_112),
.B2(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_39),
.B1(n_69),
.B2(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_76),
.B1(n_43),
.B2(n_48),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_101),
.B1(n_108),
.B2(n_52),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_76),
.B1(n_56),
.B2(n_52),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_11),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_11),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_18),
.C(n_23),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_93),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_94),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_144),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_94),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_39),
.B(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_149),
.B1(n_153),
.B2(n_159),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_96),
.CI(n_106),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_126),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_108),
.B1(n_69),
.B2(n_35),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_108),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_124),
.B1(n_123),
.B2(n_142),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_165),
.B(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_47),
.B1(n_14),
.B2(n_36),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_162),
.B1(n_161),
.B2(n_152),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_144),
.C(n_134),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_123),
.A2(n_22),
.B(n_1),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_136),
.B(n_131),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_140),
.C(n_133),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_178),
.C(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_187),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_117),
.C(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_132),
.C(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_153),
.C(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_168),
.C(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_152),
.B1(n_170),
.B2(n_165),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_160),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_198),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_180),
.A2(n_147),
.B1(n_146),
.B2(n_156),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_202),
.C(n_208),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_204),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_170),
.B1(n_22),
.B2(n_12),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_27),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_28),
.C(n_27),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_208),
.C(n_196),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_219),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_215),
.C(n_17),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_195),
.A2(n_190),
.B(n_182),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_2),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_171),
.C(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_189),
.B1(n_175),
.B2(n_188),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_220),
.B1(n_200),
.B2(n_203),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_2),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_171),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_26),
.C(n_24),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_223),
.C(n_21),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_26),
.C(n_24),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_1),
.B(n_2),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_2),
.B(n_3),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_192),
.B(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_233),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_202),
.B1(n_4),
.B2(n_5),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_231),
.B(n_234),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_210),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_236),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_218),
.C(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_4),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_239),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_246),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_244),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_217),
.B1(n_214),
.B2(n_12),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_4),
.B(n_5),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_17),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_4),
.B(n_5),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_16),
.C(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_256),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_21),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_21),
.C(n_6),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_21),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_252),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_251),
.B(n_250),
.Y(n_264)
);

NAND4xp25_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_245),
.C(n_6),
.D(n_7),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_260),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_6),
.B(n_8),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_262),
.C(n_261),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_9),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_9),
.C(n_10),
.Y(n_273)
);


endmodule