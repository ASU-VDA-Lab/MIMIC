module fake_jpeg_18637_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NAND3xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_2),
.C(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx11_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_0),
.B(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_1),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_12),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_28),
.B1(n_24),
.B2(n_16),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_19),
.B1(n_25),
.B2(n_8),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_29),
.Y(n_46)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_47),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.C(n_40),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_49),
.C(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_48),
.Y(n_70)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_31),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_17),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_24),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_21),
.C(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_49),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_60)
);

A2O1A1O1Ixp25_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_25),
.B(n_19),
.C(n_9),
.D(n_11),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_4),
.B1(n_6),
.B2(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_6),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_45),
.Y(n_75)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_48),
.C(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_56),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_73),
.B1(n_68),
.B2(n_70),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_81),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.C(n_76),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_65),
.C(n_63),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_91),
.C(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_77),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_91),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_96),
.C(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_98),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_88),
.B(n_74),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_67),
.C(n_47),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);


endmodule