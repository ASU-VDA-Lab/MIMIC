module fake_netlist_6_3426_n_697 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_697);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_697;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_694;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_663;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_10),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_91),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_55),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_136),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_50),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_14),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_24),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_17),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_49),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_38),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_56),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_32),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_12),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_14),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_70),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_53),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_8),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_121),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_73),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_23),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_77),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_61),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_96),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_39),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_22),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_36),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

AOI22x1_ASAP7_75t_SL g192 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_176),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_1),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_2),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_159),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_3),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_160),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_18),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_19),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_9),
.B(n_10),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_182),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_221),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_190),
.Y(n_245)
);

AND3x2_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_160),
.C(n_188),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_153),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_20),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_189),
.B(n_185),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_144),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_145),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_21),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_146),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_222),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_205),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_193),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_252),
.B(n_208),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_238),
.B(n_256),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_193),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_203),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_261),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_246),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_253),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_219),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_232),
.B(n_223),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_247),
.B(n_223),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_210),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_213),
.B1(n_188),
.B2(n_198),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_206),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_262),
.A2(n_183),
.B1(n_161),
.B2(n_162),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_206),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g305 ( 
.A(n_248),
.B(n_224),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_267),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_237),
.B(n_204),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_229),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_204),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_199),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_244),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_262),
.A2(n_180),
.B1(n_163),
.B2(n_170),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_229),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_229),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_270),
.B(n_148),
.Y(n_321)
);

BUFx6f_ASAP7_75t_SL g322 ( 
.A(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_233),
.B(n_258),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_229),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_230),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_230),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_174),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_255),
.B(n_178),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_282),
.A2(n_217),
.B(n_263),
.C(n_236),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_306),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_278),
.A2(n_265),
.B(n_264),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_277),
.A2(n_290),
.B(n_292),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_283),
.A2(n_234),
.B(n_239),
.C(n_236),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_224),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g347 ( 
.A1(n_305),
.A2(n_235),
.B(n_224),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_253),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_286),
.B(n_197),
.C(n_196),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_288),
.A2(n_253),
.B1(n_179),
.B2(n_230),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_230),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_192),
.Y(n_354)
);

CKINVDCx8_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_196),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_195),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_284),
.B(n_11),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_195),
.B(n_12),
.C(n_13),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_25),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_26),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_307),
.A2(n_85),
.B(n_139),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_294),
.Y(n_367)
);

BUFx4f_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_287),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_86),
.B(n_137),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_302),
.A2(n_82),
.B1(n_135),
.B2(n_27),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_296),
.B(n_15),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_16),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_320),
.A2(n_87),
.B(n_28),
.Y(n_375)
);

AOI21xp33_ASAP7_75t_L g376 ( 
.A1(n_316),
.A2(n_16),
.B(n_140),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_29),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_299),
.B(n_30),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_300),
.B(n_31),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_333),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_309),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_382)
);

OAI321xp33_ASAP7_75t_L g383 ( 
.A1(n_309),
.A2(n_37),
.A3(n_40),
.B1(n_41),
.B2(n_42),
.C(n_43),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_327),
.A2(n_44),
.B(n_45),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_311),
.B(n_325),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_46),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_329),
.B(n_47),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_L g390 ( 
.A1(n_326),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_327),
.A2(n_54),
.B(n_57),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_318),
.B(n_58),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_318),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_330),
.B(n_328),
.Y(n_394)
);

AO31x2_ASAP7_75t_L g395 ( 
.A1(n_348),
.A2(n_319),
.A3(n_300),
.B(n_322),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_335),
.B(n_300),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_342),
.A2(n_300),
.B(n_322),
.Y(n_398)
);

O2A1O1Ixp5_ASAP7_75t_L g399 ( 
.A1(n_353),
.A2(n_300),
.B(n_60),
.C(n_62),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_368),
.A2(n_59),
.B(n_65),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_338),
.A2(n_67),
.B(n_69),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_71),
.B(n_72),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_358),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_78),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_354),
.A2(n_79),
.B(n_80),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_88),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_368),
.A2(n_90),
.B(n_92),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_357),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_345),
.A2(n_93),
.B(n_94),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_355),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_100),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_377),
.A2(n_134),
.B(n_103),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_345),
.A2(n_102),
.B(n_104),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_107),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_367),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_369),
.B(n_108),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_352),
.A2(n_109),
.B(n_110),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_337),
.A2(n_111),
.B(n_112),
.Y(n_421)
);

AND3x4_ASAP7_75t_L g422 ( 
.A(n_350),
.B(n_351),
.C(n_334),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_386),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_337),
.A2(n_113),
.B(n_114),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_344),
.A2(n_391),
.B(n_380),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_378),
.A2(n_133),
.B(n_117),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_381),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_383),
.A2(n_115),
.B(n_118),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_336),
.B(n_349),
.Y(n_429)
);

AO31x2_ASAP7_75t_L g430 ( 
.A1(n_390),
.A2(n_375),
.A3(n_372),
.B(n_388),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_336),
.B(n_119),
.Y(n_431)
);

AOI21xp33_ASAP7_75t_L g432 ( 
.A1(n_359),
.A2(n_126),
.B(n_127),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_346),
.A2(n_129),
.B(n_130),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_346),
.B(n_132),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_392),
.A2(n_374),
.B(n_379),
.Y(n_436)
);

AO31x2_ASAP7_75t_L g437 ( 
.A1(n_362),
.A2(n_364),
.A3(n_385),
.B(n_370),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_371),
.A2(n_373),
.B(n_382),
.C(n_366),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_393),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_360),
.A2(n_363),
.B(n_389),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_360),
.A2(n_363),
.B(n_347),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_360),
.A2(n_290),
.B(n_277),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_363),
.B(n_340),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_397),
.Y(n_446)
);

BUFx2_ASAP7_75t_R g447 ( 
.A(n_417),
.Y(n_447)
);

AO21x2_ASAP7_75t_L g448 ( 
.A1(n_425),
.A2(n_438),
.B(n_410),
.Y(n_448)
);

AO21x2_ASAP7_75t_L g449 ( 
.A1(n_401),
.A2(n_398),
.B(n_432),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_422),
.A2(n_406),
.B1(n_419),
.B2(n_428),
.Y(n_450)
);

AOI22x1_ASAP7_75t_L g451 ( 
.A1(n_443),
.A2(n_416),
.B1(n_420),
.B2(n_423),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_413),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_415),
.A2(n_426),
.B(n_431),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_399),
.A2(n_396),
.B(n_435),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_403),
.B(n_411),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_441),
.A2(n_440),
.B(n_408),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_402),
.A2(n_400),
.B(n_407),
.Y(n_460)
);

O2A1O1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_405),
.A2(n_427),
.B(n_433),
.C(n_404),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_444),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_402),
.A2(n_424),
.B(n_434),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_395),
.B(n_437),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_395),
.A2(n_437),
.B(n_430),
.Y(n_467)
);

NAND2x1p5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_395),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_404),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_412),
.A2(n_396),
.B(n_342),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_437),
.A2(n_436),
.B(n_394),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_409),
.B(n_335),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_427),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

AO21x2_ASAP7_75t_L g478 ( 
.A1(n_425),
.A2(n_438),
.B(n_410),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_425),
.A2(n_410),
.B(n_394),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_425),
.A2(n_410),
.B(n_394),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_282),
.C(n_210),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_409),
.A2(n_283),
.B(n_282),
.C(n_372),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_484),
.A2(n_471),
.B(n_473),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_472),
.A2(n_449),
.B(n_478),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_467),
.A2(n_472),
.B(n_469),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_449),
.A2(n_478),
.B(n_448),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

AO21x2_ASAP7_75t_L g497 ( 
.A1(n_449),
.A2(n_448),
.B(n_478),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_455),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_481),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_463),
.Y(n_502)
);

CKINVDCx6p67_ASAP7_75t_R g503 ( 
.A(n_445),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_450),
.B(n_483),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_452),
.A2(n_448),
.B1(n_470),
.B2(n_464),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_462),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_452),
.A2(n_447),
.B1(n_459),
.B2(n_451),
.Y(n_507)
);

CKINVDCx12_ASAP7_75t_R g508 ( 
.A(n_445),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_468),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_468),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_464),
.A2(n_451),
.B1(n_457),
.B2(n_479),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_445),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_461),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_504),
.A2(n_464),
.B1(n_457),
.B2(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_492),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_511),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_506),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_486),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_495),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_486),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_482),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_489),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_504),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_482),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_464),
.Y(n_533)
);

NAND2x1_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_457),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_464),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_509),
.B(n_479),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_458),
.B1(n_479),
.B2(n_456),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_466),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_456),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_509),
.B(n_456),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_503),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_503),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_502),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_509),
.B(n_460),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_509),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_494),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_490),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_496),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_544),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_548),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_493),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_546),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_531),
.B(n_493),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_535),
.B(n_505),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_516),
.B(n_496),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_547),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_516),
.B(n_497),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_519),
.B(n_507),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_527),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_537),
.B(n_497),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_497),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_528),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_547),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_544),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_530),
.B(n_509),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_533),
.B(n_509),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_521),
.B(n_488),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_522),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_551),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_522),
.B(n_488),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_526),
.B(n_488),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_518),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_551),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_512),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_525),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_525),
.B(n_512),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_540),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_526),
.B(n_510),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_557),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_561),
.Y(n_586)
);

HB1xp67_ASAP7_75t_SL g587 ( 
.A(n_569),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_573),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_580),
.B(n_544),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_561),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_568),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_556),
.B(n_541),
.Y(n_592)
);

NOR2x1_ASAP7_75t_SL g593 ( 
.A(n_560),
.B(n_548),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_552),
.B(n_519),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_564),
.B(n_549),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_580),
.B(n_549),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_556),
.B(n_541),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_575),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_558),
.B(n_532),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_580),
.B(n_536),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_555),
.B(n_545),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_579),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_571),
.B(n_517),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_555),
.B(n_545),
.Y(n_607)
);

AND2x4_ASAP7_75t_SL g608 ( 
.A(n_555),
.B(n_539),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_517),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_579),
.Y(n_610)
);

AOI21x1_ASAP7_75t_L g611 ( 
.A1(n_563),
.A2(n_534),
.B(n_538),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_588),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_558),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

OAI21xp33_ASAP7_75t_L g615 ( 
.A1(n_609),
.A2(n_562),
.B(n_559),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_594),
.B(n_562),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_591),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_592),
.B(n_565),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_565),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_606),
.B(n_555),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_597),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_600),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_604),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_605),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_621),
.A2(n_585),
.B(n_595),
.Y(n_626)
);

AOI221xp5_ASAP7_75t_L g627 ( 
.A1(n_615),
.A2(n_599),
.B1(n_602),
.B2(n_598),
.C(n_610),
.Y(n_627)
);

AND2x4_ASAP7_75t_SL g628 ( 
.A(n_619),
.B(n_589),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_614),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_614),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_621),
.B(n_612),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_616),
.B(n_536),
.Y(n_632)
);

OAI31xp33_ASAP7_75t_L g633 ( 
.A1(n_612),
.A2(n_559),
.A3(n_520),
.B(n_553),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_623),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_623),
.Y(n_635)
);

INVx8_ASAP7_75t_L g636 ( 
.A(n_631),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_628),
.B(n_596),
.Y(n_637)
);

OAI32xp33_ASAP7_75t_L g638 ( 
.A1(n_626),
.A2(n_613),
.A3(n_624),
.B1(n_622),
.B2(n_625),
.Y(n_638)
);

AOI21xp33_ASAP7_75t_L g639 ( 
.A1(n_632),
.A2(n_599),
.B(n_618),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_629),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_638),
.A2(n_627),
.B1(n_631),
.B2(n_634),
.C(n_630),
.Y(n_641)
);

AOI221xp5_ASAP7_75t_L g642 ( 
.A1(n_639),
.A2(n_617),
.B1(n_633),
.B2(n_635),
.C(n_620),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_640),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_636),
.B(n_633),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_636),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_637),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_SL g647 ( 
.A(n_644),
.B(n_520),
.C(n_587),
.Y(n_647)
);

OA22x2_ASAP7_75t_L g648 ( 
.A1(n_645),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_646),
.B(n_578),
.C(n_570),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_643),
.Y(n_650)
);

OAI21xp33_ASAP7_75t_SL g651 ( 
.A1(n_648),
.A2(n_650),
.B(n_647),
.Y(n_651)
);

NAND2x1_ASAP7_75t_SL g652 ( 
.A(n_649),
.B(n_587),
.Y(n_652)
);

NOR2x1_ASAP7_75t_L g653 ( 
.A(n_650),
.B(n_489),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_653),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_651),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_652),
.B(n_542),
.C(n_543),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_651),
.A2(n_603),
.B1(n_607),
.B2(n_608),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_654),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_655),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_657),
.B(n_543),
.C(n_542),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_656),
.B(n_555),
.C(n_583),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_655),
.Y(n_662)
);

NOR4xp25_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_514),
.C(n_583),
.D(n_523),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_L g664 ( 
.A(n_654),
.B(n_611),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_655),
.A2(n_607),
.B1(n_603),
.B2(n_608),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_658),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_659),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_662),
.Y(n_668)
);

AOI221xp5_ASAP7_75t_SL g669 ( 
.A1(n_663),
.A2(n_598),
.B1(n_584),
.B2(n_582),
.C(n_573),
.Y(n_669)
);

NAND4xp75_ASAP7_75t_L g670 ( 
.A(n_664),
.B(n_514),
.C(n_508),
.D(n_582),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_665),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_661),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_660),
.A2(n_508),
.B1(n_603),
.B2(n_607),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_667),
.Y(n_674)
);

OAI211xp5_ASAP7_75t_L g675 ( 
.A1(n_668),
.A2(n_489),
.B(n_513),
.C(n_460),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_671),
.A2(n_465),
.B(n_453),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_666),
.Y(n_677)
);

OA22x2_ASAP7_75t_L g678 ( 
.A1(n_672),
.A2(n_588),
.B1(n_572),
.B2(n_554),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_670),
.Y(n_679)
);

OAI22x1_ASAP7_75t_L g680 ( 
.A1(n_673),
.A2(n_559),
.B1(n_572),
.B2(n_529),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_674),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_673),
.B(n_669),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_677),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_676),
.A2(n_465),
.B(n_453),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_SL g685 ( 
.A1(n_678),
.A2(n_680),
.B1(n_675),
.B2(n_529),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_683),
.B(n_529),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_681),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_682),
.A2(n_584),
.B1(n_572),
.B2(n_566),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_685),
.Y(n_689)
);

INVxp33_ASAP7_75t_SL g690 ( 
.A(n_687),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_689),
.A2(n_684),
.B1(n_566),
.B2(n_576),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_SL g692 ( 
.A1(n_686),
.A2(n_684),
.B1(n_593),
.B2(n_523),
.Y(n_692)
);

AOI21xp33_ASAP7_75t_SL g693 ( 
.A1(n_690),
.A2(n_688),
.B(n_577),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_691),
.A2(n_577),
.B1(n_581),
.B2(n_574),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_694),
.A2(n_692),
.B(n_534),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_695),
.B(n_693),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_696),
.A2(n_581),
.B1(n_554),
.B2(n_574),
.Y(n_697)
);


endmodule