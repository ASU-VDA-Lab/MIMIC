module real_aes_9213_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g541 ( .A1(n_0), .A2(n_189), .B(n_542), .C(n_545), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_1), .B(n_530), .Y(n_546) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_3), .A2(n_751), .B1(n_754), .B2(n_755), .Y(n_750) );
INVx1_ASAP7_75t_L g755 ( .A(n_3), .Y(n_755) );
INVx1_ASAP7_75t_L g207 ( .A(n_4), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_5), .B(n_178), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_6), .A2(n_445), .B(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_7), .A2(n_154), .B(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_8), .A2(n_36), .B1(n_134), .B2(n_143), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_9), .B(n_154), .Y(n_218) );
AND2x6_ASAP7_75t_L g152 ( .A(n_10), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_11), .A2(n_152), .B(n_448), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_12), .B(n_37), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_12), .B(n_37), .Y(n_434) );
INVx1_ASAP7_75t_L g150 ( .A(n_13), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_14), .B(n_141), .Y(n_161) );
INVx1_ASAP7_75t_L g199 ( .A(n_15), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_16), .B(n_178), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_17), .B(n_155), .Y(n_223) );
AO32x2_ASAP7_75t_L g186 ( .A1(n_18), .A2(n_151), .A3(n_154), .B1(n_187), .B2(n_191), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_19), .B(n_143), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_20), .B(n_155), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_21), .A2(n_53), .B1(n_134), .B2(n_143), .Y(n_190) );
AOI22xp33_ASAP7_75t_SL g140 ( .A1(n_22), .A2(n_82), .B1(n_141), .B2(n_143), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_23), .B(n_143), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_24), .A2(n_151), .B(n_448), .C(n_450), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_25), .A2(n_151), .B(n_448), .C(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_26), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_27), .B(n_146), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_28), .A2(n_445), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_29), .B(n_146), .Y(n_184) );
INVx2_ASAP7_75t_L g136 ( .A(n_30), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_31), .A2(n_469), .B(n_478), .C(n_480), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_32), .B(n_143), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_33), .B(n_146), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_34), .A2(n_74), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_34), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_35), .B(n_163), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_38), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_39), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_40), .B(n_178), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_41), .B(n_445), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_42), .A2(n_469), .B(n_478), .C(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_43), .A2(n_124), .B1(n_428), .B2(n_429), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_43), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_43), .A2(n_80), .B1(n_428), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_44), .A2(n_103), .B1(n_116), .B2(n_762), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_45), .B(n_143), .Y(n_213) );
INVx1_ASAP7_75t_L g543 ( .A(n_46), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_47), .A2(n_90), .B1(n_134), .B2(n_137), .Y(n_133) );
INVx1_ASAP7_75t_L g516 ( .A(n_48), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_49), .B(n_143), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_50), .B(n_143), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_51), .B(n_445), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_52), .B(n_205), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g227 ( .A1(n_54), .A2(n_59), .B1(n_141), .B2(n_143), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_55), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_56), .B(n_143), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_57), .B(n_143), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_58), .Y(n_759) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_61), .B(n_445), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_62), .B(n_530), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_63), .A2(n_202), .B(n_205), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_64), .B(n_143), .Y(n_208) );
INVx1_ASAP7_75t_L g149 ( .A(n_65), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_66), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_67), .B(n_178), .Y(n_482) );
AO32x2_ASAP7_75t_L g131 ( .A1(n_68), .A2(n_132), .A3(n_145), .B1(n_151), .B2(n_154), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_69), .B(n_144), .Y(n_506) );
INVx1_ASAP7_75t_L g241 ( .A(n_70), .Y(n_241) );
INVx1_ASAP7_75t_L g176 ( .A(n_71), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_72), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_73), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_75), .A2(n_448), .B(n_465), .C(n_469), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_76), .B(n_141), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_77), .Y(n_525) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_79), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_80), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_81), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_83), .B(n_134), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_84), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_85), .B(n_141), .Y(n_181) );
INVx2_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_87), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_88), .B(n_138), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_89), .B(n_141), .Y(n_214) );
INVx2_ASAP7_75t_L g112 ( .A(n_91), .Y(n_112) );
OR2x2_ASAP7_75t_L g432 ( .A(n_91), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g749 ( .A(n_91), .B(n_743), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_92), .A2(n_101), .B1(n_141), .B2(n_142), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_93), .B(n_445), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_94), .Y(n_481) );
INVxp67_ASAP7_75t_L g528 ( .A(n_95), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_96), .B(n_141), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g466 ( .A(n_98), .Y(n_466) );
INVx1_ASAP7_75t_L g502 ( .A(n_99), .Y(n_502) );
AND2x2_ASAP7_75t_L g518 ( .A(n_100), .B(n_146), .Y(n_518) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g762 ( .A(n_105), .Y(n_762) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g433 ( .A(n_111), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g730 ( .A(n_112), .B(n_433), .Y(n_730) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_112), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO221x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_744), .B1(n_747), .B2(n_756), .C(n_758), .Y(n_116) );
OAI222xp33_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_121), .B1(n_731), .B2(n_732), .C1(n_738), .C2(n_739), .Y(n_117) );
INVx1_ASAP7_75t_L g731 ( .A(n_118), .Y(n_731) );
INVxp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_430), .B1(n_435), .B2(n_728), .Y(n_122) );
INVx1_ASAP7_75t_L g734 ( .A(n_123), .Y(n_734) );
INVx2_ASAP7_75t_L g429 ( .A(n_124), .Y(n_429) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XOR2x2_ASAP7_75t_L g751 ( .A(n_125), .B(n_752), .Y(n_751) );
AND3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_348), .C(n_396), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_276), .C(n_321), .D(n_335), .Y(n_126) );
OAI311xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_192), .A3(n_219), .B1(n_229), .C1(n_244), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_156), .Y(n_128) );
OAI21xp33_ASAP7_75t_L g229 ( .A1(n_129), .A2(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g337 ( .A(n_129), .B(n_264), .Y(n_337) );
AND2x2_ASAP7_75t_L g394 ( .A(n_129), .B(n_280), .Y(n_394) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g287 ( .A(n_130), .B(n_185), .Y(n_287) );
AND2x2_ASAP7_75t_L g344 ( .A(n_130), .B(n_292), .Y(n_344) );
INVx1_ASAP7_75t_L g385 ( .A(n_130), .Y(n_385) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_131), .Y(n_253) );
AND2x2_ASAP7_75t_L g294 ( .A(n_131), .B(n_185), .Y(n_294) );
AND2x2_ASAP7_75t_L g298 ( .A(n_131), .B(n_186), .Y(n_298) );
INVx1_ASAP7_75t_L g310 ( .A(n_131), .Y(n_310) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_138), .B1(n_140), .B2(n_144), .Y(n_132) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx3_ASAP7_75t_L g137 ( .A(n_135), .Y(n_137) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
AND2x6_ASAP7_75t_L g448 ( .A(n_135), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_137), .Y(n_483) );
INVx2_ASAP7_75t_L g545 ( .A(n_137), .Y(n_545) );
INVx2_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_138), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_138), .A2(n_189), .B1(n_226), .B2(n_227), .Y(n_225) );
INVx4_ASAP7_75t_L g544 ( .A(n_138), .Y(n_544) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g144 ( .A(n_139), .Y(n_144) );
INVx1_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
AND2x2_ASAP7_75t_L g446 ( .A(n_139), .B(n_206), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_139), .Y(n_449) );
INVx2_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_143), .Y(n_468) );
INVx5_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
INVx1_ASAP7_75t_L g455 ( .A(n_145), .Y(n_455) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_146), .A2(n_158), .B(n_168), .Y(n_157) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_146), .A2(n_173), .B(n_184), .Y(n_172) );
INVx1_ASAP7_75t_L g458 ( .A(n_146), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_146), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_146), .A2(n_513), .B(n_514), .Y(n_512) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x2_ASAP7_75t_L g155 ( .A(n_147), .B(n_148), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NAND3xp33_ASAP7_75t_L g224 ( .A(n_151), .B(n_225), .C(n_228), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_151), .A2(n_237), .B(n_240), .Y(n_236) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g158 ( .A1(n_152), .A2(n_159), .B(n_164), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_152), .A2(n_174), .B(n_179), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_152), .A2(n_198), .B(n_203), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_152), .A2(n_212), .B(n_215), .Y(n_211) );
AND2x4_ASAP7_75t_L g445 ( .A(n_152), .B(n_446), .Y(n_445) );
INVx4_ASAP7_75t_SL g470 ( .A(n_152), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_152), .B(n_446), .Y(n_503) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_154), .A2(n_211), .B(n_218), .Y(n_210) );
INVx4_ASAP7_75t_L g228 ( .A(n_154), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_154), .A2(n_493), .B(n_494), .Y(n_492) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_154), .Y(n_522) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_169), .Y(n_156) );
AND2x2_ASAP7_75t_L g231 ( .A(n_157), .B(n_185), .Y(n_231) );
INVx2_ASAP7_75t_L g265 ( .A(n_157), .Y(n_265) );
AND2x2_ASAP7_75t_L g280 ( .A(n_157), .B(n_186), .Y(n_280) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_157), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_157), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g300 ( .A(n_157), .B(n_263), .Y(n_300) );
INVx1_ASAP7_75t_L g312 ( .A(n_157), .Y(n_312) );
INVx1_ASAP7_75t_L g353 ( .A(n_157), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_157), .B(n_253), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .Y(n_164) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_167), .A2(n_204), .B(n_241), .C(n_242), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g169 ( .A(n_170), .B(n_185), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g230 ( .A(n_171), .B(n_231), .Y(n_230) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_171), .Y(n_258) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_171), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g315 ( .A(n_171), .B(n_185), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_171), .B(n_310), .Y(n_373) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g263 ( .A(n_172), .Y(n_263) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_172), .Y(n_279) );
OR2x2_ASAP7_75t_L g352 ( .A(n_172), .B(n_353), .Y(n_352) );
O2A1O1Ixp5_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_178), .Y(n_174) );
INVx2_ASAP7_75t_L g189 ( .A(n_178), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_178), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_178), .A2(n_238), .B(n_239), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_178), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g452 ( .A(n_183), .Y(n_452) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx2_ASAP7_75t_L g259 ( .A(n_186), .Y(n_259) );
AND2x2_ASAP7_75t_L g264 ( .A(n_186), .B(n_265), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_189), .A2(n_204), .B(n_207), .C(n_208), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_189), .A2(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g196 ( .A(n_191), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_191), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_192), .B(n_247), .Y(n_410) );
INVx1_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_L g380 ( .A(n_193), .B(n_221), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_210), .Y(n_193) );
AND2x2_ASAP7_75t_L g256 ( .A(n_194), .B(n_247), .Y(n_256) );
INVx2_ASAP7_75t_L g268 ( .A(n_194), .Y(n_268) );
AND2x2_ASAP7_75t_L g302 ( .A(n_194), .B(n_250), .Y(n_302) );
AND2x2_ASAP7_75t_L g369 ( .A(n_194), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_195), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g249 ( .A(n_195), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g289 ( .A(n_195), .B(n_210), .Y(n_289) );
AND2x2_ASAP7_75t_L g306 ( .A(n_195), .B(n_307), .Y(n_306) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_209), .Y(n_195) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_196), .A2(n_236), .B(n_243), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .C(n_202), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_200), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_200), .A2(n_506), .B(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_202), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_204), .A2(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g232 ( .A(n_210), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g250 ( .A(n_210), .Y(n_250) );
AND2x2_ASAP7_75t_L g255 ( .A(n_210), .B(n_235), .Y(n_255) );
AND2x2_ASAP7_75t_L g328 ( .A(n_210), .B(n_307), .Y(n_328) );
AND2x2_ASAP7_75t_L g393 ( .A(n_210), .B(n_383), .Y(n_393) );
OAI311xp33_ASAP7_75t_L g276 ( .A1(n_219), .A2(n_277), .A3(n_281), .B1(n_283), .C1(n_303), .Y(n_276) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g288 ( .A(n_220), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g347 ( .A(n_220), .B(n_255), .Y(n_347) );
AND2x2_ASAP7_75t_L g421 ( .A(n_220), .B(n_302), .Y(n_421) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_221), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g356 ( .A(n_221), .Y(n_356) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
NOR2x1_ASAP7_75t_L g319 ( .A(n_222), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g376 ( .A(n_222), .B(n_250), .Y(n_376) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
AO21x1_ASAP7_75t_L g272 ( .A1(n_225), .A2(n_228), .B(n_273), .Y(n_272) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_228), .A2(n_463), .B(n_472), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_228), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_228), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_228), .A2(n_501), .B(n_508), .Y(n_500) );
INVx3_ASAP7_75t_L g530 ( .A(n_228), .Y(n_530) );
AND2x2_ASAP7_75t_L g251 ( .A(n_231), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g304 ( .A(n_231), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g384 ( .A(n_231), .B(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_232), .A2(n_264), .B1(n_284), .B2(n_288), .C(n_290), .Y(n_283) );
INVx1_ASAP7_75t_L g408 ( .A(n_233), .Y(n_408) );
OR2x2_ASAP7_75t_L g374 ( .A(n_234), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g269 ( .A(n_235), .B(n_250), .Y(n_269) );
OR2x2_ASAP7_75t_L g271 ( .A(n_235), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
INVx2_ASAP7_75t_L g307 ( .A(n_235), .Y(n_307) );
AND2x2_ASAP7_75t_L g334 ( .A(n_235), .B(n_272), .Y(n_334) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_235), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_251), .B1(n_254), .B2(n_257), .C(n_260), .Y(n_244) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g345 ( .A(n_247), .B(n_255), .Y(n_345) );
AND2x2_ASAP7_75t_L g395 ( .A(n_247), .B(n_249), .Y(n_395) );
INVx2_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g282 ( .A(n_249), .B(n_253), .Y(n_282) );
AND2x2_ASAP7_75t_L g361 ( .A(n_249), .B(n_334), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_250), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
OAI21xp33_ASAP7_75t_L g330 ( .A1(n_251), .A2(n_331), .B(n_333), .Y(n_330) );
OR2x2_ASAP7_75t_L g274 ( .A(n_252), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g340 ( .A(n_252), .B(n_300), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_252), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g317 ( .A(n_253), .B(n_286), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_253), .B(n_400), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_254), .B(n_280), .Y(n_390) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g313 ( .A(n_255), .B(n_268), .Y(n_313) );
INVx1_ASAP7_75t_L g329 ( .A(n_256), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_266), .B1(n_270), .B2(n_274), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
INVx1_ASAP7_75t_L g305 ( .A(n_263), .Y(n_305) );
INVx1_ASAP7_75t_L g275 ( .A(n_264), .Y(n_275) );
AND2x2_ASAP7_75t_L g346 ( .A(n_264), .B(n_292), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_264), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
OR2x2_ASAP7_75t_L g270 ( .A(n_267), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_267), .B(n_383), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_267), .B(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g417 ( .A(n_269), .B(n_369), .Y(n_417) );
INVx1_ASAP7_75t_SL g383 ( .A(n_271), .Y(n_383) );
AND2x2_ASAP7_75t_L g323 ( .A(n_272), .B(n_307), .Y(n_323) );
INVx1_ASAP7_75t_L g370 ( .A(n_272), .Y(n_370) );
OAI222xp33_ASAP7_75t_L g411 ( .A1(n_277), .A2(n_367), .B1(n_412), .B2(n_413), .C1(n_416), .C2(n_418), .Y(n_411) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
AND2x2_ASAP7_75t_L g343 ( .A(n_280), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_280), .B(n_385), .Y(n_412) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_282), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g387 ( .A(n_284), .Y(n_387) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g325 ( .A(n_287), .Y(n_325) );
AND2x2_ASAP7_75t_L g404 ( .A(n_287), .B(n_365), .Y(n_404) );
AND2x2_ASAP7_75t_L g427 ( .A(n_287), .B(n_311), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_289), .B(n_323), .Y(n_322) );
OAI32xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .A3(n_295), .B1(n_297), .B2(n_301), .Y(n_290) );
BUFx2_ASAP7_75t_L g365 ( .A(n_292), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_293), .B(n_311), .Y(n_392) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g331 ( .A(n_294), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g399 ( .A(n_294), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g388 ( .A(n_295), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g359 ( .A(n_298), .B(n_332), .Y(n_359) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OAI221xp5_ASAP7_75t_SL g321 ( .A1(n_300), .A2(n_322), .B1(n_324), .B2(n_326), .C(n_330), .Y(n_321) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g333 ( .A(n_302), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g339 ( .A(n_302), .B(n_323), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_306), .B1(n_308), .B2(n_313), .C(n_314), .Y(n_303) );
INVx1_ASAP7_75t_L g422 ( .A(n_304), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_305), .B(n_399), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_306), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_311), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g377 ( .A(n_311), .Y(n_377) );
BUFx3_ASAP7_75t_L g400 ( .A(n_312), .Y(n_400) );
INVx1_ASAP7_75t_SL g341 ( .A(n_313), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_313), .B(n_355), .Y(n_354) );
AOI21xp33_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_316), .B(n_318), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_315), .A2(n_416), .B1(n_420), .B2(n_422), .C(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g362 ( .A(n_320), .B(n_323), .Y(n_362) );
INVx1_ASAP7_75t_L g426 ( .A(n_320), .Y(n_426) );
INVx2_ASAP7_75t_L g415 ( .A(n_323), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_323), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g368 ( .A(n_328), .B(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_338), .B1(n_340), .B2(n_341), .C(n_342), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B1(n_346), .B2(n_347), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_344), .A2(n_406), .B1(n_407), .B2(n_409), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_347), .A2(n_424), .B(n_427), .Y(n_423) );
NOR4xp25_ASAP7_75t_SL g348 ( .A(n_349), .B(n_357), .C(n_366), .D(n_386), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_363), .B2(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_374), .B2(n_377), .C(n_378), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g389 ( .A(n_369), .Y(n_389) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI21xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_381), .B(n_384), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_390), .C(n_391), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_394), .B2(n_395), .Y(n_391) );
CKINVDCx14_ASAP7_75t_R g401 ( .A(n_395), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_411), .C(n_419), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B1(n_402), .B2(n_403), .C(n_405), .Y(n_397) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g735 ( .A(n_431), .Y(n_735) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g743 ( .A(n_433), .Y(n_743) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g736 ( .A(n_436), .Y(n_736) );
AND3x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_632), .C(n_689), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_577), .C(n_613), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_486), .B(n_532), .C(n_564), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_459), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g535 ( .A(n_441), .B(n_536), .Y(n_535) );
INVx5_ASAP7_75t_L g563 ( .A(n_441), .Y(n_563) );
AND2x2_ASAP7_75t_L g636 ( .A(n_441), .B(n_552), .Y(n_636) );
AND2x2_ASAP7_75t_L g674 ( .A(n_441), .B(n_580), .Y(n_674) );
AND2x2_ASAP7_75t_L g694 ( .A(n_441), .B(n_537), .Y(n_694) );
OR2x6_ASAP7_75t_L g441 ( .A(n_442), .B(n_456), .Y(n_441) );
AOI21xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_447), .B(n_455), .Y(n_442) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx5_ASAP7_75t_L g479 ( .A(n_448), .Y(n_479) );
INVx2_ASAP7_75t_L g454 ( .A(n_452), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_454), .A2(n_481), .B(n_482), .C(n_483), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_454), .A2(n_483), .B(n_516), .C(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_459), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_460), .Y(n_575) );
AND2x2_ASAP7_75t_L g589 ( .A(n_460), .B(n_536), .Y(n_589) );
INVx1_ASAP7_75t_L g612 ( .A(n_460), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_460), .B(n_563), .Y(n_651) );
OR2x2_ASAP7_75t_L g688 ( .A(n_460), .B(n_534), .Y(n_688) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_461), .Y(n_624) );
AND2x2_ASAP7_75t_L g631 ( .A(n_461), .B(n_537), .Y(n_631) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g552 ( .A(n_462), .B(n_537), .Y(n_552) );
BUFx2_ASAP7_75t_L g580 ( .A(n_462), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_470), .A2(n_479), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g539 ( .A1(n_470), .A2(n_479), .B(n_540), .C(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
BUFx2_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
AND2x2_ASAP7_75t_L g713 ( .A(n_474), .B(n_567), .Y(n_713) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_519), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_488), .A2(n_614), .B1(n_621), .B2(n_622), .C(n_625), .Y(n_613) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
AND2x2_ASAP7_75t_L g520 ( .A(n_489), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_489), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g548 ( .A(n_490), .B(n_499), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_490), .B(n_500), .Y(n_558) );
OR2x2_ASAP7_75t_L g569 ( .A(n_490), .B(n_521), .Y(n_569) );
AND2x2_ASAP7_75t_L g572 ( .A(n_490), .B(n_560), .Y(n_572) );
AND2x2_ASAP7_75t_L g588 ( .A(n_490), .B(n_510), .Y(n_588) );
OR2x2_ASAP7_75t_L g604 ( .A(n_490), .B(n_500), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_490), .B(n_521), .Y(n_666) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_491), .B(n_510), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_491), .B(n_500), .Y(n_661) );
OR2x2_ASAP7_75t_L g582 ( .A(n_498), .B(n_569), .Y(n_582) );
INVx2_ASAP7_75t_L g608 ( .A(n_498), .Y(n_608) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
AND2x2_ASAP7_75t_L g531 ( .A(n_499), .B(n_511), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_499), .B(n_521), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_499), .B(n_511), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_499), .B(n_560), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_499), .A2(n_691), .B1(n_693), .B2(n_695), .C(n_698), .Y(n_690) );
INVx5_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_500), .B(n_521), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_510), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_510), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g576 ( .A(n_510), .B(n_548), .Y(n_576) );
OR2x2_ASAP7_75t_L g620 ( .A(n_510), .B(n_521), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_510), .B(n_572), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_510), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g685 ( .A(n_510), .B(n_686), .Y(n_685) );
INVx5_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_SL g549 ( .A(n_511), .B(n_520), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_511), .A2(n_554), .B(n_557), .C(n_561), .Y(n_553) );
OR2x2_ASAP7_75t_L g591 ( .A(n_511), .B(n_587), .Y(n_591) );
OR2x2_ASAP7_75t_L g627 ( .A(n_511), .B(n_569), .Y(n_627) );
OAI311xp33_ASAP7_75t_L g633 ( .A1(n_511), .A2(n_572), .A3(n_634), .B1(n_637), .C1(n_644), .Y(n_633) );
AND2x2_ASAP7_75t_L g684 ( .A(n_511), .B(n_521), .Y(n_684) );
AND2x2_ASAP7_75t_L g692 ( .A(n_511), .B(n_547), .Y(n_692) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_511), .Y(n_710) );
AND2x2_ASAP7_75t_L g727 ( .A(n_511), .B(n_548), .Y(n_727) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
AND2x2_ASAP7_75t_L g555 ( .A(n_520), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g711 ( .A(n_520), .Y(n_711) );
AND2x2_ASAP7_75t_L g547 ( .A(n_521), .B(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g560 ( .A(n_521), .Y(n_560) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_521), .Y(n_603) );
INVxp67_ASAP7_75t_L g642 ( .A(n_521), .Y(n_642) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_529), .Y(n_521) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_530), .A2(n_538), .B(n_546), .Y(n_537) );
AND2x2_ASAP7_75t_L g720 ( .A(n_531), .B(n_568), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_547), .B1(n_549), .B2(n_550), .C(n_553), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_534), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g573 ( .A(n_534), .B(n_563), .Y(n_573) );
AND2x2_ASAP7_75t_L g581 ( .A(n_534), .B(n_536), .Y(n_581) );
OR2x2_ASAP7_75t_L g593 ( .A(n_534), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_534), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g635 ( .A(n_534), .B(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_534), .Y(n_655) );
AND2x2_ASAP7_75t_L g707 ( .A(n_534), .B(n_631), .Y(n_707) );
OAI31xp33_ASAP7_75t_L g715 ( .A1(n_534), .A2(n_584), .A3(n_683), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_535), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g679 ( .A(n_535), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_535), .B(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g567 ( .A(n_536), .B(n_563), .Y(n_567) );
INVx1_ASAP7_75t_L g654 ( .A(n_536), .Y(n_654) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g704 ( .A(n_537), .B(n_563), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_SL g714 ( .A(n_547), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_548), .B(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_549), .A2(n_661), .B1(n_699), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g562 ( .A(n_552), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g621 ( .A(n_552), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_552), .B(n_573), .Y(n_726) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g696 ( .A(n_555), .B(n_697), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_556), .A2(n_615), .B(n_617), .Y(n_614) );
OR2x2_ASAP7_75t_L g622 ( .A(n_556), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g643 ( .A(n_556), .B(n_631), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_556), .B(n_654), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_556), .B(n_694), .Y(n_693) );
OAI221xp5_ASAP7_75t_SL g670 ( .A1(n_557), .A2(n_671), .B1(n_676), .B2(n_679), .C(n_680), .Y(n_670) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OR2x2_ASAP7_75t_L g647 ( .A(n_558), .B(n_620), .Y(n_647) );
INVx1_ASAP7_75t_L g686 ( .A(n_558), .Y(n_686) );
INVx2_ASAP7_75t_L g662 ( .A(n_559), .Y(n_662) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g601 ( .A(n_563), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_563), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_563), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g718 ( .A(n_563), .B(n_688), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B1(n_570), .B2(n_573), .C1(n_574), .C2(n_576), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g574 ( .A(n_567), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_567), .A2(n_617), .B1(n_645), .B2(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_567), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_576), .A2(n_606), .B(n_609), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_582), .B(n_583), .C(n_605), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_581), .A2(n_584), .B1(n_589), .B2(n_590), .C(n_592), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_581), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g675 ( .A(n_581), .Y(n_675) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
AND2x2_ASAP7_75t_L g677 ( .A(n_586), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g594 ( .A(n_589), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_589), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_599), .B2(n_602), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_596), .B(n_608), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_597), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g697 ( .A(n_601), .Y(n_697) );
AND2x2_ASAP7_75t_L g716 ( .A(n_601), .B(n_631), .Y(n_716) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_608), .B(n_665), .Y(n_724) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_611), .B(n_679), .Y(n_722) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g645 ( .A(n_623), .Y(n_645) );
BUFx2_ASAP7_75t_L g669 ( .A(n_624), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_628), .B(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_648), .C(n_670), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_652), .B(n_656), .C(n_659), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_649), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp67_ASAP7_75t_SL g653 ( .A(n_654), .B(n_655), .Y(n_653) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_SL g678 ( .A(n_658), .Y(n_678) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_667), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g683 ( .A(n_661), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_685), .B2(n_687), .Y(n_680) );
INVx2_ASAP7_75t_SL g701 ( .A(n_688), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_705), .C(n_717), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_701), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B1(n_712), .B2(n_714), .C(n_715), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_706), .A2(n_718), .B(n_719), .C(n_721), .Y(n_717) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_725), .B2(n_727), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g737 ( .A(n_729), .Y(n_737) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g757 ( .A(n_745), .Y(n_757) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g761 ( .A(n_749), .Y(n_761) );
INVx1_ASAP7_75t_L g754 ( .A(n_751), .Y(n_754) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule