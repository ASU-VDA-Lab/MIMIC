module fake_jpeg_22076_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp67_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_35),
.B(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_1),
.Y(n_53)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_32),
.B1(n_28),
.B2(n_22),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_51),
.B(n_2),
.Y(n_107)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_17),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_21),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_68),
.B(n_55),
.C(n_34),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_22),
.B1(n_28),
.B2(n_32),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_74),
.B1(n_23),
.B2(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_29),
.B1(n_19),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_18),
.B1(n_60),
.B2(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_34),
.B1(n_24),
.B2(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_33),
.C(n_20),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_23),
.Y(n_94)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_48),
.B1(n_18),
.B2(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_72),
.B1(n_61),
.B2(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_17),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_99),
.Y(n_136)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_23),
.B1(n_34),
.B2(n_17),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_74),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_43),
.CI(n_34),
.CON(n_108),
.SN(n_108)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_74),
.B(n_66),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_113),
.B(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_115),
.B1(n_87),
.B2(n_89),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_137),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_80),
.B(n_66),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_131),
.C(n_139),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_108),
.B1(n_109),
.B2(n_54),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_88),
.B1(n_83),
.B2(n_5),
.Y(n_157)
);

XNOR2x2_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_50),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_81),
.B1(n_52),
.B2(n_65),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_128),
.B1(n_111),
.B2(n_87),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_77),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_132),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_134),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_81),
.B(n_43),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_56),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_56),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_17),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_17),
.B(n_4),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_153),
.Y(n_179)
);

OR2x2_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_154),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_89),
.B1(n_90),
.B2(n_96),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_158),
.B1(n_147),
.B2(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_162),
.C(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_163),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_3),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_88),
.B1(n_83),
.B2(n_7),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_114),
.B1(n_119),
.B2(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_14),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_181),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_182),
.B(n_153),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_112),
.B(n_113),
.C(n_138),
.D(n_125),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_142),
.B(n_159),
.C(n_163),
.D(n_117),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_125),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_116),
.B1(n_128),
.B2(n_117),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_142),
.C(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_120),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

OAI321xp33_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_163),
.A3(n_182),
.B1(n_180),
.B2(n_178),
.C(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_197),
.C(n_198),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_157),
.B1(n_160),
.B2(n_175),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_165),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_148),
.B1(n_159),
.B2(n_127),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_195),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_139),
.B(n_129),
.C(n_121),
.D(n_120),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_176),
.C(n_181),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_210),
.B(n_8),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_168),
.B1(n_177),
.B2(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_190),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_172),
.C(n_171),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.C(n_188),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_172),
.C(n_134),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_200),
.B1(n_201),
.B2(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_197),
.C(n_189),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_186),
.B(n_4),
.C(n_7),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_9),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_127),
.C(n_8),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_3),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_9),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_226),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_221),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_219),
.B(n_220),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_218),
.B1(n_207),
.B2(n_202),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_9),
.C(n_10),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_215),
.C(n_217),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_231),
.A2(n_232),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_234),
.C(n_11),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_223),
.B(n_10),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_238),
.B(n_14),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_11),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_11),
.B(n_13),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.Y(n_244)
);


endmodule