module real_jpeg_11736_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_37),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_18),
.B(n_20),
.C(n_24),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_9),
.B(n_31),
.C(n_53),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_9),
.A2(n_68),
.B(n_70),
.Y(n_98)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_72),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_71),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_61),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_61),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_38),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_26),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_18),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g43 ( 
.A1(n_18),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_43)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_21),
.B(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_27),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_22),
.A2(n_23),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_23),
.B(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_34),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_27),
.A2(n_34),
.B(n_89),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_28),
.B(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_28),
.A2(n_35),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_30),
.A2(n_31),
.B1(n_53),
.B2(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_30),
.B(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_45),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_55),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_64),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.C(n_67),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_85),
.B(n_103),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_82),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_93),
.B(n_102),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_91),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_101),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);


endmodule