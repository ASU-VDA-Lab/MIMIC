module real_jpeg_14988_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_28),
.B1(n_46),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_51),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_28),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_23),
.B1(n_28),
.B2(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_23),
.B1(n_56),
.B2(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_10),
.B(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_54),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_10),
.B(n_35),
.C(n_83),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_10),
.B(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_84),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_24),
.B(n_59),
.C(n_175),
.Y(n_174)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_116),
.B1(n_196),
.B2(n_197),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_14),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_114),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_101),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_16),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_68),
.B2(n_69),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_20),
.A2(n_21),
.B1(n_30),
.B2(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.C(n_26),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_23),
.A2(n_56),
.B(n_60),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_24),
.A2(n_25),
.B1(n_59),
.B2(n_60),
.Y(n_67)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B(n_37),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_32),
.B(n_128),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_32),
.A2(n_40),
.B(n_110),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_33),
.A2(n_40),
.B(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AO22x1_ASAP7_75t_L g84 ( 
.A1(n_34),
.A2(n_35),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_35),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_37),
.B(n_159),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_40),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_40),
.B(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_62),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_57),
.B(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_61),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_92),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.C(n_87),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_78),
.B1(n_87),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_80),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_80),
.B(n_100),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_84),
.B(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_84),
.B(n_98),
.Y(n_182)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_95),
.B(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_107),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_102),
.A2(n_103),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_106),
.B(n_107),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_107),
.A2(n_180),
.B1(n_186),
.B2(n_187),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_111),
.CI(n_112),
.CON(n_107),
.SN(n_107)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_109),
.B(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_190),
.B(n_195),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_178),
.B(n_189),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_162),
.B(n_177),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_144),
.B(n_161),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_138),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_129),
.B1(n_130),
.B2(n_137),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_135),
.C(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_155),
.B(n_160),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_151),
.B(n_154),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_158),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_164),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);


endmodule