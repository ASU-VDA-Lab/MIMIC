module fake_jpeg_378_n_72 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_67;
wire n_66;

INVx1_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_22),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_26),
.B(n_22),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_28),
.B(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_38),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_1),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_43),
.B(n_45),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_58),
.C(n_2),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_44),
.C(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_12),
.Y(n_55)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_47),
.B(n_48),
.C(n_4),
.D(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_60),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_47),
.B(n_13),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_19),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_61),
.B(n_4),
.C(n_6),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_65),
.A3(n_66),
.B1(n_23),
.B2(n_8),
.C1(n_9),
.C2(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_65),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_16),
.A3(n_15),
.B1(n_14),
.B2(n_8),
.Y(n_70)
);

A2O1A1O1Ixp25_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_3),
.B(n_6),
.C(n_7),
.D(n_9),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_23),
.Y(n_72)
);


endmodule