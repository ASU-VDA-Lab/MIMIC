module real_jpeg_25693_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_47),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_2),
.B(n_66),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_2),
.B(n_49),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_2),
.B(n_33),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_27),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_5),
.B(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_5),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_33),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_5),
.B(n_52),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_5),
.B(n_49),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_47),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_5),
.B(n_66),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_6),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_6),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_6),
.B(n_33),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_6),
.B(n_52),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_8),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_33),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_8),
.B(n_52),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_8),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_8),
.B(n_49),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_8),
.B(n_47),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_8),
.B(n_66),
.Y(n_288)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_10),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_10),
.B(n_17),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_10),
.B(n_33),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_10),
.B(n_52),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_11),
.B(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_11),
.B(n_47),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_52),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_11),
.B(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_11),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_11),
.B(n_66),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_27),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_11),
.B(n_43),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_12),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_12),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_12),
.B(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_66),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_27),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_13),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_13),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_13),
.B(n_52),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_15),
.B(n_47),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_16),
.B(n_52),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_16),
.B(n_49),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_16),
.B(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_16),
.B(n_17),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_16),
.B(n_47),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_16),
.B(n_66),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_16),
.B(n_27),
.Y(n_282)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_17),
.Y(n_163)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_17),
.Y(n_209)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_17),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_94),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_21),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_70),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_22),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_23),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_60),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_SL g92 ( 
.A(n_30),
.B(n_83),
.C(n_93),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_30),
.A2(n_38),
.B1(n_82),
.B2(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_32),
.B(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_36),
.Y(n_172)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_39),
.B(n_45),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_40),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_41),
.A2(n_42),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_43),
.Y(n_265)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_45),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_52),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_54),
.B(n_70),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_55),
.A2(n_56),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_62),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_57),
.B(n_59),
.CI(n_62),
.CON(n_310),
.SN(n_310)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_61),
.B(n_63),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_73),
.C(n_75),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_65),
.A2(n_69),
.B1(n_74),
.B2(n_339),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_69),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_76),
.A2(n_77),
.B1(n_94),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_88),
.C(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_80),
.B(n_83),
.C(n_84),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_85),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_99),
.SN(n_99)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_94),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_101),
.C(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_96),
.B(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_98),
.B(n_99),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_99),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_108),
.C(n_111),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_117),
.Y(n_358)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.CI(n_120),
.CON(n_117),
.SN(n_117)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_350),
.C(n_351),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_342),
.C(n_343),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_327),
.C(n_328),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_305),
.C(n_306),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_271),
.C(n_272),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_239),
.C(n_240),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_214),
.C(n_215),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_174),
.C(n_186),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_158),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_153),
.C(n_158),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_148),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_159),
.B(n_167),
.C(n_168),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_173),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_185),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_179),
.B1(n_185),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_210),
.C(n_211),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.C(n_200),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_193),
.C(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.C(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_228),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_229),
.C(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_223),
.C(n_224),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_222),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_224),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.CI(n_227),
.CON(n_224),
.SN(n_224)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_226),
.C(n_227),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_238),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_236),
.B2(n_237),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_232),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.C(n_237),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_255),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_244),
.C(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_251),
.C(n_254),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g360 ( 
.A(n_246),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.CI(n_249),
.CON(n_246),
.SN(n_246)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_248),
.C(n_249),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_263),
.C(n_269),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_263),
.B1(n_269),
.B2(n_270),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_261),
.B(n_262),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_295),
.C(n_296),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_263),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_291),
.B2(n_304),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_292),
.C(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_277),
.C(n_284),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_284),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_280),
.C(n_283),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_289),
.C(n_290),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_297),
.B(n_323),
.C(n_324),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.CI(n_303),
.CON(n_297),
.SN(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_325),
.B2(n_326),
.Y(n_306)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_317),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_317),
.C(n_325),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_310),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_320),
.C(n_321),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_331),
.C(n_341),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_341),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_334),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_334),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.CI(n_337),
.CON(n_334),
.SN(n_334)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_336),
.C(n_337),
.Y(n_349)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_347),
.C(n_349),
.Y(n_350)
);


endmodule