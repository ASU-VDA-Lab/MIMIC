module fake_netlist_1_6786_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
NAND2xp33_ASAP7_75t_R g12 ( .A(n_7), .B(n_10), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
BUFx10_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_17), .B(n_2), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_13), .B(n_2), .C(n_4), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_11), .A2(n_6), .B(n_8), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_14), .B(n_5), .Y(n_22) );
A2O1A1Ixp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_19), .B(n_18), .C(n_21), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_18), .B(n_15), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_16), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_24), .B(n_11), .Y(n_27) );
AOI21xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_23), .B(n_12), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx2_ASAP7_75t_SL g30 ( .A(n_29), .Y(n_30) );
AOI322xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_5), .A3(n_9), .B1(n_16), .B2(n_26), .C1(n_27), .C2(n_29), .Y(n_31) );
CKINVDCx16_ASAP7_75t_R g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
BUFx2_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
OAI21xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_26), .B(n_27), .Y(n_35) );
OAI22xp5_ASAP7_75t_SL g36 ( .A1(n_32), .A2(n_27), .B1(n_26), .B2(n_16), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_27), .B1(n_34), .B2(n_35), .Y(n_37) );
endmodule