module real_jpeg_21026_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_240;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx13_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_52),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_35),
.B1(n_43),
.B2(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_3),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_112),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_112),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_3),
.A2(n_43),
.B1(n_51),
.B2(n_112),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_4),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_43),
.B1(n_51),
.B2(n_147),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_147),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_6),
.A2(n_103),
.B(n_154),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_8),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_141),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_141),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_43),
.B1(n_51),
.B2(n_141),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_9),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_14),
.B(n_47),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_9),
.A2(n_43),
.B1(n_51),
.B2(n_145),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_79),
.B1(n_202),
.B2(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_9),
.B(n_27),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_27),
.B(n_229),
.Y(n_233)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_43),
.B1(n_51),
.B2(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_63),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_13),
.A2(n_32),
.B1(n_43),
.B2(n_51),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_13),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_43),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_92),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_92),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_19),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_66),
.CI(n_75),
.CON(n_19),
.SN(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_33),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_23),
.A2(n_88),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_23),
.B(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_23),
.A2(n_88),
.B1(n_111),
.B2(n_160),
.Y(n_273)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_25),
.B(n_30),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_24),
.B(n_90),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_24),
.A2(n_36),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_25),
.B(n_27),
.Y(n_151)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_26),
.A2(n_37),
.B1(n_144),
.B2(n_151),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g228 ( 
.A1(n_26),
.A2(n_43),
.A3(n_58),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_27),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_30),
.B(n_145),
.CON(n_144),
.SN(n_144)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_53),
.B2(n_54),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_49),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_42),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_42),
.A2(n_45),
.B1(n_84),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_42),
.A2(n_49),
.B(n_85),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_42),
.A2(n_45),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_42),
.A2(n_45),
.B1(n_198),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_42),
.A2(n_45),
.B1(n_220),
.B2(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_42),
.A2(n_70),
.B(n_236),
.Y(n_251)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_45),
.A2(n_72),
.B(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_45),
.B(n_145),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_46),
.B(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_80),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_48),
.A2(n_51),
.B(n_145),
.C(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_71),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_51),
.B(n_57),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_55),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_55),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_55),
.A2(n_64),
.B(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_56),
.A2(n_60),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_56),
.A2(n_60),
.B1(n_140),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_56),
.A2(n_60),
.B1(n_174),
.B2(n_233),
.Y(n_232)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_60),
.A2(n_68),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_60),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_60),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_65),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_86),
.B(n_87),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_77),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_86),
.B1(n_87),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_78),
.A2(n_83),
.B1(n_86),
.B2(n_290),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_79),
.A2(n_130),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_79),
.A2(n_188),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_79),
.A2(n_105),
.B(n_190),
.Y(n_221)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_80),
.B(n_145),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_82),
.A2(n_132),
.B(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_83),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_91),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_111),
.B(n_113),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_98),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_93),
.B(n_97),
.Y(n_297)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_98),
.A2(n_99),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.C(n_114),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_100),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_101),
.B(n_107),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_106),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_293),
.B(n_298),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_281),
.B(n_292),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_178),
.B(n_260),
.C(n_280),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_167),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_124),
.B(n_167),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_148),
.B2(n_166),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_127),
.B(n_135),
.C(n_166),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_128),
.B(n_134),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_143),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_149),
.B(n_157),
.C(n_162),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_168),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_176),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_173),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_175),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_259),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_253),
.B(n_258),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_241),
.B(n_252),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_223),
.B(n_240),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_211),
.B(n_222),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_199),
.B(n_210),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_191),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_205),
.B(n_209),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_219),
.C(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_225),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_231),
.B1(n_238),
.B2(n_239),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_243),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_250),
.C(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_262),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_278),
.B2(n_279),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.C(n_279),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_277),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_275),
.C(n_277),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_289),
.C(n_291),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);


endmodule