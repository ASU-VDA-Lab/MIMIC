module real_aes_597_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g207 ( .A(n_0), .B(n_154), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_2), .B(n_138), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_3), .B(n_156), .Y(n_547) );
INVx1_ASAP7_75t_L g145 ( .A(n_4), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_5), .B(n_138), .Y(n_137) );
NAND2xp33_ASAP7_75t_SL g251 ( .A(n_6), .B(n_144), .Y(n_251) );
INVx1_ASAP7_75t_L g243 ( .A(n_7), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_8), .Y(n_109) );
AND2x2_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g485 ( .A(n_10), .B(n_249), .Y(n_485) );
AND2x2_ASAP7_75t_L g549 ( .A(n_11), .B(n_183), .Y(n_549) );
INVx2_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_13), .B(n_156), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_14), .Y(n_111) );
AOI221x1_ASAP7_75t_L g246 ( .A1(n_15), .A2(n_147), .B1(n_247), .B2(n_249), .C(n_250), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_16), .B(n_138), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_17), .B(n_138), .Y(n_504) );
INVx1_ASAP7_75t_L g113 ( .A(n_18), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_19), .A2(n_64), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_19), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_20), .A2(n_91), .B1(n_138), .B2(n_187), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_21), .A2(n_147), .B(n_152), .Y(n_146) );
AOI221xp5_ASAP7_75t_SL g217 ( .A1(n_22), .A2(n_35), .B1(n_138), .B2(n_147), .C(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_23), .B(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g135 ( .A(n_24), .B(n_90), .Y(n_135) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_24), .A2(n_90), .B(n_134), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_25), .B(n_156), .Y(n_234) );
INVxp67_ASAP7_75t_L g245 ( .A(n_26), .Y(n_245) );
AND2x2_ASAP7_75t_L g178 ( .A(n_27), .B(n_168), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_28), .A2(n_147), .B(n_206), .Y(n_205) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_29), .A2(n_249), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_30), .B(n_156), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_31), .A2(n_147), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_32), .B(n_156), .Y(n_520) );
AND2x2_ASAP7_75t_L g144 ( .A(n_33), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g148 ( .A(n_33), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g195 ( .A(n_33), .Y(n_195) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_34), .B(n_108), .C(n_110), .Y(n_107) );
OR2x6_ASAP7_75t_L g120 ( .A(n_34), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_36), .B(n_138), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_37), .A2(n_82), .B1(n_147), .B2(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_38), .B(n_156), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_39), .B(n_138), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_40), .B(n_154), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_41), .A2(n_147), .B(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_42), .A2(n_50), .B1(n_774), .B2(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_42), .Y(n_775) );
AND2x2_ASAP7_75t_L g210 ( .A(n_43), .B(n_168), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_44), .B(n_154), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_45), .B(n_168), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_46), .B(n_138), .Y(n_528) );
INVx1_ASAP7_75t_L g141 ( .A(n_47), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_47), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_48), .A2(n_125), .B1(n_445), .B2(n_446), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_48), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_49), .B(n_156), .Y(n_483) );
INVx1_ASAP7_75t_L g774 ( .A(n_50), .Y(n_774) );
AND2x2_ASAP7_75t_L g495 ( .A(n_51), .B(n_168), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_52), .B(n_138), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_53), .B(n_154), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_54), .B(n_154), .Y(n_519) );
AND2x2_ASAP7_75t_L g169 ( .A(n_55), .B(n_168), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_56), .B(n_138), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_57), .B(n_156), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_58), .B(n_138), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_59), .A2(n_147), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_60), .B(n_154), .Y(n_165) );
AND2x2_ASAP7_75t_SL g235 ( .A(n_61), .B(n_133), .Y(n_235) );
AND2x2_ASAP7_75t_L g510 ( .A(n_62), .B(n_133), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_63), .A2(n_147), .B(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_64), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_65), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_66), .B(n_183), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_67), .B(n_154), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_68), .B(n_154), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_69), .A2(n_93), .B1(n_147), .B2(n_193), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_70), .B(n_156), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_71), .Y(n_785) );
INVx1_ASAP7_75t_L g143 ( .A(n_72), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_72), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_73), .B(n_154), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_74), .A2(n_147), .B(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_75), .A2(n_147), .B(n_473), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_76), .A2(n_147), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g522 ( .A(n_77), .B(n_133), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_78), .B(n_168), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_79), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_79), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_80), .B(n_138), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_81), .A2(n_84), .B1(n_138), .B2(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_83), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_85), .B(n_154), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_86), .B(n_154), .Y(n_220) );
AND2x2_ASAP7_75t_L g476 ( .A(n_87), .B(n_183), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_88), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_89), .A2(n_147), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_92), .B(n_156), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_94), .A2(n_147), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_95), .B(n_156), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_96), .B(n_138), .Y(n_209) );
INVxp67_ASAP7_75t_L g248 ( .A(n_97), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_98), .B(n_156), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_99), .A2(n_147), .B(n_232), .Y(n_231) );
BUFx2_ASAP7_75t_L g509 ( .A(n_100), .Y(n_509) );
BUFx2_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_102), .A2(n_770), .B1(n_777), .B2(n_780), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_114), .B(n_784), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
BUFx4f_ASAP7_75t_SL g787 ( .A(n_106), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_107), .B(n_112), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_111), .B(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_SL g460 ( .A(n_111), .B(n_120), .Y(n_460) );
OR2x6_ASAP7_75t_SL g769 ( .A(n_111), .B(n_119), .Y(n_769) );
OR2x2_ASAP7_75t_L g783 ( .A(n_111), .B(n_120), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_113), .B(n_122), .Y(n_121) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_452), .Y(n_114) );
AO21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_124), .B(n_447), .Y(n_115) );
NOR2x1_ASAP7_75t_R g116 ( .A(n_117), .B(n_123), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx3_ASAP7_75t_L g451 ( .A(n_118), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_123), .Y(n_454) );
INVx2_ASAP7_75t_L g445 ( .A(n_125), .Y(n_445) );
XNOR2x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_442), .Y(n_125) );
INVx3_ASAP7_75t_SL g458 ( .A(n_126), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g777 ( .A1(n_126), .A2(n_462), .B1(n_778), .B2(n_779), .Y(n_777) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_372), .Y(n_126) );
NOR4xp25_ASAP7_75t_SL g127 ( .A(n_128), .B(n_265), .C(n_309), .D(n_336), .Y(n_127) );
OAI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_226), .B1(n_236), .B2(n_253), .C(n_255), .Y(n_128) );
AOI32xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_179), .A3(n_199), .B1(n_211), .B2(n_222), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_130), .B(n_408), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_130), .A2(n_378), .B1(n_436), .B2(n_439), .Y(n_435) );
AND2x4_ASAP7_75t_SL g130 ( .A(n_131), .B(n_159), .Y(n_130) );
INVx5_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
OR2x2_ASAP7_75t_L g254 ( .A(n_131), .B(n_224), .Y(n_254) );
AND2x4_ASAP7_75t_L g256 ( .A(n_131), .B(n_171), .Y(n_256) );
INVx2_ASAP7_75t_L g271 ( .A(n_131), .Y(n_271) );
OR2x2_ASAP7_75t_L g283 ( .A(n_131), .B(n_180), .Y(n_283) );
AND2x2_ASAP7_75t_L g290 ( .A(n_131), .B(n_170), .Y(n_290) );
AND2x2_ASAP7_75t_SL g332 ( .A(n_131), .B(n_213), .Y(n_332) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_131), .Y(n_389) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g158 ( .A(n_134), .B(n_135), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_158), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g252 ( .A(n_139), .Y(n_252) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x6_ASAP7_75t_L g154 ( .A(n_140), .B(n_149), .Y(n_154) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g156 ( .A(n_142), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
AND2x2_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
INVx2_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
AND2x4_ASAP7_75t_L g193 ( .A(n_150), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_154), .B(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_157), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_157), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_157), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_157), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_157), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_157), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_157), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_157), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_157), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_157), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_157), .A2(n_546), .B(n_547), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_158), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_158), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_158), .B(n_248), .Y(n_247) );
NOR3xp33_ASAP7_75t_L g250 ( .A(n_158), .B(n_251), .C(n_252), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_158), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_158), .A2(n_528), .B(n_529), .Y(n_527) );
INVx3_ASAP7_75t_SL g284 ( .A(n_159), .Y(n_284) );
AND2x2_ASAP7_75t_L g303 ( .A(n_159), .B(n_225), .Y(n_303) );
AOI32xp33_ASAP7_75t_L g418 ( .A1(n_159), .A2(n_289), .A3(n_319), .B1(n_349), .B2(n_384), .Y(n_418) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_170), .Y(n_159) );
AND2x2_ASAP7_75t_L g258 ( .A(n_160), .B(n_180), .Y(n_258) );
OR2x2_ASAP7_75t_L g274 ( .A(n_160), .B(n_171), .Y(n_274) );
INVx1_ASAP7_75t_L g297 ( .A(n_160), .Y(n_297) );
INVx2_ASAP7_75t_L g313 ( .A(n_160), .Y(n_313) );
AND2x2_ASAP7_75t_L g350 ( .A(n_160), .B(n_213), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_160), .B(n_171), .Y(n_369) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_160), .Y(n_438) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_167), .B(n_169), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_167), .A2(n_172), .B(n_178), .Y(n_171) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_167), .A2(n_172), .B(n_178), .Y(n_224) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_167), .A2(n_543), .B(n_549), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_168), .A2(n_217), .B(n_221), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_168), .A2(n_471), .B(n_472), .Y(n_470) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_168), .A2(n_489), .B(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g405 ( .A(n_171), .B(n_180), .Y(n_405) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_171), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_177), .Y(n_172) );
OR2x2_ASAP7_75t_L g253 ( .A(n_179), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g259 ( .A(n_179), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g272 ( .A(n_179), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g434 ( .A(n_179), .B(n_303), .Y(n_434) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g363 ( .A(n_180), .B(n_313), .Y(n_363) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_181), .Y(n_213) );
AOI21x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_185), .B(n_198), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_183), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_183), .A2(n_504), .B(n_505), .Y(n_503) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx3_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_192), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_187), .A2(n_193), .B1(n_242), .B2(n_244), .Y(n_241) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_191), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2x1p5_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_199), .B(n_330), .Y(n_432) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_200), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g215 ( .A(n_201), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g237 ( .A(n_201), .Y(n_237) );
AND2x2_ASAP7_75t_L g263 ( .A(n_201), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_201), .B(n_239), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_201), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g321 ( .A(n_201), .Y(n_321) );
OR2x2_ASAP7_75t_L g340 ( .A(n_201), .B(n_267), .Y(n_340) );
INVx1_ASAP7_75t_L g347 ( .A(n_201), .Y(n_347) );
NOR2xp33_ASAP7_75t_R g399 ( .A(n_201), .B(n_228), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_201), .B(n_240), .Y(n_403) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21x1_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_210), .Y(n_202) );
INVx4_ASAP7_75t_L g249 ( .A(n_203), .Y(n_249) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_203), .A2(n_479), .B(n_485), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_211), .A2(n_262), .A3(n_427), .B1(n_428), .B2(n_429), .Y(n_426) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx2_ASAP7_75t_L g293 ( .A(n_213), .Y(n_293) );
AND2x4_ASAP7_75t_L g312 ( .A(n_213), .B(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_213), .B(n_284), .Y(n_341) );
OR2x2_ASAP7_75t_L g395 ( .A(n_213), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g353 ( .A(n_214), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g411 ( .A(n_214), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_215), .B(n_228), .Y(n_377) );
AND2x2_ASAP7_75t_L g414 ( .A(n_215), .B(n_380), .Y(n_414) );
INVx2_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
INVx2_ASAP7_75t_L g267 ( .A(n_216), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_216), .B(n_228), .Y(n_287) );
INVx1_ASAP7_75t_L g318 ( .A(n_216), .Y(n_318) );
OR2x2_ASAP7_75t_L g344 ( .A(n_216), .B(n_228), .Y(n_344) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_216), .Y(n_396) );
BUFx3_ASAP7_75t_L g425 ( .A(n_216), .Y(n_425) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g294 ( .A(n_223), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_223), .B(n_312), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_223), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_224), .B(n_297), .Y(n_296) );
OAI21xp33_ASAP7_75t_L g326 ( .A1(n_224), .A2(n_293), .B(n_311), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g348 ( .A1(n_225), .A2(n_349), .A3(n_351), .B1(n_353), .B2(n_355), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_225), .B(n_312), .Y(n_421) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g354 ( .A(n_227), .Y(n_354) );
NOR2x1p5_ASAP7_75t_L g424 ( .A(n_227), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g238 ( .A(n_228), .B(n_239), .Y(n_238) );
AND2x4_ASAP7_75t_SL g262 ( .A(n_228), .B(n_240), .Y(n_262) );
OR2x2_ASAP7_75t_L g266 ( .A(n_228), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g301 ( .A(n_228), .Y(n_301) );
AND2x2_ASAP7_75t_L g319 ( .A(n_228), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g330 ( .A(n_228), .B(n_240), .Y(n_330) );
OR2x2_ASAP7_75t_L g392 ( .A(n_228), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g409 ( .A(n_228), .B(n_340), .Y(n_409) );
INVx1_ASAP7_75t_L g441 ( .A(n_228), .Y(n_441) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_237), .B(n_318), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_238), .B(n_352), .Y(n_351) );
AOI222xp33_ASAP7_75t_L g356 ( .A1(n_238), .A2(n_357), .B1(n_362), .B2(n_364), .C1(n_367), .C2(n_370), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_238), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_238), .B(n_263), .Y(n_384) );
AND2x2_ASAP7_75t_L g346 ( .A(n_239), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g361 ( .A(n_239), .B(n_266), .Y(n_361) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_240), .B(n_267), .Y(n_299) );
AND2x4_ASAP7_75t_L g320 ( .A(n_240), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g380 ( .A(n_240), .B(n_301), .Y(n_380) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_246), .Y(n_240) );
INVx3_ASAP7_75t_L g515 ( .A(n_249), .Y(n_515) );
INVx1_ASAP7_75t_SL g260 ( .A(n_254), .Y(n_260) );
NAND2xp33_ASAP7_75t_SL g429 ( .A(n_254), .B(n_284), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_259), .C(n_261), .Y(n_255) );
INVx2_ASAP7_75t_SL g306 ( .A(n_256), .Y(n_306) );
AND2x2_ASAP7_75t_L g310 ( .A(n_257), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_258), .B(n_306), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_258), .A2(n_296), .B(n_332), .C(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g408 ( .A(n_258), .B(n_389), .Y(n_408) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x4_ASAP7_75t_L g307 ( .A(n_262), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g412 ( .A(n_262), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .B(n_275), .C(n_302), .Y(n_265) );
INVx2_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
OR2x2_ASAP7_75t_L g324 ( .A(n_266), .B(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_267), .Y(n_308) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_270), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g362 ( .A(n_270), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_270), .B(n_350), .Y(n_416) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_272), .A2(n_375), .B1(n_376), .B2(n_378), .C1(n_381), .C2(n_384), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_273), .A2(n_338), .B1(n_341), .B2(n_342), .C(n_348), .Y(n_337) );
AND2x2_ASAP7_75t_L g375 ( .A(n_273), .B(n_332), .Y(n_375) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp33_ASAP7_75t_SL g288 ( .A(n_274), .B(n_289), .Y(n_288) );
AOI221x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B1(n_285), .B2(n_288), .C(n_291), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g428 ( .A(n_278), .B(n_366), .Y(n_428) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g286 ( .A(n_279), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OAI32xp33_ASAP7_75t_L g394 ( .A1(n_284), .A2(n_325), .A3(n_395), .B1(n_397), .B2(n_401), .Y(n_394) );
OAI21xp33_ASAP7_75t_SL g413 ( .A1(n_285), .A2(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI21xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B(n_298), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g295 ( .A(n_293), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g368 ( .A(n_293), .B(n_369), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_297), .A2(n_323), .B1(n_326), .B2(n_327), .C(n_331), .Y(n_322) );
INVx1_ASAP7_75t_L g398 ( .A(n_297), .Y(n_398) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_297), .Y(n_404) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OAI21xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_306), .B(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_314), .B(n_322), .Y(n_309) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_316), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g335 ( .A(n_318), .Y(n_335) );
INVx1_ASAP7_75t_L g325 ( .A(n_320), .Y(n_325) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_320), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_320), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_320), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_335), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_337), .B(n_356), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g352 ( .A(n_340), .Y(n_352) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_SL g366 ( .A(n_344), .Y(n_366) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_346), .B(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_347), .Y(n_360) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_358), .B(n_361), .Y(n_357) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g371 ( .A(n_363), .Y(n_371) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g390 ( .A(n_369), .Y(n_390) );
NOR4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_406), .C(n_417), .D(n_430), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_385), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_375), .A2(n_386), .B(n_391), .C(n_394), .Y(n_385) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_390), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g397 ( .A1(n_388), .A2(n_398), .B(n_399), .C(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
OAI21xp33_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_404), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_405), .B(n_437), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_409), .B1(n_410), .B2(n_411), .C(n_413), .Y(n_406) );
INVx1_ASAP7_75t_SL g410 ( .A(n_408), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_419), .C(n_426), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp33_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
CKINVDCx11_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_770), .B(n_776), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI22x1_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_459), .B1(n_461), .B2(n_767), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
CKINVDCx11_ASAP7_75t_R g778 ( .A(n_460), .Y(n_778) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_692), .Y(n_462) );
NOR2xp67_ASAP7_75t_L g463 ( .A(n_464), .B(n_611), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_555), .C(n_565), .D(n_582), .E(n_598), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_491), .B1(n_533), .B2(n_537), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g539 ( .A(n_469), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g557 ( .A(n_469), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g578 ( .A(n_469), .B(n_579), .Y(n_578) );
INVx4_ASAP7_75t_L g592 ( .A(n_469), .Y(n_592) );
AND2x2_ASAP7_75t_L g601 ( .A(n_469), .B(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_SL g623 ( .A(n_469), .B(n_541), .Y(n_623) );
BUFx2_ASAP7_75t_L g666 ( .A(n_469), .Y(n_666) );
AND2x2_ASAP7_75t_L g681 ( .A(n_469), .B(n_478), .Y(n_681) );
OR2x2_ASAP7_75t_L g713 ( .A(n_469), .B(n_714), .Y(n_713) );
NOR4xp25_ASAP7_75t_L g762 ( .A(n_469), .B(n_763), .C(n_764), .D(n_765), .Y(n_762) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
AOI31xp33_ASAP7_75t_L g630 ( .A1(n_477), .A2(n_631), .A3(n_633), .B(n_635), .Y(n_630) );
INVx2_ASAP7_75t_SL g747 ( .A(n_477), .Y(n_747) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
INVx2_ASAP7_75t_L g554 ( .A(n_478), .Y(n_554) );
AND2x2_ASAP7_75t_L g558 ( .A(n_478), .B(n_542), .Y(n_558) );
INVx2_ASAP7_75t_L g581 ( .A(n_478), .Y(n_581) );
AND2x2_ASAP7_75t_L g600 ( .A(n_478), .B(n_541), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_484), .Y(n_479) );
AND2x2_ASAP7_75t_L g552 ( .A(n_486), .B(n_553), .Y(n_552) );
BUFx3_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
INVx2_ASAP7_75t_L g577 ( .A(n_486), .Y(n_577) );
AND2x2_ASAP7_75t_L g632 ( .A(n_486), .B(n_592), .Y(n_632) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
AND2x4_ASAP7_75t_L g603 ( .A(n_487), .B(n_488), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_523), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_511), .Y(n_492) );
OR2x2_ASAP7_75t_L g533 ( .A(n_493), .B(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g684 ( .A(n_493), .Y(n_684) );
OR2x2_ASAP7_75t_L g732 ( .A(n_493), .B(n_733), .Y(n_732) );
NAND2x1_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
OR2x2_ASAP7_75t_SL g524 ( .A(n_494), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g562 ( .A(n_494), .Y(n_562) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_494), .Y(n_606) );
INVx2_ASAP7_75t_L g614 ( .A(n_494), .Y(n_614) );
OR2x2_ASAP7_75t_L g649 ( .A(n_494), .B(n_513), .Y(n_649) );
AND2x2_ASAP7_75t_L g761 ( .A(n_494), .B(n_616), .Y(n_761) );
AND2x2_ASAP7_75t_L g766 ( .A(n_494), .B(n_526), .Y(n_766) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
OR2x2_ASAP7_75t_L g525 ( .A(n_502), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g590 ( .A(n_502), .B(n_512), .Y(n_590) );
OR2x2_ASAP7_75t_L g597 ( .A(n_502), .B(n_562), .Y(n_597) );
NOR2x1_ASAP7_75t_SL g616 ( .A(n_502), .B(n_536), .Y(n_616) );
BUFx2_ASAP7_75t_L g648 ( .A(n_502), .Y(n_648) );
AND2x2_ASAP7_75t_L g657 ( .A(n_502), .B(n_562), .Y(n_657) );
AND2x2_ASAP7_75t_L g690 ( .A(n_502), .B(n_610), .Y(n_690) );
INVx2_ASAP7_75t_SL g699 ( .A(n_502), .Y(n_699) );
AND2x2_ASAP7_75t_L g702 ( .A(n_502), .B(n_513), .Y(n_702) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_511), .B(n_567), .C(n_652), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_511), .B(n_614), .Y(n_717) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_512), .B(n_699), .Y(n_720) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_513), .Y(n_564) );
AND2x2_ASAP7_75t_L g608 ( .A(n_513), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g673 ( .A(n_513), .B(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_522), .Y(n_514) );
AO21x1_ASAP7_75t_SL g536 ( .A1(n_515), .A2(n_516), .B(n_522), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
AND2x4_ASAP7_75t_L g568 ( .A(n_523), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g704 ( .A(n_525), .B(n_649), .Y(n_704) );
AND2x2_ASAP7_75t_L g535 ( .A(n_526), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_526), .Y(n_589) );
INVx2_ASAP7_75t_L g610 ( .A(n_526), .Y(n_610) );
INVx1_ASAP7_75t_L g674 ( .A(n_526), .Y(n_674) );
INVx2_ASAP7_75t_L g756 ( .A(n_533), .Y(n_756) );
OR2x2_ASAP7_75t_L g620 ( .A(n_534), .B(n_597), .Y(n_620) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g760 ( .A(n_535), .B(n_657), .Y(n_760) );
AND2x2_ASAP7_75t_L g653 ( .A(n_536), .B(n_610), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_550), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_539), .A2(n_667), .B1(n_684), .B2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g580 ( .A(n_541), .Y(n_580) );
AND2x2_ASAP7_75t_L g634 ( .A(n_541), .B(n_554), .Y(n_634) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_541), .Y(n_661) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_542), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_552), .B(n_666), .Y(n_665) );
OAI32xp33_ASAP7_75t_L g682 ( .A1(n_552), .A2(n_683), .A3(n_685), .B1(n_686), .B2(n_688), .Y(n_682) );
BUFx2_ASAP7_75t_L g567 ( .A(n_553), .Y(n_567) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g709 ( .A(n_554), .B(n_603), .Y(n_709) );
OR4x1_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .C(n_560), .D(n_563), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_556), .A2(n_647), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_557), .Y(n_749) );
AND2x2_ASAP7_75t_L g591 ( .A(n_558), .B(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g671 ( .A(n_558), .Y(n_671) );
INVx1_ASAP7_75t_L g687 ( .A(n_558), .Y(n_687) );
INVx1_ASAP7_75t_L g722 ( .A(n_558), .Y(n_722) );
OR2x2_ASAP7_75t_L g679 ( .A(n_559), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g723 ( .A(n_559), .B(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_560), .A2(n_597), .B1(n_641), .B2(n_660), .Y(n_662) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g706 ( .A(n_561), .B(n_615), .Y(n_706) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g573 ( .A(n_562), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g588 ( .A(n_562), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g569 ( .A(n_563), .Y(n_569) );
NAND4xp25_ASAP7_75t_L g696 ( .A(n_563), .B(n_567), .C(n_648), .D(n_660), .Y(n_696) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g733 ( .A(n_564), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B1(n_570), .B2(n_574), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_566), .A2(n_567), .B1(n_717), .B2(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx3_ASAP7_75t_L g595 ( .A(n_572), .Y(n_595) );
AOI32xp33_ASAP7_75t_L g711 ( .A1(n_572), .A2(n_712), .A3(n_716), .B1(n_721), .B2(n_725), .Y(n_711) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_575), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g670 ( .A(n_575), .B(n_671), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_575), .A2(n_583), .B1(n_695), .B2(n_700), .C(n_703), .Y(n_694) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g627 ( .A(n_576), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g742 ( .A(n_576), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_577), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g584 ( .A(n_579), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_579), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_SL g642 ( .A(n_580), .Y(n_642) );
INVx1_ASAP7_75t_L g626 ( .A(n_581), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B1(n_591), .B2(n_593), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g728 ( .A(n_584), .B(n_658), .Y(n_728) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g668 ( .A(n_587), .Y(n_668) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_592), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_592), .B(n_629), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g641 ( .A(n_592), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_592), .B(n_634), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_593), .A2(n_753), .B1(n_754), .B2(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OR2x2_ASAP7_75t_L g635 ( .A(n_595), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g645 ( .A(n_595), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_595), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_595), .B(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_SL g700 ( .A(n_595), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g676 ( .A(n_597), .B(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g618 ( .A(n_600), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_601), .A2(n_638), .B1(n_645), .B2(n_650), .Y(n_637) );
INVx3_ASAP7_75t_L g640 ( .A(n_603), .Y(n_640) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI32xp33_ASAP7_75t_SL g695 ( .A1(n_606), .A2(n_666), .A3(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g615 ( .A(n_609), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g611 ( .A(n_612), .B(n_637), .C(n_654), .D(n_669), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_617), .B1(n_619), .B2(n_621), .C(n_630), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx2_ASAP7_75t_L g652 ( .A(n_614), .Y(n_652) );
AND2x2_ASAP7_75t_L g701 ( .A(n_614), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_614), .B(n_653), .Y(n_739) );
AND2x2_ASAP7_75t_L g750 ( .A(n_614), .B(n_673), .Y(n_750) );
INVx2_ASAP7_75t_L g636 ( .A(n_616), .Y(n_636) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B(n_627), .Y(n_621) );
AND2x2_ASAP7_75t_L g753 ( .A(n_622), .B(n_624), .Y(n_753) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_623), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g730 ( .A(n_628), .Y(n_730) );
INVx1_ASAP7_75t_L g715 ( .A(n_629), .Y(n_715) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_632), .B(n_687), .Y(n_686) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_633), .B(n_640), .Y(n_644) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g743 ( .A(n_634), .Y(n_743) );
INVx1_ASAP7_75t_L g725 ( .A(n_636), .Y(n_725) );
OR2x2_ASAP7_75t_L g741 ( .A(n_636), .B(n_652), .Y(n_741) );
NAND2xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_643), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g658 ( .A(n_640), .Y(n_658) );
AND2x2_ASAP7_75t_L g663 ( .A(n_640), .B(n_653), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_640), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g737 ( .A(n_641), .Y(n_737) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_646), .A2(n_727), .B1(n_729), .B2(n_731), .Y(n_726) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g691 ( .A(n_649), .Y(n_691) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g677 ( .A(n_653), .Y(n_677) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .A3(n_659), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_667), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g705 ( .A1(n_655), .A2(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_657), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g729 ( .A(n_658), .B(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_665), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g685 ( .A(n_666), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_666), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B1(n_675), .B2(n_678), .C(n_682), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_671), .A2(n_758), .B1(n_760), .B2(n_761), .C(n_762), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_673), .B(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g724 ( .A(n_674), .Y(n_724) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_678), .A2(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp33_ASAP7_75t_SL g758 ( .A(n_687), .B(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
NOR4xp75_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .C(n_734), .D(n_751), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_705), .Y(n_693) );
INVx1_ASAP7_75t_L g764 ( .A(n_702), .Y(n_764) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g736 ( .A(n_709), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g763 ( .A(n_709), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_726), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g759 ( .A(n_730), .Y(n_759) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND3x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_744), .C(n_748), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B(n_740), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_757), .Y(n_751) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g779 ( .A(n_768), .Y(n_779) );
CKINVDCx11_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
endmodule