module fake_jpeg_30940_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_48),
.B1(n_51),
.B2(n_55),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_77),
.C(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_45),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_45),
.B1(n_44),
.B2(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_47),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_3),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_52),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_92),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_90),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_89),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_40),
.B1(n_22),
.B2(n_24),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_0),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_19),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_3),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_1),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_69),
.C(n_26),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_17),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_79),
.B1(n_89),
.B2(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_108),
.B1(n_10),
.B2(n_15),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_7),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_32),
.B(n_13),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_117),
.B(n_33),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_34),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_105),
.C(n_102),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_10),
.B(n_16),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_100),
.B1(n_106),
.B2(n_93),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_31),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_129),
.B(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_130),
.A2(n_122),
.B1(n_116),
.B2(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_132),
.B1(n_116),
.B2(n_128),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.C(n_127),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_125),
.B(n_118),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_35),
.C(n_36),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_37),
.Y(n_138)
);


endmodule