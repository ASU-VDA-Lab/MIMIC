module real_jpeg_12118_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_314, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_314;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_59),
.B1(n_64),
.B2(n_98),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_98),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_39),
.B1(n_59),
.B2(n_64),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_7),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_253)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_9),
.A2(n_54),
.B1(n_59),
.B2(n_64),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_10),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_59),
.B1(n_64),
.B2(n_139),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_139),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_139),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_12),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_12),
.A2(n_44),
.B1(n_59),
.B2(n_64),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_13),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_13),
.B(n_59),
.C(n_63),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_49),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_13),
.A2(n_142),
.B(n_145),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_33),
.B(n_48),
.C(n_173),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_13),
.B(n_25),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_59),
.B1(n_64),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_14),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_144),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_144),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_144),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_59),
.B1(n_64),
.B2(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_16),
.A2(n_29),
.B1(n_59),
.B2(n_64),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_16),
.A2(n_29),
.B1(n_50),
.B2(n_51),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_16),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_112),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_20),
.B(n_99),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_80),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_21),
.B(n_72),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_71),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_22),
.A2(n_23),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_23),
.B(n_41),
.C(n_56),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_24),
.A2(n_31),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_26),
.B1(n_32),
.B2(n_36),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_26),
.A2(n_30),
.B(n_127),
.C(n_218),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_26),
.A2(n_33),
.A3(n_36),
.B1(n_219),
.B2(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_30),
.A2(n_31),
.B1(n_38),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_30),
.A2(n_31),
.B1(n_246),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_30),
.A2(n_266),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_31),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_31),
.B(n_97),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_31),
.A2(n_94),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_32),
.B(n_34),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_52),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_45),
.B(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_47),
.A2(n_50),
.B(n_127),
.Y(n_173)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_49),
.B(n_180),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_51),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_74),
.B1(n_76),
.B2(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_56),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_65),
.B(n_67),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_65),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_57),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_57),
.A2(n_65),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_57),
.A2(n_65),
.B1(n_225),
.B2(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_57),
.A2(n_65),
.B1(n_91),
.B2(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_68),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_138),
.B(n_140),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_58),
.B(n_127),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_58),
.A2(n_140),
.B(n_224),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_64),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_65),
.B(n_129),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_72),
.A2(n_73),
.B(n_77),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_74),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_74),
.A2(n_76),
.B1(n_193),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_74),
.A2(n_179),
.B(n_222),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_268),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_76),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_76),
.A2(n_194),
.B(n_268),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_126),
.B(n_128),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_78),
.A2(n_128),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_80),
.B(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_93),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_81),
.A2(n_82),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_83),
.A2(n_84),
.B1(n_93),
.B2(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_85),
.A2(n_86),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_85),
.B(n_146),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_85),
.A2(n_86),
.B1(n_236),
.B2(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_86),
.B(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_86),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_88),
.A2(n_142),
.B1(n_159),
.B2(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_93),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_308),
.B(n_312),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_295),
.B(n_307),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_278),
.B(n_294),
.Y(n_116)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_238),
.A3(n_271),
.B1(n_276),
.B2(n_277),
.C(n_314),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_210),
.B(n_237),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_187),
.B(n_209),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_168),
.B(n_186),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_147),
.B(n_167),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_159),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_130),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_137),
.C(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_142),
.A2(n_159),
.B1(n_175),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_142),
.A2(n_159),
.B1(n_201),
.B2(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_155),
.B(n_166),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_153),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_161),
.B(n_165),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_158),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_160),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_181),
.C(n_185),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_174),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_202),
.B2(n_203),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_205),
.C(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_196),
.C(n_200),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_212),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_228),
.C(n_229),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_220),
.B2(n_226),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_221),
.C(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_255),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_249),
.C(n_254),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_240),
.A2(n_241),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_247),
.C(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_254),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_252),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_263),
.C(n_270),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_261),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_293),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_293),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_289),
.C(n_292),
.Y(n_306)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_306),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.C(n_306),
.Y(n_311)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_311),
.Y(n_312)
);


endmodule