module fake_jpeg_12094_n_203 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_9),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_89),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_71),
.Y(n_87)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_94),
.Y(n_102)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_78),
.B1(n_82),
.B2(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_77),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_73),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_0),
.C(n_4),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_59),
.B1(n_69),
.B2(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_109),
.B1(n_82),
.B2(n_60),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_59),
.B1(n_91),
.B2(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_63),
.Y(n_121)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_80),
.B(n_75),
.C(n_58),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_72),
.B1(n_83),
.B2(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_120),
.B1(n_126),
.B2(n_130),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_82),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_67),
.C(n_62),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_6),
.C(n_7),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_72),
.B1(n_83),
.B2(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_4),
.Y(n_133)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_81),
.B1(n_60),
.B2(n_68),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_66),
.B1(n_1),
.B2(n_2),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_28),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_138),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_6),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_113),
.B(n_8),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_8),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_29),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_10),
.C(n_11),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_10),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_22),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_150),
.B1(n_149),
.B2(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_166),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_13),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_162),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_14),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_167),
.B(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_141),
.B1(n_41),
.B2(n_43),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_23),
.B(n_24),
.C(n_25),
.D(n_26),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_30),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_34),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_35),
.B(n_37),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_135),
.B(n_149),
.Y(n_173)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_40),
.C(n_46),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_183),
.C(n_169),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_49),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_160),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_182),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_163),
.A3(n_164),
.B1(n_158),
.B2(n_162),
.C1(n_56),
.C2(n_54),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_192),
.A2(n_193),
.B1(n_187),
.B2(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_178),
.C(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_186),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_194),
.B(n_192),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_176),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_174),
.Y(n_203)
);


endmodule