module fake_netlist_5_1840_n_296 (n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_48, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_296);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_296;

wire n_137;
wire n_210;
wire n_168;
wire n_294;
wire n_260;
wire n_164;
wire n_286;
wire n_91;
wire n_208;
wire n_82;
wire n_122;
wire n_194;
wire n_282;
wire n_142;
wire n_176;
wire n_214;
wire n_140;
wire n_248;
wire n_124;
wire n_86;
wire n_146;
wire n_136;
wire n_268;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_237;
wire n_90;
wire n_241;
wire n_127;
wire n_101;
wire n_75;
wire n_180;
wire n_184;
wire n_226;
wire n_235;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_281;
wire n_207;
wire n_240;
wire n_114;
wire n_57;
wire n_96;
wire n_189;
wire n_220;
wire n_291;
wire n_165;
wire n_111;
wire n_231;
wire n_108;
wire n_229;
wire n_257;
wire n_213;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_197;
wire n_107;
wire n_58;
wire n_69;
wire n_236;
wire n_116;
wire n_195;
wire n_227;
wire n_117;
wire n_249;
wire n_271;
wire n_284;
wire n_233;
wire n_94;
wire n_203;
wire n_245;
wire n_274;
wire n_205;
wire n_123;
wire n_113;
wire n_139;
wire n_105;
wire n_280;
wire n_246;
wire n_80;
wire n_179;
wire n_125;
wire n_269;
wire n_167;
wire n_128;
wire n_73;
wire n_234;
wire n_277;
wire n_92;
wire n_267;
wire n_149;
wire n_120;
wire n_285;
wire n_232;
wire n_135;
wire n_156;
wire n_126;
wire n_254;
wire n_225;
wire n_84;
wire n_202;
wire n_130;
wire n_266;
wire n_272;
wire n_219;
wire n_157;
wire n_258;
wire n_265;
wire n_79;
wire n_193;
wire n_293;
wire n_131;
wire n_151;
wire n_173;
wire n_192;
wire n_244;
wire n_251;
wire n_53;
wire n_160;
wire n_198;
wire n_223;
wire n_288;
wire n_247;
wire n_188;
wire n_190;
wire n_201;
wire n_292;
wire n_158;
wire n_263;
wire n_224;
wire n_100;
wire n_154;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_228;
wire n_264;
wire n_283;
wire n_109;
wire n_112;
wire n_212;
wire n_85;
wire n_159;
wire n_163;
wire n_276;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_243;
wire n_239;
wire n_275;
wire n_175;
wire n_252;
wire n_169;
wire n_59;
wire n_262;
wire n_255;
wire n_133;
wire n_238;
wire n_215;
wire n_295;
wire n_55;
wire n_196;
wire n_99;
wire n_211;
wire n_218;
wire n_181;
wire n_49;
wire n_290;
wire n_54;
wire n_147;
wire n_221;
wire n_178;
wire n_67;
wire n_121;
wire n_242;
wire n_76;
wire n_200;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_161;
wire n_209;
wire n_259;
wire n_273;
wire n_287;
wire n_270;
wire n_222;
wire n_230;
wire n_81;
wire n_118;
wire n_89;
wire n_279;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_253;
wire n_261;
wire n_72;
wire n_186;
wire n_174;
wire n_199;
wire n_289;
wire n_134;
wire n_187;
wire n_104;
wire n_191;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_141;
wire n_97;
wire n_166;
wire n_206;
wire n_217;
wire n_171;
wire n_153;
wire n_145;
wire n_256;
wire n_204;
wire n_50;
wire n_250;
wire n_52;
wire n_278;
wire n_88;
wire n_110;
wire n_216;

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_31),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_12),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_0),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_51),
.B(n_0),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NAND2x1p5_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_21),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_74),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_60),
.C(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_60),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_57),
.B1(n_74),
.B2(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_73),
.Y(n_113)
);

AND2x4_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_62),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_2),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_7),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_8),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_9),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_81),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

OR2x6_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_92),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_98),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_142),
.A2(n_129),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_110),
.B1(n_129),
.B2(n_124),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_125),
.B(n_99),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_84),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_84),
.Y(n_158)
);

AND2x4_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_146),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_97),
.B1(n_102),
.B2(n_100),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_84),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_103),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_91),
.B(n_90),
.C(n_103),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_155),
.B(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_146),
.B1(n_131),
.B2(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_156),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

AO21x2_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_131),
.B(n_130),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_130),
.B(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_157),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_130),
.B(n_133),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_159),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_184),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_183),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_142),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_142),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_197),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_191),
.B1(n_182),
.B2(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_173),
.B(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

OAI222xp33_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_136),
.B1(n_107),
.B2(n_161),
.C1(n_171),
.C2(n_182),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_170),
.B(n_187),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

AOI211xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_148),
.B(n_136),
.C(n_152),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_182),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_196),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_196),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

AO21x2_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_170),
.B(n_187),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_219),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_169),
.B1(n_168),
.B2(n_195),
.C(n_180),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_207),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

AND2x4_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_217),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_211),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_211),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_214),
.Y(n_244)
);

NOR2x1_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_217),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NAND2x1_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_214),
.B1(n_213),
.B2(n_176),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_229),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_169),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_202),
.Y(n_265)
);

AOI211xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_252),
.B(n_249),
.C(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_250),
.Y(n_267)
);

XOR2x2_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_245),
.Y(n_268)
);

NAND4xp25_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_240),
.C(n_199),
.D(n_177),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_10),
.Y(n_270)
);

AOI211x1_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_255),
.B(n_259),
.C(n_265),
.Y(n_271)
);

OAI211xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_261),
.B(n_256),
.C(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_263),
.B(n_262),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_270),
.B(n_260),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_271),
.B1(n_176),
.B2(n_216),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NAND4xp25_ASAP7_75t_SL g282 ( 
.A(n_280),
.B(n_11),
.C(n_13),
.D(n_15),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_16),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_216),
.C(n_133),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_26),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

OAI22x1_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_291),
.B1(n_290),
.B2(n_286),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_178),
.B(n_34),
.Y(n_293)
);

NOR4xp25_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_28),
.C(n_41),
.D(n_43),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_294),
.B(n_293),
.Y(n_296)
);


endmodule