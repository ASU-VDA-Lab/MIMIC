module real_jpeg_25897_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_0),
.A2(n_40),
.B1(n_42),
.B2(n_60),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_0),
.A2(n_27),
.B1(n_34),
.B2(n_60),
.Y(n_223)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_2),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_62),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_2),
.B(n_40),
.C(n_84),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_2),
.A2(n_63),
.B1(n_68),
.B2(n_185),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_2),
.B(n_126),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_2),
.A2(n_40),
.B1(n_42),
.B2(n_185),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_2),
.B(n_27),
.C(n_45),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_2),
.A2(n_26),
.B(n_272),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_27),
.B1(n_34),
.B2(n_49),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_49),
.B1(n_63),
.B2(n_68),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_3),
.A2(n_49),
.B1(n_76),
.B2(n_77),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_76),
.B1(n_78),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_5),
.A2(n_63),
.B1(n_68),
.B2(n_161),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_161),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_5),
.A2(n_27),
.B1(n_34),
.B2(n_161),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_58),
.B1(n_78),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_8),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_63),
.B1(n_68),
.B2(n_111),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_111),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_8),
.A2(n_27),
.B1(n_34),
.B2(n_111),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_63),
.B1(n_68),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_11),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_88),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_11),
.A2(n_27),
.B1(n_34),
.B2(n_88),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_39),
.B1(n_63),
.B2(n_68),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_13),
.A2(n_39),
.B1(n_78),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_13),
.A2(n_27),
.B1(n_34),
.B2(n_39),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_14),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_14),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_35),
.B1(n_63),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_14),
.A2(n_35),
.B1(n_58),
.B2(n_77),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_15),
.A2(n_59),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_15),
.A2(n_63),
.B1(n_68),
.B2(n_73),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_15),
.A2(n_40),
.B1(n_42),
.B2(n_73),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_15),
.A2(n_27),
.B1(n_34),
.B2(n_73),
.Y(n_242)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_16),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_355),
.B(n_358),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_350),
.B(n_354),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_337),
.B(n_349),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_136),
.A3(n_151),
.B(n_334),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_115),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_22),
.B(n_115),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.C(n_95),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_23),
.A2(n_79),
.B1(n_80),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_23),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_51),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_24),
.A2(n_25),
.B(n_53),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_25),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_25),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_26),
.A2(n_33),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_100),
.B1(n_101),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_26),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_26),
.A2(n_101),
.B1(n_190),
.B2(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_26),
.B(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_26),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_29),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_31),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_34),
.B(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_38),
.A2(n_43),
.B1(n_50),
.B2(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_40),
.A2(n_42),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_40),
.B(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_43),
.A2(n_50),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_43),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_43),
.A2(n_50),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_47),
.A2(n_91),
.B1(n_105),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_171),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_47),
.A2(n_210),
.B(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_47),
.B(n_185),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_50),
.B(n_211),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_55),
.A2(n_61),
.B1(n_112),
.B2(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_57),
.B(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_59),
.A2(n_184),
.B(n_185),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_61),
.A2(n_112),
.B1(n_134),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_61),
.A2(n_69),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_62),
.A2(n_74),
.B1(n_110),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_62),
.A2(n_74),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_62),
.A2(n_74),
.B1(n_345),
.B2(n_352),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_62),
.A2(n_74),
.B(n_352),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_68),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_63),
.A2(n_67),
.B(n_184),
.C(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_63),
.B(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_67),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_SL g186 ( 
.A(n_66),
.B(n_68),
.C(n_78),
.Y(n_186)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_74),
.A2(n_114),
.B(n_213),
.Y(n_212)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_94),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_82),
.A2(n_83),
.B1(n_128),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_82),
.A2(n_178),
.B(n_180),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_82),
.A2(n_180),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_107),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_83),
.A2(n_164),
.B(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_89),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_91),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_91),
.A2(n_260),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_95),
.A2(n_96),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.C(n_108),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_97),
.A2(n_98),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_99),
.Y(n_173)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_101),
.Y(n_301)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_106),
.B(n_108),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_133),
.B2(n_135),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_126),
.B1(n_179),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_125),
.A2(n_126),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_126),
.B(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_130),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_130),
.B(n_143),
.C(n_148),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_135),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_133),
.B(n_139),
.C(n_142),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_137),
.A2(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_150),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_138),
.B(n_150),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_144),
.Y(n_344)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_149),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_327),
.B(n_333),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_199),
.B(n_326),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_192),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_154),
.B(n_192),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_172),
.C(n_174),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_155),
.A2(n_156),
.B1(n_172),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_166),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_162),
.C(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_170),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_172),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_174),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_181),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_177),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_181),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_185),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_188),
.A2(n_284),
.B1(n_286),
.B2(n_288),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_194),
.B(n_195),
.C(n_198),
.Y(n_332)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_230),
.B(n_320),
.C(n_325),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_224),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_214),
.C(n_217),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_202),
.A2(n_203),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.C(n_212),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_217),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_313),
.B(n_319),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_261),
.B(n_312),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_250),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_235),
.B(n_250),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_243),
.C(n_247),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_242),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_243),
.A2(n_247),
.B1(n_248),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_251),
.B(n_257),
.C(n_258),
.Y(n_318)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_306),
.B(n_311),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_281),
.B(n_305),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_275),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_275),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_291),
.B(n_304),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_289),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_297),
.B(n_303),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_318),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_332),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_339),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_343),
.B1(n_346),
.B2(n_347),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_341),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_343),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_346),
.C(n_348),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_353),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_356),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_351),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_360),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_359),
.Y(n_358)
);


endmodule