module real_jpeg_7747_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_1),
.A2(n_16),
.B(n_31),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_2),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_2),
.A2(n_22),
.B1(n_64),
.B2(n_67),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_2),
.A2(n_22),
.B1(n_46),
.B2(n_47),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_54),
.B1(n_64),
.B2(n_67),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_54),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_9),
.A2(n_33),
.B1(n_64),
.B2(n_67),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_10),
.A2(n_56),
.B1(n_64),
.B2(n_67),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_11),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_64),
.B1(n_67),
.B2(n_91),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_91),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_12),
.A2(n_64),
.B1(n_67),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_12),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_108),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_108),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_108),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_13),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_156),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_156),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_156),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_14),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_14),
.A2(n_64),
.B1(n_67),
.B2(n_103),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_103),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_103),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_16),
.A2(n_47),
.B(n_59),
.C(n_88),
.D(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_16),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_45),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_16),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_16),
.A2(n_109),
.B(n_112),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_16),
.A2(n_30),
.B(n_41),
.C(n_144),
.D(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_16),
.B(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_34),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_16),
.A2(n_23),
.B1(n_24),
.B2(n_125),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_77),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_75),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_35),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_32),
.B2(n_34),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_21),
.A2(n_25),
.B1(n_34),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_23),
.A2(n_27),
.B(n_125),
.C(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_25),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_25),
.B(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_26),
.A2(n_29),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_26),
.A2(n_29),
.B1(n_215),
.B2(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_26),
.A2(n_206),
.B(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_26),
.A2(n_29),
.B1(n_53),
.B2(n_288),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_29),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_29),
.A2(n_216),
.B(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_34),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_70),
.C(n_72),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_36),
.A2(n_37),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_51),
.C(n_57),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_38),
.A2(n_39),
.B1(n_57),
.B2(n_313),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_40),
.A2(n_49),
.B1(n_165),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_40),
.A2(n_201),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_45),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_41),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_41),
.A2(n_45),
.B1(n_241),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_41),
.A2(n_45),
.B1(n_260),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_42),
.B(n_47),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_44),
.A2(n_46),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_49),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_49),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_49),
.A2(n_166),
.B(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_51),
.A2(n_52),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_57),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_57),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_58),
.A2(n_68),
.B1(n_102),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_58),
.A2(n_142),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_58),
.A2(n_68),
.B1(n_198),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_58),
.A2(n_68),
.B1(n_226),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_58),
.A2(n_68),
.B1(n_235),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_59),
.A2(n_63),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_67),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_64),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_67),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_68),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_68),
.A2(n_104),
.B(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_69),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_70),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_331),
.B(n_337),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_304),
.A3(n_324),
.B1(n_329),
.B2(n_330),
.C(n_339),
.Y(n_78)
);

AOI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_252),
.A3(n_292),
.B1(n_298),
.B2(n_303),
.C(n_340),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_209),
.C(n_248),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_180),
.B(n_208),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_159),
.B(n_179),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_136),
.B(n_158),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_114),
.B(n_135),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_96),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_86),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_89),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_101),
.C(n_106),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B(n_112),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_109),
.A2(n_127),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_109),
.A2(n_127),
.B1(n_191),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_109),
.A2(n_127),
.B1(n_224),
.B2(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_109),
.A2(n_127),
.B(n_233),
.Y(n_265)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_111),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_113),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_111),
.B1(n_155),
.B2(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_122),
.B(n_134),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_120),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_129),
.B(n_133),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_126),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_127),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_128),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_138),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_157),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_148),
.C(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_153),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_175),
.C(n_177),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_172),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_169),
.C(n_170),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_195),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_194),
.C(n_195),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_210),
.A2(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_228),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_211),
.B(n_228),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.C(n_227),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_220),
.C(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_227),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_246),
.B2(n_247),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_236),
.C(n_247),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_242),
.C(n_245),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_250),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_270),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_253),
.B(n_270),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_263),
.C(n_269),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_254),
.A2(n_255),
.B1(n_263),
.B2(n_297),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_263),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_265),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_283),
.B(n_287),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_267),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_290),
.B2(n_291),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_281),
.B2(n_282),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_273),
.B(n_282),
.C(n_291),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_278),
.B(n_280),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_279),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_280),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_280),
.A2(n_306),
.B1(n_315),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_289),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_285),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_299),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_317),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_317),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_315),
.C(n_316),
.Y(n_305)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_308),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_313),
.C(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_319),
.C(n_323),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_311),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_336),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_336),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule