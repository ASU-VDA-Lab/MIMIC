module fake_netlist_1_1279_n_716 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_716);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx3_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_34), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_19), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_75), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_7), .Y(n_84) );
INVx1_ASAP7_75t_SL g85 ( .A(n_26), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_61), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_32), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_73), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_9), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_18), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_39), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_68), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_22), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_78), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_0), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_66), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_74), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_60), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_59), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_13), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_24), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_13), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_45), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_47), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_20), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_29), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_69), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_8), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_31), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_10), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_30), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_1), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_51), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_37), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_76), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_108), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_106), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVxp33_ASAP7_75t_SL g138 ( .A(n_116), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_116), .B(n_2), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_118), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_118), .B(n_4), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_121), .B(n_4), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_84), .B(n_5), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_109), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_107), .B(n_5), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_90), .B(n_6), .Y(n_153) );
OR2x2_ASAP7_75t_L g154 ( .A(n_99), .B(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_82), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_80), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_104), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_101), .Y(n_162) );
BUFx10_ASAP7_75t_L g163 ( .A(n_81), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_127), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_113), .B(n_7), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_83), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_86), .Y(n_168) );
INVx5_ASAP7_75t_L g169 ( .A(n_105), .Y(n_169) );
BUFx8_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_94), .B(n_9), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_152), .B(n_110), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_144), .B(n_120), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_129), .B(n_81), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_144), .B(n_100), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_131), .B(n_126), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_169), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_146), .B(n_123), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_163), .B(n_93), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_163), .B(n_93), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
AND2x6_ASAP7_75t_L g189 ( .A(n_153), .B(n_105), .Y(n_189) );
INVxp33_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_163), .B(n_124), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_138), .B(n_102), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_152), .B(n_111), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_154), .A2(n_125), .B1(n_124), .B2(n_89), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_161), .A2(n_122), .B1(n_119), .B2(n_96), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_131), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_131), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_130), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_158), .B(n_97), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_141), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_158), .B(n_98), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_133), .B(n_103), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_133), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_152), .B(n_112), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_152), .B(n_115), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_170), .Y(n_213) );
INVx5_ASAP7_75t_L g214 ( .A(n_157), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_166), .B(n_117), .Y(n_215) );
INVxp33_ASAP7_75t_SL g216 ( .A(n_128), .Y(n_216) );
INVx6_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
BUFx10_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
BUFx4f_ASAP7_75t_L g219 ( .A(n_134), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_148), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_132), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_170), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_168), .B(n_117), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_136), .B(n_114), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_134), .A2(n_100), .B1(n_95), .B2(n_89), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_135), .B(n_95), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_157), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_142), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_132), .Y(n_231) );
INVx5_ASAP7_75t_L g232 ( .A(n_157), .Y(n_232) );
NOR2xp33_ASAP7_75t_SL g233 ( .A(n_170), .B(n_85), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_135), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_169), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_169), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_218), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_218), .B(n_168), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_204), .Y(n_240) );
NAND3xp33_ASAP7_75t_SL g241 ( .A(n_220), .B(n_145), .C(n_154), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_220), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_215), .B(n_137), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_213), .B(n_165), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_190), .B(n_137), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_225), .B(n_143), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_190), .B(n_143), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_199), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_200), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g251 ( .A(n_183), .B(n_151), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_228), .B(n_151), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_203), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_234), .B(n_155), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_228), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_179), .B(n_155), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_228), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_222), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_207), .B(n_171), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_216), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_213), .B(n_149), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_226), .A2(n_164), .B1(n_139), .B2(n_167), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
INVx5_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_226), .B(n_139), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_224), .A2(n_160), .B(n_167), .Y(n_266) );
INVx8_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_214), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_207), .B(n_164), .Y(n_269) );
BUFx12f_ASAP7_75t_L g270 ( .A(n_226), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_208), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_222), .Y(n_272) );
OR2x6_ASAP7_75t_L g273 ( .A(n_226), .B(n_139), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_230), .A2(n_160), .B1(n_167), .B2(n_162), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_189), .A2(n_164), .B1(n_159), .B2(n_162), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_177), .B(n_139), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_175), .B(n_159), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_189), .A2(n_162), .B1(n_160), .B2(n_159), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_192), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_180), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_180), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_223), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_173), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_180), .Y(n_285) );
BUFx12f_ASAP7_75t_L g286 ( .A(n_211), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_176), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_189), .A2(n_169), .B1(n_156), .B2(n_150), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_196), .A2(n_156), .B1(n_150), .B2(n_12), .Y(n_289) );
NAND2xp33_ASAP7_75t_L g290 ( .A(n_223), .B(n_156), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_207), .B(n_156), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_219), .A2(n_156), .B(n_150), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_178), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_216), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_219), .B(n_156), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_233), .A2(n_150), .B1(n_11), .B2(n_15), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_189), .A2(n_150), .B1(n_11), .B2(n_15), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_188), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_219), .B(n_44), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_214), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_193), .B(n_46), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_173), .A2(n_41), .B(n_70), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_191), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_229), .Y(n_304) );
NOR2x1p5_ASAP7_75t_L g305 ( .A(n_211), .B(n_10), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_238), .A2(n_173), .B(n_182), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_262), .A2(n_182), .B(n_195), .C(n_194), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_246), .B(n_227), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_248), .B(n_186), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_281), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_258), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_251), .A2(n_182), .B1(n_195), .B2(n_187), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_256), .A2(n_195), .B(n_205), .C(n_202), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_247), .A2(n_209), .B(n_174), .C(n_194), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_189), .B1(n_210), .B2(n_209), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
AOI21x1_ASAP7_75t_L g321 ( .A1(n_245), .A2(n_174), .B(n_172), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
NOR2x1_ASAP7_75t_SL g323 ( .A(n_286), .B(n_232), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_293), .A2(n_303), .B1(n_298), .B2(n_271), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_253), .Y(n_325) );
AOI21x1_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_172), .B(n_184), .Y(n_326) );
NAND2x2_ASAP7_75t_L g327 ( .A(n_305), .B(n_197), .Y(n_327) );
BUFx8_ASAP7_75t_SL g328 ( .A(n_260), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_258), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_294), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_252), .A2(n_214), .B(n_232), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_241), .B(n_16), .Y(n_332) );
INVx8_ASAP7_75t_L g333 ( .A(n_267), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_253), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_280), .B(n_210), .Y(n_335) );
BUFx12f_ASAP7_75t_L g336 ( .A(n_243), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_257), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_278), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_259), .A2(n_214), .B1(n_232), .B2(n_210), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_272), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_244), .B(n_210), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_265), .Y(n_342) );
HB1xp67_ASAP7_75t_SL g343 ( .A(n_255), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_261), .A2(n_214), .B(n_232), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_272), .Y(n_346) );
OAI22xp5_ASAP7_75t_SL g347 ( .A1(n_270), .A2(n_232), .B1(n_17), .B2(n_16), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_237), .B(n_181), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_269), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_254), .A2(n_235), .B(n_236), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_265), .A2(n_210), .B1(n_217), .B2(n_236), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_275), .B(n_259), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_267), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_263), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_239), .B(n_210), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_267), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_277), .B(n_185), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_269), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_321), .A2(n_302), .B(n_299), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_338), .A2(n_254), .B1(n_276), .B2(n_279), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_328), .Y(n_363) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_347), .A2(n_266), .B1(n_304), .B2(n_242), .C1(n_249), .C2(n_250), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_327), .A2(n_265), .B1(n_273), .B2(n_274), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_312), .B(n_273), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_311), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_327), .A2(n_273), .B1(n_301), .B2(n_289), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_307), .A2(n_299), .B(n_266), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_264), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_306), .A2(n_295), .B(n_288), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_308), .B(n_264), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_324), .A2(n_291), .B(n_296), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_324), .A2(n_291), .B(n_297), .Y(n_374) );
INVxp67_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
AO32x2_ASAP7_75t_L g377 ( .A1(n_314), .A2(n_185), .A3(n_181), .B1(n_17), .B2(n_283), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_337), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_315), .A2(n_231), .B(n_201), .C(n_206), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_350), .A2(n_268), .B(n_300), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g381 ( .A1(n_315), .A2(n_221), .B(n_201), .C(n_206), .Y(n_381) );
OAI22x1_ASAP7_75t_L g382 ( .A1(n_332), .A2(n_264), .B1(n_23), .B2(n_25), .Y(n_382) );
OA21x2_ASAP7_75t_L g383 ( .A1(n_316), .A2(n_231), .B(n_221), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_310), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_344), .A2(n_184), .B(n_283), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_309), .A2(n_290), .B(n_283), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g387 ( .A(n_336), .B(n_264), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_333), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_328), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_352), .B(n_185), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_349), .A2(n_217), .B1(n_181), .B2(n_235), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_364), .B(n_358), .Y(n_392) );
AOI22xp5_ASAP7_75t_SL g393 ( .A1(n_363), .A2(n_343), .B1(n_335), .B2(n_354), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_384), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_378), .B(n_320), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_375), .A2(n_341), .B1(n_333), .B2(n_318), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_390), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_380), .A2(n_346), .B(n_344), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_316), .B(n_357), .C(n_317), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_372), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_365), .A2(n_335), .B1(n_319), .B2(n_322), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_366), .A2(n_317), .B1(n_357), .B2(n_351), .C(n_339), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_362), .A2(n_354), .B1(n_334), .B2(n_325), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_360), .A2(n_355), .B(n_348), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_382), .A2(n_331), .B1(n_345), .B2(n_348), .C(n_340), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_329), .B1(n_340), .B2(n_346), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_386), .A2(n_313), .B(n_311), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_379), .A2(n_313), .B(n_311), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_359), .B(n_323), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_370), .A2(n_329), .B1(n_313), .B2(n_311), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_388), .B(n_313), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_388), .A2(n_356), .B1(n_353), .B2(n_217), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_388), .A2(n_356), .B1(n_353), .B2(n_212), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_363), .A2(n_356), .B1(n_353), .B2(n_212), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_359), .B(n_356), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_367), .B(n_353), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_404), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_420), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_415), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_394), .B(n_377), .Y(n_424) );
AND2x4_ASAP7_75t_SL g425 ( .A(n_415), .B(n_367), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_404), .Y(n_426) );
INVx4_ASAP7_75t_L g427 ( .A(n_420), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_411), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_411), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_392), .A2(n_389), .B1(n_377), .B2(n_367), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_419), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_410), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_400), .Y(n_437) );
AOI21x1_ASAP7_75t_L g438 ( .A1(n_412), .A2(n_383), .B(n_380), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_410), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_397), .B(n_383), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_409), .B(n_373), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_420), .B(n_385), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_395), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_413), .B(n_373), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_419), .B(n_385), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_419), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
AO31x2_ASAP7_75t_L g450 ( .A1(n_399), .A2(n_381), .A3(n_379), .B(n_391), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_403), .B(n_377), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_408), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_401), .B(n_381), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_402), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_393), .B(n_369), .Y(n_456) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_455), .A2(n_389), .B1(n_396), .B2(n_387), .C1(n_393), .C2(n_407), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_428), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_428), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_455), .A2(n_406), .B1(n_418), .B2(n_414), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_428), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_429), .B(n_369), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_429), .B(n_374), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_442), .B(n_374), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_426), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_421), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_421), .Y(n_469) );
AO21x1_ASAP7_75t_L g470 ( .A1(n_430), .A2(n_452), .B(n_456), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_442), .B(n_361), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_442), .B(n_361), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_447), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_440), .B(n_445), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_424), .B(n_371), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_456), .B(n_371), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_425), .Y(n_479) );
AND2x4_ASAP7_75t_SL g480 ( .A(n_427), .B(n_417), .Y(n_480) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_430), .A2(n_416), .B(n_212), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_446), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_21), .Y(n_484) );
AOI21xp5_ASAP7_75t_SL g485 ( .A1(n_445), .A2(n_27), .B(n_28), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_431), .B(n_33), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_435), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_440), .B(n_35), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_455), .A2(n_212), .B1(n_38), .B2(n_40), .C(n_48), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_445), .B(n_437), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_423), .A2(n_36), .B1(n_49), .B2(n_50), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_436), .B(n_71), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_423), .B(n_52), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_423), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_454), .A2(n_55), .B1(n_56), .B2(n_57), .C(n_62), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_432), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_491), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_504), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_491), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_482), .B(n_443), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_465), .B(n_443), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_465), .B(n_456), .Y(n_513) );
NOR2xp67_ASAP7_75t_L g514 ( .A(n_506), .B(n_439), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_487), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_467), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_458), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_477), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_498), .B(n_448), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_498), .B(n_448), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_501), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_465), .B(n_456), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_495), .B(n_452), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_501), .B(n_427), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_477), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_505), .Y(n_527) );
AO21x1_ASAP7_75t_L g528 ( .A1(n_489), .A2(n_452), .B(n_427), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_505), .B(n_448), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_479), .B(n_427), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_495), .B(n_439), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_479), .B(n_451), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_474), .B(n_436), .Y(n_533) );
AOI211xp5_ASAP7_75t_L g534 ( .A1(n_470), .A2(n_434), .B(n_454), .C(n_451), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_467), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_459), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_475), .B(n_451), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_475), .B(n_451), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_466), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_474), .B(n_441), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_474), .B(n_441), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_493), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_476), .B(n_441), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_473), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_477), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_436), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_476), .B(n_449), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_457), .B(n_434), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_492), .B(n_444), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_482), .B(n_449), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_493), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_473), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_459), .B(n_422), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_473), .B(n_422), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_464), .B(n_422), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_464), .B(n_422), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_458), .B(n_450), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_471), .B(n_444), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_471), .B(n_444), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_458), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_461), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_471), .B(n_444), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_472), .B(n_492), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_461), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_461), .B(n_450), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_514), .B(n_470), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_564), .B(n_502), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_522), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_559), .B(n_502), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_508), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_508), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_550), .B(n_497), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_559), .B(n_497), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_524), .B(n_472), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_550), .B(n_478), .Y(n_576) );
AND2x4_ASAP7_75t_SL g577 ( .A(n_550), .B(n_487), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_524), .B(n_472), .Y(n_578) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_539), .B(n_487), .Y(n_579) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_545), .B(n_500), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_560), .B(n_478), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_546), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_560), .B(n_478), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_563), .B(n_478), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_564), .B(n_466), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_563), .B(n_463), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_518), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_516), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_543), .B(n_463), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_516), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_512), .B(n_463), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_535), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_552), .B(n_462), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_518), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_531), .B(n_462), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_549), .A2(n_457), .B1(n_481), .B2(n_460), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_509), .B(n_489), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_535), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_531), .B(n_462), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_510), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_526), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_525), .A2(n_481), .B1(n_506), .B2(n_484), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_511), .B(n_468), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_513), .B(n_500), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_512), .B(n_484), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_513), .B(n_484), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_548), .B(n_503), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_548), .B(n_503), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_521), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_561), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_511), .B(n_466), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_523), .B(n_503), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_527), .Y(n_613) );
NAND2xp33_ASAP7_75t_SL g614 ( .A(n_526), .B(n_481), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_523), .B(n_468), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_534), .A2(n_499), .B1(n_481), .B2(n_490), .C(n_485), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_544), .B(n_499), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_536), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_569), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_619), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_567), .A2(n_528), .B(n_530), .C(n_515), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_569), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_591), .B(n_544), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_600), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_567), .A2(n_528), .B(n_540), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_579), .A2(n_480), .B1(n_547), .B2(n_532), .Y(n_627) );
OAI22xp33_ASAP7_75t_SL g628 ( .A1(n_587), .A2(n_551), .B1(n_554), .B2(n_557), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_576), .B(n_533), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_579), .A2(n_557), .B1(n_556), .B2(n_554), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_614), .A2(n_496), .B(n_480), .Y(n_632) );
AOI21xp33_ASAP7_75t_SL g633 ( .A1(n_580), .A2(n_551), .B(n_556), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_597), .A2(n_537), .B1(n_538), .B2(n_536), .C(n_555), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_575), .B(n_547), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_580), .A2(n_529), .B1(n_519), .B2(n_520), .C1(n_553), .C2(n_541), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_581), .B(n_541), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_613), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_596), .A2(n_562), .B1(n_517), .B2(n_558), .Y(n_639) );
NOR4xp25_ASAP7_75t_L g640 ( .A(n_582), .B(n_542), .C(n_533), .D(n_566), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_578), .B(n_566), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_571), .Y(n_642) );
AOI221x1_ASAP7_75t_L g643 ( .A1(n_614), .A2(n_499), .B1(n_496), .B2(n_507), .C(n_517), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_572), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g646 ( .A1(n_601), .A2(n_480), .A3(n_558), .B(n_542), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_602), .A2(n_468), .B1(n_490), .B2(n_507), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g648 ( .A1(n_577), .A2(n_496), .A3(n_425), .B1(n_494), .B2(n_507), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_607), .B(n_488), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_608), .B(n_488), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_606), .A2(n_488), .B(n_486), .C(n_483), .Y(n_651) );
AOI221x1_ASAP7_75t_L g652 ( .A1(n_594), .A2(n_597), .B1(n_618), .B2(n_598), .C(n_592), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_594), .A2(n_486), .B(n_483), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_610), .B(n_486), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_616), .A2(n_483), .B1(n_425), .B2(n_432), .C1(n_450), .C2(n_438), .Y(n_655) );
OAI222xp33_ASAP7_75t_L g656 ( .A1(n_568), .A2(n_438), .B1(n_450), .B2(n_432), .C1(n_65), .C2(n_63), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_620), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_625), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_631), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_638), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_654), .Y(n_662) );
AOI211xp5_ASAP7_75t_SL g663 ( .A1(n_639), .A2(n_606), .B(n_604), .C(n_610), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_640), .B(n_577), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_629), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_642), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_621), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_634), .B(n_586), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_629), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_644), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_639), .A2(n_604), .B(n_573), .C(n_576), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_645), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_622), .A2(n_593), .B1(n_590), .B2(n_589), .C(n_603), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_636), .B(n_615), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_636), .B(n_599), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_655), .B(n_611), .C(n_617), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_633), .B(n_573), .Y(n_677) );
NOR2x1p5_ASAP7_75t_L g678 ( .A(n_641), .B(n_573), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_652), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_666), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_676), .B(n_635), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_670), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_672), .Y(n_683) );
NAND2xp33_ASAP7_75t_SL g684 ( .A(n_664), .B(n_630), .Y(n_684) );
NAND2xp33_ASAP7_75t_R g685 ( .A(n_664), .B(n_626), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_663), .A2(n_632), .B1(n_643), .B2(n_647), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_662), .Y(n_687) );
AOI221xp5_ASAP7_75t_SL g688 ( .A1(n_679), .A2(n_628), .B1(n_651), .B2(n_624), .C(n_637), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_677), .B(n_576), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_675), .A2(n_655), .B(n_627), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_679), .A2(n_646), .B(n_656), .C(n_653), .Y(n_691) );
OAI322xp33_ASAP7_75t_SL g692 ( .A1(n_674), .A2(n_595), .A3(n_649), .B1(n_650), .B2(n_648), .C1(n_605), .C2(n_574), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_671), .B(n_612), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_680), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_689), .B(n_678), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_684), .A2(n_673), .B1(n_668), .B2(n_667), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_688), .A2(n_669), .A3(n_665), .B1(n_667), .B2(n_661), .C1(n_660), .C2(n_659), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_681), .B(n_662), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_693), .A2(n_658), .B1(n_657), .B2(n_585), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_687), .Y(n_700) );
OAI31xp33_ASAP7_75t_L g701 ( .A1(n_686), .A2(n_570), .A3(n_583), .B(n_584), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_696), .B(n_690), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_697), .B(n_686), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_699), .A2(n_691), .B1(n_692), .B2(n_685), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_699), .A2(n_695), .B1(n_698), .B2(n_700), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_694), .Y(n_706) );
XNOR2x1_ASAP7_75t_L g707 ( .A(n_704), .B(n_701), .Y(n_707) );
XNOR2xp5_ASAP7_75t_L g708 ( .A(n_702), .B(n_682), .Y(n_708) );
OR3x1_ASAP7_75t_L g709 ( .A(n_703), .B(n_685), .C(n_683), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_707), .Y(n_710) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_709), .B(n_705), .Y(n_711) );
OAI22x1_ASAP7_75t_L g712 ( .A1(n_710), .A2(n_708), .B1(n_706), .B2(n_612), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_712), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_711), .B1(n_612), .B2(n_432), .Y(n_714) );
AO221x1_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_711), .B1(n_432), .B2(n_64), .C(n_450), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_432), .B1(n_450), .B2(n_710), .C(n_709), .Y(n_716) );
endmodule