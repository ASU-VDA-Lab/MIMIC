module fake_jpeg_26258_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_15),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_26),
.B1(n_39),
.B2(n_18),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_63),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_28),
.B1(n_19),
.B2(n_32),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_42),
.A3(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_18),
.B1(n_22),
.B2(n_31),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_22),
.B1(n_31),
.B2(n_28),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_73),
.B1(n_59),
.B2(n_58),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_19),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_91),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_56),
.B1(n_55),
.B2(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_89),
.B1(n_59),
.B2(n_75),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_44),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_18),
.B1(n_16),
.B2(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_20),
.B(n_16),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_111),
.B1(n_69),
.B2(n_27),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_54),
.B(n_1),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_97),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_55),
.C(n_58),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_104),
.B1(n_92),
.B2(n_117),
.Y(n_136)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_46),
.C(n_47),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_70),
.C(n_85),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_75),
.B1(n_65),
.B2(n_76),
.Y(n_125)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_126),
.B(n_30),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_81),
.B1(n_73),
.B2(n_47),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_129),
.B1(n_130),
.B2(n_135),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_86),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_134),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_112),
.B1(n_102),
.B2(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_131),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_115),
.B1(n_110),
.B2(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_67),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_20),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_67),
.B1(n_76),
.B2(n_69),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_109),
.B1(n_108),
.B2(n_113),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_31),
.B1(n_12),
.B2(n_14),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_99),
.C(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_32),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_148),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_158),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_157),
.B1(n_160),
.B2(n_0),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_98),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_153),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_99),
.A3(n_93),
.B1(n_96),
.B2(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_113),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_30),
.B1(n_29),
.B2(n_86),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_19),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_37),
.B1(n_32),
.B2(n_19),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_170),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_37),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_174),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_29),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_118),
.A2(n_37),
.A3(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_144),
.B(n_127),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_187),
.B(n_195),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_185),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_148),
.A2(n_122),
.B1(n_132),
.B2(n_127),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_188),
.B1(n_193),
.B2(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_123),
.C(n_133),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_13),
.C(n_11),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_133),
.B(n_142),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_143),
.B1(n_142),
.B2(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_191),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_164),
.A2(n_143),
.B1(n_140),
.B2(n_137),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_14),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_158),
.B1(n_146),
.B2(n_149),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_212),
.B1(n_182),
.B2(n_188),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_170),
.B1(n_163),
.B2(n_171),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_200),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_175),
.B1(n_155),
.B2(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_210),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_152),
.B1(n_155),
.B2(n_167),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_172),
.B(n_161),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_1),
.B(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_196),
.C(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_10),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_10),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_10),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_224),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_13),
.B1(n_9),
.B2(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_225),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_9),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_1),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_239),
.B1(n_242),
.B2(n_207),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_189),
.C(n_183),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_240),
.C(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_176),
.B1(n_201),
.B2(n_197),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_212),
.B1(n_204),
.B2(n_217),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_222),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_246),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_179),
.B1(n_181),
.B2(n_195),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_190),
.C(n_177),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_199),
.B(n_194),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_207),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_179),
.B(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_237),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_215),
.C(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_252),
.C(n_255),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_232),
.B1(n_229),
.B2(n_246),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_221),
.C(n_218),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_244),
.B1(n_236),
.B2(n_234),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_228),
.B(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_226),
.C(n_217),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_224),
.C(n_2),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_237),
.C(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_4),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_232),
.C(n_243),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_234),
.CI(n_233),
.CON(n_273),
.SN(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_4),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_6),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_250),
.B1(n_256),
.B2(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_247),
.B(n_5),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_273),
.C(n_269),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_282),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_7),
.B1(n_8),
.B2(n_265),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_274),
.C(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_291),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_265),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_264),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_284),
.B(n_281),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_298),
.B(n_290),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_290),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_287),
.B(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_300),
.B(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_294),
.C(n_297),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_283),
.B1(n_279),
.B2(n_276),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_307),
.A2(n_8),
.B(n_299),
.Y(n_308)
);


endmodule