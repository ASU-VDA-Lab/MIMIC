module fake_jpeg_4502_n_138 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx4_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_22),
.Y(n_34)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_8),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_33),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_31),
.B1(n_24),
.B2(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_22),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_10),
.B1(n_24),
.B2(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_40),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_21),
.B1(n_27),
.B2(n_22),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_21),
.B1(n_27),
.B2(n_22),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_49),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_35),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_28),
.B(n_44),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_59),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_68),
.B1(n_71),
.B2(n_21),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_72),
.C(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_40),
.B1(n_58),
.B2(n_39),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_45),
.B(n_50),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_51),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_45),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_51),
.B(n_55),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_52),
.A3(n_49),
.B1(n_36),
.B2(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_83),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_49),
.B(n_34),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_70),
.B1(n_19),
.B2(n_16),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_47),
.B(n_19),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.C(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_47),
.B1(n_10),
.B2(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_26),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_78),
.A3(n_77),
.B1(n_81),
.B2(n_82),
.C1(n_88),
.C2(n_79),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_96),
.C(n_92),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_11),
.C(n_20),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_82),
.C(n_86),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_59),
.B(n_53),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_94),
.B1(n_97),
.B2(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_101),
.B1(n_98),
.B2(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_20),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_114),
.B1(n_107),
.B2(n_103),
.Y(n_120)
);

NAND4xp25_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_101),
.C(n_59),
.D(n_53),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_116),
.B(n_117),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_109),
.C(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_20),
.B1(n_11),
.B2(n_2),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_104),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_9),
.B(n_8),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_11),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_0),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_122),
.B1(n_9),
.B2(n_7),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_102),
.A3(n_11),
.B1(n_9),
.B2(n_7),
.C(n_4),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_0),
.B(n_1),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.C(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_11),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_127),
.B(n_2),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_2),
.B(n_3),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_118),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_5),
.B(n_134),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_124),
.B(n_3),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_137),
.B(n_5),
.Y(n_138)
);


endmodule