module fake_netlist_1_4159_n_534 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_534);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_534;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g72 ( .A(n_50), .Y(n_72) );
INVx2_ASAP7_75t_L g73 ( .A(n_54), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_71), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_65), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_7), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_53), .Y(n_77) );
BUFx3_ASAP7_75t_L g78 ( .A(n_21), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_47), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_20), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_32), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_51), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_13), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_30), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_6), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_9), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_10), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_48), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_13), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_63), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_68), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_42), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_45), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_55), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_1), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_70), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_69), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_11), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_23), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_59), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_17), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_66), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_78), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_83), .B(n_0), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_78), .B(n_0), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_76), .B(n_1), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_72), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_79), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_84), .B(n_2), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_82), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_72), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_86), .B(n_2), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_115), .B(n_85), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_125), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_115), .A2(n_106), .B1(n_95), .B2(n_104), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_112), .B(n_86), .Y(n_134) );
INVx2_ASAP7_75t_SL g135 ( .A(n_111), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_125), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx2_ASAP7_75t_SL g138 ( .A(n_111), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_110), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_111), .B(n_89), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_125), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_111), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_114), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_109), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
INVx1_ASAP7_75t_SL g146 ( .A(n_110), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_112), .B(n_95), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_118), .B(n_73), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_118), .B(n_73), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_111), .B(n_89), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_120), .A2(n_102), .B1(n_106), .B2(n_104), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_130), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_139), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_140), .B(n_117), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
BUFx4f_ASAP7_75t_L g161 ( .A(n_140), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_139), .B(n_117), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_140), .B(n_120), .Y(n_163) );
BUFx8_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_140), .A2(n_130), .B1(n_110), .B2(n_113), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_140), .B(n_121), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_146), .B(n_121), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_140), .A2(n_130), .B1(n_113), .B2(n_128), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_140), .B(n_122), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_140), .B(n_122), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
INVxp67_ASAP7_75t_SL g175 ( .A(n_142), .Y(n_175) );
NOR2xp67_ASAP7_75t_L g176 ( .A(n_142), .B(n_108), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_134), .B(n_130), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_146), .B(n_123), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_151), .B(n_123), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_142), .B(n_130), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_151), .B(n_128), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_134), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_177), .A2(n_151), .B1(n_142), .B2(n_135), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_174), .Y(n_190) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_174), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_177), .A2(n_151), .B1(n_135), .B2(n_138), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_167), .A2(n_155), .B(n_138), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_183), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_177), .A2(n_151), .B1(n_135), .B2(n_138), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_170), .A2(n_155), .B1(n_133), .B2(n_152), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_183), .Y(n_199) );
INVxp67_ASAP7_75t_SL g200 ( .A(n_164), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_183), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_164), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_170), .A2(n_155), .B1(n_133), .B2(n_152), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
INVx1_ASAP7_75t_SL g205 ( .A(n_188), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_177), .B(n_134), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_166), .A2(n_151), .B1(n_131), .B2(n_147), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_169), .B(n_147), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_181), .A2(n_151), .B1(n_131), .B2(n_147), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_174), .Y(n_211) );
BUFx16f_ASAP7_75t_R g212 ( .A(n_164), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_162), .A2(n_151), .B1(n_150), .B2(n_145), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_156), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_167), .A2(n_144), .B(n_153), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_157), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_160), .Y(n_218) );
BUFx2_ASAP7_75t_R g219 ( .A(n_159), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_159), .A2(n_80), .B1(n_90), .B2(n_148), .Y(n_220) );
OR2x2_ASAP7_75t_L g221 ( .A(n_187), .B(n_148), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_208), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_205), .B(n_163), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_206), .B(n_160), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_202), .B(n_161), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_197), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_206), .A2(n_164), .B1(n_161), .B2(n_187), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_208), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_219), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_210), .A2(n_176), .B(n_150), .C(n_184), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_206), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_202), .B(n_174), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_221), .Y(n_233) );
OAI221xp5_ASAP7_75t_L g234 ( .A1(n_209), .A2(n_186), .B1(n_172), .B2(n_184), .C(n_163), .Y(n_234) );
CKINVDCx14_ASAP7_75t_R g235 ( .A(n_212), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_211), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_220), .A2(n_161), .B1(n_173), .B2(n_172), .Y(n_237) );
NAND2x1_ASAP7_75t_L g238 ( .A(n_204), .B(n_157), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_196), .A2(n_161), .B1(n_173), .B2(n_168), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_203), .A2(n_176), .B1(n_113), .B2(n_186), .Y(n_242) );
AOI22xp33_ASAP7_75t_SL g243 ( .A1(n_218), .A2(n_87), .B1(n_185), .B2(n_174), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_215), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_168), .B1(n_175), .B2(n_174), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_218), .Y(n_246) );
OAI221xp5_ASAP7_75t_L g247 ( .A1(n_207), .A2(n_186), .B1(n_88), .B2(n_124), .C(n_98), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_226), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g250 ( .A1(n_247), .A2(n_210), .B1(n_213), .B2(n_200), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_230), .A2(n_193), .B(n_213), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_233), .B(n_215), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_241), .B(n_217), .Y(n_253) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_241), .A2(n_217), .A3(n_214), .B(n_119), .Y(n_254) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_226), .A2(n_124), .B1(n_102), .B2(n_189), .C(n_154), .Y(n_255) );
OAI222xp33_ASAP7_75t_L g256 ( .A1(n_242), .A2(n_93), .B1(n_103), .B2(n_101), .C1(n_99), .C2(n_97), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_242), .A2(n_221), .B1(n_192), .B2(n_195), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_235), .A2(n_199), .B1(n_198), .B2(n_194), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_244), .B(n_165), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_154), .B1(n_182), .B2(n_171), .C(n_178), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_224), .A2(n_199), .B1(n_198), .B2(n_194), .Y(n_261) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_107), .B(n_93), .C(n_103), .Y(n_262) );
OAI21xp33_ASAP7_75t_L g263 ( .A1(n_239), .A2(n_109), .B(n_216), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_244), .A2(n_185), .B1(n_191), .B2(n_211), .Y(n_264) );
OAI21xp33_ASAP7_75t_SL g265 ( .A1(n_222), .A2(n_171), .B(n_182), .Y(n_265) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_222), .A2(n_97), .B(n_99), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_222), .B(n_165), .Y(n_267) );
OAI211xp5_ASAP7_75t_L g268 ( .A1(n_243), .A2(n_101), .B(n_105), .C(n_109), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_238), .B(n_116), .C(n_114), .Y(n_269) );
OAI211xp5_ASAP7_75t_SL g270 ( .A1(n_223), .A2(n_105), .B(n_129), .C(n_126), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_254), .Y(n_271) );
OAI211xp5_ASAP7_75t_L g272 ( .A1(n_258), .A2(n_229), .B(n_223), .C(n_246), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_267), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_249), .B(n_100), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_252), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_253), .Y(n_276) );
OAI221xp5_ASAP7_75t_L g277 ( .A1(n_255), .A2(n_227), .B1(n_245), .B2(n_234), .C(n_238), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g278 ( .A(n_265), .B(n_248), .C(n_228), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_252), .B(n_228), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_250), .A2(n_232), .B1(n_225), .B2(n_248), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
AOI33xp33_ASAP7_75t_L g282 ( .A1(n_249), .A2(n_129), .A3(n_126), .B1(n_127), .B2(n_119), .B3(n_145), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_254), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_225), .B1(n_248), .B2(n_228), .C(n_201), .Y(n_285) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_251), .A2(n_127), .B(n_129), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_257), .A2(n_232), .B1(n_225), .B2(n_201), .Y(n_287) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_267), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_254), .B(n_232), .Y(n_289) );
AOI222xp33_ASAP7_75t_L g290 ( .A1(n_256), .A2(n_178), .B1(n_232), .B2(n_81), .C1(n_179), .C2(n_180), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_254), .Y(n_291) );
NAND4xp25_ASAP7_75t_SL g292 ( .A(n_265), .B(n_3), .C(n_4), .D(n_5), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_292), .A2(n_251), .B1(n_261), .B2(n_270), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_275), .B(n_266), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_278), .A2(n_268), .B(n_263), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_281), .B(n_276), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_275), .B(n_259), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_288), .B(n_259), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_276), .B(n_266), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_289), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_266), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_271), .B(n_269), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_284), .B(n_269), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_289), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_272), .B(n_3), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_284), .B(n_240), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_290), .A2(n_260), .B1(n_264), .B2(n_263), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_283), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_279), .B(n_264), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_279), .B(n_4), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_291), .Y(n_315) );
OAI31xp33_ASAP7_75t_L g316 ( .A1(n_277), .A2(n_165), .A3(n_180), .B(n_179), .Y(n_316) );
AND2x4_ASAP7_75t_SL g317 ( .A(n_281), .B(n_236), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_286), .Y(n_319) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_286), .B(n_240), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_273), .B(n_81), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_313), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_308), .A2(n_274), .B1(n_81), .B2(n_287), .C(n_280), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_301), .B(n_273), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_313), .Y(n_326) );
NAND4xp25_ASAP7_75t_SL g327 ( .A(n_301), .B(n_282), .C(n_285), .D(n_8), .Y(n_327) );
OAI211xp5_ASAP7_75t_L g328 ( .A1(n_321), .A2(n_273), .B(n_81), .C(n_91), .Y(n_328) );
NAND2xp33_ASAP7_75t_SL g329 ( .A(n_314), .B(n_273), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_311), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_306), .B(n_273), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_316), .A2(n_286), .B1(n_81), .B2(n_240), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_81), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_311), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
AOI211x1_ASAP7_75t_L g337 ( .A1(n_296), .A2(n_5), .B(n_6), .C(n_8), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_315), .B(n_119), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_315), .B(n_126), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_127), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_307), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_294), .B(n_9), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_297), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_296), .B(n_10), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_314), .B(n_11), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_307), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_302), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_303), .B(n_114), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_298), .B(n_12), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_298), .B(n_12), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g357 ( .A(n_316), .B(n_75), .C(n_92), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_309), .B(n_114), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_309), .B(n_114), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_299), .B(n_14), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_321), .B(n_14), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_312), .B(n_15), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_309), .B(n_116), .Y(n_364) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_322), .B(n_236), .Y(n_365) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_293), .B(n_15), .C(n_16), .D(n_17), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_353), .B(n_312), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_331), .B(n_322), .Y(n_368) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_362), .A2(n_322), .B(n_310), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_342), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_353), .B(n_318), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_343), .B(n_299), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_343), .B(n_309), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_325), .B(n_317), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_354), .B(n_318), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_331), .B(n_305), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_330), .Y(n_378) );
NOR2x2_ASAP7_75t_L g379 ( .A(n_366), .B(n_16), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_325), .B(n_317), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_354), .B(n_319), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_358), .B(n_293), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_358), .B(n_304), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_334), .B(n_305), .Y(n_385) );
INVxp33_ASAP7_75t_SL g386 ( .A(n_346), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_363), .B(n_317), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_304), .Y(n_388) );
XNOR2x1_ASAP7_75t_L g389 ( .A(n_363), .B(n_18), .Y(n_389) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_324), .A2(n_310), .B(n_295), .C(n_320), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_365), .A2(n_320), .B(n_319), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_335), .B(n_305), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_352), .B(n_305), .Y(n_394) );
AOI322xp5_ASAP7_75t_L g395 ( .A1(n_329), .A2(n_304), .A3(n_19), .B1(n_20), .B2(n_22), .C1(n_23), .C2(n_18), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_340), .B(n_19), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_361), .B(n_22), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_349), .B(n_295), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_341), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_334), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_337), .B(n_114), .C(n_116), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_349), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_359), .B(n_116), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_351), .B(n_116), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_116), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_351), .B(n_116), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_323), .B(n_236), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_350), .B(n_236), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_323), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_350), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_326), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_360), .B(n_24), .Y(n_413) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_348), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_326), .B(n_236), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_345), .A2(n_94), .B1(n_96), .B2(n_143), .C(n_137), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_336), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_336), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_370), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_383), .B(n_347), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_398), .B(n_347), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_389), .A2(n_357), .B(n_328), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_374), .B(n_333), .Y(n_423) );
XOR2x2_ASAP7_75t_L g424 ( .A(n_386), .B(n_356), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_403), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_SL g427 ( .A1(n_397), .A2(n_355), .B(n_327), .C(n_360), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_371), .B(n_344), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_380), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_371), .B(n_344), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_367), .B(n_375), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_369), .B(n_332), .C(n_333), .D(n_365), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_401), .A2(n_364), .B(n_348), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_393), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
NAND3x1_ASAP7_75t_L g437 ( .A(n_381), .B(n_333), .C(n_339), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_400), .B(n_364), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_382), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_382), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_414), .Y(n_442) );
OAI211xp5_ASAP7_75t_SL g443 ( .A1(n_395), .A2(n_143), .B(n_364), .C(n_180), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_375), .B(n_339), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_405), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_394), .B(n_364), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_372), .B(n_338), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_373), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_384), .B(n_338), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_402), .B(n_25), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_390), .A2(n_191), .B(n_190), .C(n_185), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_392), .B(n_26), .Y(n_454) );
XNOR2x1_ASAP7_75t_L g455 ( .A(n_396), .B(n_27), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_368), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_392), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g460 ( .A(n_368), .B(n_191), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_387), .B(n_28), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_417), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_418), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_394), .B(n_29), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g466 ( .A(n_413), .B(n_31), .Y(n_466) );
NOR3x1_ASAP7_75t_L g467 ( .A(n_379), .B(n_33), .C(n_34), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_377), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_385), .A2(n_185), .B1(n_190), .B2(n_211), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_377), .B(n_37), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_391), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_409), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_388), .B(n_38), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_385), .A2(n_185), .B1(n_190), .B2(n_211), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_404), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_406), .B(n_39), .Y(n_476) );
AO221x1_ASAP7_75t_L g477 ( .A1(n_408), .A2(n_185), .B1(n_41), .B2(n_43), .C(n_44), .Y(n_477) );
OAI21xp33_ASAP7_75t_SL g478 ( .A1(n_408), .A2(n_40), .B(n_46), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_416), .A2(n_179), .B(n_143), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_415), .B(n_49), .Y(n_480) );
OAI31xp33_ASAP7_75t_L g481 ( .A1(n_415), .A2(n_143), .A3(n_153), .B(n_144), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_411), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_376), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_370), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_383), .B(n_52), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_411), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_368), .Y(n_487) );
AOI322xp5_ASAP7_75t_L g488 ( .A1(n_383), .A2(n_56), .A3(n_57), .B1(n_58), .B2(n_60), .C1(n_61), .C2(n_62), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_390), .A2(n_137), .B1(n_153), .B2(n_144), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_394), .B(n_64), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_376), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_383), .A2(n_137), .B1(n_153), .B2(n_144), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_370), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_478), .A2(n_419), .B(n_484), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_484), .A2(n_487), .B1(n_456), .B2(n_419), .Y(n_495) );
AOI221xp5_ASAP7_75t_SL g496 ( .A1(n_493), .A2(n_466), .B1(n_433), .B2(n_448), .C(n_432), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
O2A1O1Ixp5_ASAP7_75t_L g498 ( .A1(n_420), .A2(n_440), .B(n_439), .C(n_471), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_457), .B(n_442), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_475), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_424), .A2(n_437), .B1(n_446), .B2(n_422), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_424), .A2(n_437), .B1(n_446), .B2(n_438), .Y(n_502) );
OAI322xp33_ASAP7_75t_L g503 ( .A1(n_421), .A2(n_447), .A3(n_425), .B1(n_450), .B2(n_453), .C1(n_441), .C2(n_445), .Y(n_503) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_455), .B(n_466), .Y(n_504) );
AOI322xp5_ASAP7_75t_L g505 ( .A1(n_487), .A2(n_423), .A3(n_468), .B1(n_490), .B2(n_472), .C1(n_444), .C2(n_429), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_455), .A2(n_468), .B1(n_490), .B2(n_443), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_483), .B(n_491), .Y(n_507) );
AOI21x1_ASAP7_75t_L g508 ( .A1(n_470), .A2(n_434), .B(n_471), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_461), .A2(n_472), .B1(n_460), .B2(n_426), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g510 ( .A1(n_467), .A2(n_473), .B1(n_461), .B2(n_489), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_488), .B(n_427), .C(n_452), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_501), .A2(n_428), .B(n_431), .Y(n_512) );
NAND4xp25_ASAP7_75t_SL g513 ( .A(n_496), .B(n_467), .C(n_470), .D(n_452), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_496), .A2(n_427), .B1(n_430), .B2(n_436), .C(n_435), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_502), .A2(n_491), .B1(n_483), .B2(n_485), .C(n_465), .Y(n_515) );
AOI322xp5_ASAP7_75t_L g516 ( .A1(n_504), .A2(n_451), .A3(n_462), .B1(n_459), .B2(n_458), .C1(n_463), .C2(n_464), .Y(n_516) );
NAND3xp33_ASAP7_75t_SL g517 ( .A(n_494), .B(n_481), .C(n_473), .Y(n_517) );
AOI211x1_ASAP7_75t_L g518 ( .A1(n_495), .A2(n_469), .B(n_474), .C(n_454), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_507), .Y(n_519) );
OAI211xp5_ASAP7_75t_L g520 ( .A1(n_511), .A2(n_476), .B(n_492), .C(n_480), .Y(n_520) );
NAND3x1_ASAP7_75t_L g521 ( .A(n_514), .B(n_508), .C(n_506), .Y(n_521) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_513), .B(n_497), .Y(n_522) );
NOR3x1_ASAP7_75t_L g523 ( .A(n_517), .B(n_477), .C(n_510), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_515), .A2(n_500), .B1(n_509), .B2(n_499), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_519), .B(n_449), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_525), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_522), .A2(n_518), .B1(n_512), .B2(n_520), .Y(n_527) );
OAI222xp33_ASAP7_75t_L g528 ( .A1(n_524), .A2(n_516), .B1(n_505), .B2(n_503), .C1(n_498), .C2(n_486), .Y(n_528) );
AOI22x1_ASAP7_75t_L g529 ( .A1(n_526), .A2(n_521), .B1(n_523), .B2(n_477), .Y(n_529) );
NOR2x2_ASAP7_75t_L g530 ( .A(n_527), .B(n_486), .Y(n_530) );
XNOR2x1_ASAP7_75t_L g531 ( .A(n_529), .B(n_530), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_531), .Y(n_532) );
XNOR2xp5_ASAP7_75t_L g533 ( .A(n_532), .B(n_528), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_533), .A2(n_482), .B1(n_464), .B2(n_479), .Y(n_534) );
endmodule