module fake_jpeg_25763_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_56),
.B1(n_49),
.B2(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_52),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_77),
.B(n_1),
.C(n_2),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_76),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_56),
.B1(n_54),
.B2(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_44),
.B1(n_43),
.B2(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_49),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_52),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_57),
.B1(n_55),
.B2(n_50),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_57),
.B1(n_50),
.B2(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_96),
.B1(n_74),
.B2(n_79),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_91),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_95),
.B(n_81),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_1),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_17),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_3),
.C(n_4),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_20),
.B1(n_40),
.B2(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_86),
.B1(n_95),
.B2(n_88),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_15),
.C(n_36),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_3),
.C(n_4),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_107),
.B(n_103),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_97),
.B(n_100),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_114),
.B1(n_14),
.B2(n_32),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_96),
.B1(n_82),
.B2(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_104),
.Y(n_117)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_21),
.B1(n_41),
.B2(n_33),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_97),
.B(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_116),
.B(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_118),
.B1(n_110),
.B2(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_123),
.B1(n_122),
.B2(n_24),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_11),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_13),
.C(n_30),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_29),
.C(n_27),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_5),
.B(n_6),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_6),
.B(n_7),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_7),
.B(n_8),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_8),
.Y(n_134)
);


endmodule