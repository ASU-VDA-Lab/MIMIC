module fake_netlist_1_1084_n_652 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_652);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_652;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_17), .Y(n_78) );
INVxp33_ASAP7_75t_SL g79 ( .A(n_43), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_13), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_26), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_59), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_54), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_42), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_20), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_70), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_35), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_77), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_75), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_65), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_32), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_38), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_2), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_17), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_61), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_63), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_73), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_53), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_55), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_74), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_60), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_76), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_45), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_57), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_48), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_1), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_66), .B(n_22), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_29), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_13), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_9), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_14), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_41), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_46), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_25), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_47), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_34), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_109), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_110), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_87), .B(n_0), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_91), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_103), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_83), .B(n_1), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_90), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_83), .B(n_2), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_92), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_116), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_87), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_124), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_78), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_98), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_124), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_122), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_118), .B(n_3), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_92), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_79), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_94), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_84), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_110), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_117), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_80), .Y(n_164) );
AND3x2_ASAP7_75t_L g165 ( .A(n_82), .B(n_4), .C(n_5), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_82), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_81), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_100), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_134), .B(n_96), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_144), .B(n_123), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_167), .B(n_106), .Y(n_171) );
CKINVDCx14_ASAP7_75t_R g172 ( .A(n_155), .Y(n_172) );
AND3x4_ASAP7_75t_L g173 ( .A(n_144), .B(n_112), .C(n_99), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_144), .B(n_95), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
NAND3x1_ASAP7_75t_L g176 ( .A(n_166), .B(n_95), .C(n_96), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_134), .B(n_114), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_129), .B(n_111), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_130), .A2(n_111), .B1(n_114), .B2(n_115), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_131), .B(n_102), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_150), .B(n_115), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_152), .B(n_123), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_159), .B(n_119), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_152), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_131), .B(n_119), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_132), .B(n_121), .Y(n_199) );
OR2x2_ASAP7_75t_SL g200 ( .A(n_164), .B(n_121), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_146), .Y(n_201) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_133), .B(n_120), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_126), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_168), .B(n_104), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_132), .B(n_120), .Y(n_206) );
NAND2xp33_ASAP7_75t_L g207 ( .A(n_156), .B(n_113), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_136), .B(n_113), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g212 ( .A(n_137), .B(n_107), .C(n_97), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_146), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_139), .B(n_105), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_139), .B(n_107), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
NAND3x1_ASAP7_75t_L g220 ( .A(n_166), .B(n_94), .C(n_97), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_140), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_145), .B(n_108), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_145), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
AND2x6_ASAP7_75t_SL g225 ( .A(n_172), .B(n_135), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_179), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_213), .B(n_158), .Y(n_227) );
OR2x2_ASAP7_75t_SL g228 ( .A(n_176), .B(n_125), .Y(n_228) );
OR2x2_ASAP7_75t_SL g229 ( .A(n_176), .B(n_153), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_172), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_187), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_222), .B(n_158), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_179), .B(n_187), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_197), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_173), .A2(n_163), .B1(n_161), .B2(n_157), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_187), .B(n_142), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
XOR2xp5_ASAP7_75t_L g242 ( .A(n_181), .B(n_6), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_198), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_222), .B(n_126), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_222), .B(n_126), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_174), .B(n_165), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_200), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_199), .B(n_160), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_184), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_190), .B(n_88), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_181), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_198), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_174), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_173), .A2(n_154), .B1(n_127), .B2(n_151), .Y(n_259) );
AND3x2_ASAP7_75t_SL g260 ( .A(n_220), .B(n_160), .C(n_151), .Y(n_260) );
BUFx4f_ASAP7_75t_SL g261 ( .A(n_170), .Y(n_261) );
AOI22x1_ASAP7_75t_L g262 ( .A1(n_183), .A2(n_160), .B1(n_151), .B2(n_149), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_199), .B(n_149), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_199), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_192), .Y(n_265) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_212), .B(n_142), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_170), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_169), .Y(n_268) );
NOR2xp33_ASAP7_75t_R g269 ( .A(n_207), .B(n_142), .Y(n_269) );
NOR2xp33_ASAP7_75t_R g270 ( .A(n_207), .B(n_142), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_202), .B(n_149), .Y(n_271) );
NOR3xp33_ASAP7_75t_SL g272 ( .A(n_205), .B(n_101), .C(n_8), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_177), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_181), .A2(n_143), .B1(n_140), .B2(n_147), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g275 ( .A(n_174), .B(n_143), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_175), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_202), .B(n_143), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_194), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_171), .B(n_36), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_195), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_206), .B(n_140), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_206), .B(n_7), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_209), .B(n_147), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_209), .B(n_147), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
O2A1O1Ixp5_ASAP7_75t_L g290 ( .A1(n_280), .A2(n_205), .B(n_204), .C(n_191), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_257), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_241), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_240), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_241), .Y(n_294) );
BUFx2_ASAP7_75t_R g295 ( .A(n_230), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_247), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_240), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_247), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_231), .B(n_216), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_251), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_264), .B(n_216), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_240), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_284), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_284), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_257), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_238), .Y(n_307) );
BUFx12f_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
INVx3_ASAP7_75t_SL g309 ( .A(n_284), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_268), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_261), .A2(n_216), .B1(n_220), .B2(n_211), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_227), .B(n_224), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_251), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_235), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_234), .A2(n_191), .B(n_204), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_282), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
INVx4_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
AOI22xp5_ASAP7_75t_SL g320 ( .A1(n_242), .A2(n_215), .B1(n_185), .B2(n_223), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_233), .B(n_219), .Y(n_321) );
BUFx12f_ASAP7_75t_L g322 ( .A(n_225), .Y(n_322) );
INVxp33_ASAP7_75t_L g323 ( .A(n_235), .Y(n_323) );
AOI322xp5_ASAP7_75t_L g324 ( .A1(n_248), .A2(n_268), .A3(n_273), .B1(n_255), .B2(n_246), .C1(n_272), .C2(n_259), .Y(n_324) );
OAI21x1_ASAP7_75t_SL g325 ( .A1(n_267), .A2(n_218), .B(n_203), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_254), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_249), .A2(n_217), .B(n_183), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_239), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_279), .A2(n_196), .B1(n_217), .B2(n_210), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_265), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_239), .B(n_7), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_252), .B(n_10), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_250), .Y(n_337) );
INVx5_ASAP7_75t_L g338 ( .A(n_267), .Y(n_338) );
AND2x4_ASAP7_75t_SL g339 ( .A(n_246), .B(n_210), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_262), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_307), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_324), .B(n_274), .C(n_273), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_309), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_292), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_299), .B(n_256), .Y(n_347) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_332), .A2(n_269), .B(n_270), .C(n_248), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_307), .A2(n_253), .B1(n_237), .B2(n_287), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_294), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_294), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_316), .B(n_226), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_271), .B1(n_258), .B2(n_246), .C(n_276), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_299), .A2(n_269), .B1(n_270), .B2(n_249), .Y(n_355) );
AND2x6_ASAP7_75t_L g356 ( .A(n_289), .B(n_232), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_340), .A2(n_286), .B(n_285), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_299), .A2(n_263), .B1(n_232), .B2(n_245), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_313), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_314), .B(n_232), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_302), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_314), .B(n_236), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_291), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_303), .A2(n_263), .B1(n_244), .B2(n_277), .Y(n_365) );
AO31x2_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_186), .A3(n_196), .B(n_203), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_336), .B(n_283), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_303), .A2(n_266), .B(n_260), .C(n_186), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_318), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_304), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_333), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_320), .A2(n_275), .B1(n_260), .B2(n_228), .C(n_229), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_296), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_304), .B(n_275), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_358), .A2(n_325), .B(n_290), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_373), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_373), .B(n_296), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_349), .B(n_329), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_372), .A2(n_310), .B1(n_291), .B2(n_322), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_361), .B(n_336), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_344), .A2(n_310), .B1(n_322), .B2(n_308), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_344), .A2(n_308), .B1(n_312), .B2(n_334), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_343), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_358), .A2(n_325), .B(n_328), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g386 ( .A1(n_341), .A2(n_306), .B1(n_300), .B2(n_331), .C1(n_327), .C2(n_326), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_354), .B(n_326), .C(n_298), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_369), .A2(n_333), .B(n_298), .Y(n_388) );
OR2x6_ASAP7_75t_L g389 ( .A(n_342), .B(n_301), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_327), .B1(n_300), .B2(n_331), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_341), .A2(n_288), .B1(n_306), .B2(n_323), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_367), .A2(n_321), .B1(n_315), .B2(n_335), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_342), .A2(n_229), .B1(n_228), .B2(n_295), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_367), .A2(n_335), .B1(n_339), .B2(n_318), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_353), .A2(n_330), .B1(n_339), .B2(n_337), .C(n_318), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_367), .A2(n_289), .B1(n_305), .B2(n_297), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_319), .B1(n_293), .B2(n_221), .C(n_305), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_342), .A2(n_338), .B1(n_317), .B2(n_302), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_368), .A2(n_221), .B(n_146), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_347), .A2(n_319), .B1(n_293), .B2(n_297), .C(n_146), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_377), .B(n_350), .Y(n_404) );
AOI21x1_ASAP7_75t_L g405 ( .A1(n_401), .A2(n_370), .B(n_371), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_394), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_379), .A2(n_359), .B1(n_348), .B2(n_365), .C(n_345), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_375), .A2(n_365), .B(n_371), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_382), .A2(n_345), .B1(n_342), .B2(n_370), .C(n_350), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
NAND2xp33_ASAP7_75t_R g412 ( .A(n_389), .B(n_369), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_391), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_389), .A2(n_360), .B1(n_352), .B2(n_357), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_388), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_391), .Y(n_417) );
AO21x2_ASAP7_75t_L g418 ( .A1(n_375), .A2(n_357), .B(n_352), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_384), .B(n_362), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_378), .A3(n_387), .B(n_390), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_383), .A2(n_367), .B1(n_363), .B2(n_361), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_392), .A2(n_374), .B1(n_369), .B2(n_362), .C(n_293), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_387), .A2(n_374), .B1(n_361), .B2(n_363), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_398), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_381), .B(n_361), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_389), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_381), .A2(n_363), .B1(n_374), .B2(n_356), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_389), .A2(n_363), .B1(n_302), .B2(n_317), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_381), .B(n_362), .Y(n_434) );
OAI211xp5_ASAP7_75t_SL g435 ( .A1(n_393), .A2(n_319), .B(n_11), .C(n_12), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_413), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_404), .B(n_401), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_427), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_396), .B1(n_402), .B2(n_395), .Y(n_439) );
AND2x4_ASAP7_75t_SL g440 ( .A(n_429), .B(n_397), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_399), .B1(n_356), .B2(n_401), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_404), .B(n_401), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_409), .B(n_10), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_427), .B(n_366), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_426), .B(n_385), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_409), .B(n_366), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_406), .A2(n_356), .B1(n_400), .B2(n_351), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_429), .B(n_351), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_426), .B(n_366), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_411), .B(n_366), .Y(n_453) );
INVx5_ASAP7_75t_L g454 ( .A(n_419), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_403), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_423), .A2(n_147), .B1(n_338), .B2(n_351), .C(n_193), .Y(n_456) );
OAI33xp33_ASAP7_75t_L g457 ( .A1(n_435), .A2(n_11), .A3(n_12), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_422), .B(n_351), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_411), .B(n_15), .Y(n_459) );
INVx5_ASAP7_75t_L g460 ( .A(n_419), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_415), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_413), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_421), .Y(n_465) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_405), .A2(n_366), .B(n_351), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_431), .B(n_356), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_421), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_410), .A2(n_422), .B1(n_424), .B2(n_435), .C(n_432), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_410), .A2(n_18), .A3(n_356), .B(n_23), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_418), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
BUFx2_ASAP7_75t_SL g476 ( .A(n_419), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_428), .B(n_18), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_412), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_430), .A2(n_356), .B1(n_317), .B2(n_302), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_430), .B(n_147), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_424), .A2(n_147), .B1(n_338), .B2(n_208), .C(n_214), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_461), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_438), .B(n_428), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_450), .B(n_425), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_462), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_437), .B(n_442), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_437), .B(n_420), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_452), .B(n_434), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_469), .B(n_425), .C(n_434), .D(n_431), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_444), .B(n_416), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_462), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_465), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_457), .B(n_414), .C(n_433), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_468), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_436), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_442), .B(n_416), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_445), .B(n_408), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_445), .B(n_408), .Y(n_499) );
NAND2x1_ASAP7_75t_L g500 ( .A(n_468), .B(n_431), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_408), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_455), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_471), .B(n_408), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_448), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_473), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_463), .Y(n_507) );
HB1xp67_ASAP7_75t_SL g508 ( .A(n_476), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_444), .B(n_418), .Y(n_509) );
NOR2xp33_ASAP7_75t_R g510 ( .A(n_449), .B(n_405), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_459), .B(n_418), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_473), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_443), .B(n_418), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_478), .A2(n_356), .B(n_24), .C(n_27), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_453), .B(n_317), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
NAND2xp33_ASAP7_75t_R g517 ( .A(n_467), .B(n_21), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_470), .B(n_28), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_477), .B(n_30), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_446), .B(n_31), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_453), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_470), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_446), .B(n_33), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_440), .B(n_37), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_464), .B(n_39), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_440), .B(n_40), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_451), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_454), .B(n_44), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_464), .B(n_49), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_476), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_441), .A2(n_214), .B(n_208), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_454), .B(n_460), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_530), .A2(n_472), .B(n_447), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_487), .B(n_454), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_496), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_482), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_487), .B(n_454), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_508), .A2(n_439), .B1(n_460), .B2(n_454), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_486), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_517), .A2(n_458), .B1(n_481), .B2(n_456), .C(n_475), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_492), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_521), .B(n_475), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_494), .A2(n_480), .B(n_449), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_490), .A2(n_449), .B1(n_460), .B2(n_480), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_493), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_484), .B(n_460), .Y(n_546) );
NOR2xp33_ASAP7_75t_SL g547 ( .A(n_528), .B(n_460), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_517), .A2(n_460), .B1(n_467), .B2(n_474), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_531), .A2(n_466), .B(n_474), .Y(n_549) );
NAND4xp25_ASAP7_75t_L g550 ( .A(n_519), .B(n_479), .C(n_467), .D(n_56), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_519), .A2(n_467), .B1(n_317), .B2(n_338), .Y(n_552) );
OAI31xp33_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_466), .A3(n_52), .B(n_58), .Y(n_553) );
OAI31xp33_ASAP7_75t_L g554 ( .A1(n_514), .A2(n_466), .A3(n_64), .B(n_67), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_500), .A2(n_338), .B(n_201), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_520), .A2(n_50), .B(n_69), .C(n_72), .Y(n_556) );
AOI211xp5_ASAP7_75t_L g557 ( .A1(n_532), .A2(n_193), .B(n_201), .C(n_208), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_502), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_527), .B(n_193), .Y(n_559) );
BUFx2_ASAP7_75t_SL g560 ( .A(n_528), .Y(n_560) );
XNOR2x1_ASAP7_75t_L g561 ( .A(n_489), .B(n_193), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_528), .Y(n_564) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_525), .B(n_201), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_483), .Y(n_566) );
BUFx3_ASAP7_75t_L g567 ( .A(n_523), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_523), .A2(n_208), .B(n_214), .C(n_515), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_505), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_506), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
NAND2xp33_ASAP7_75t_SL g572 ( .A(n_510), .B(n_214), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_522), .Y(n_573) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_513), .A2(n_511), .B(n_526), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_491), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_510), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_497), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_488), .B(n_498), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_483), .Y(n_579) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_550), .B(n_524), .Y(n_580) );
XNOR2x1_ASAP7_75t_L g581 ( .A(n_561), .B(n_485), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_572), .B(n_509), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_577), .B(n_563), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_536), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_578), .B(n_498), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_533), .A2(n_499), .B1(n_503), .B2(n_529), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_539), .Y(n_588) );
XNOR2xp5_ASAP7_75t_L g589 ( .A(n_534), .B(n_499), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_545), .Y(n_591) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_543), .A2(n_503), .B1(n_518), .B2(n_504), .C1(n_507), .C2(n_516), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_537), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_551), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_566), .Y(n_595) );
XNOR2xp5_ASAP7_75t_L g596 ( .A(n_575), .B(n_518), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_546), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_566), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_579), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_560), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_576), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_558), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_535), .B(n_504), .Y(n_603) );
XNOR2x2_ASAP7_75t_L g604 ( .A(n_540), .B(n_507), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_569), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_574), .A2(n_516), .B(n_540), .C(n_568), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_548), .A2(n_554), .B(n_553), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_570), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_571), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_562), .B(n_573), .Y(n_610) );
AO22x1_ASAP7_75t_L g611 ( .A1(n_600), .A2(n_567), .B1(n_538), .B2(n_564), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_610), .B(n_542), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_593), .B(n_544), .Y(n_613) );
NAND4xp75_ASAP7_75t_L g614 ( .A(n_607), .B(n_565), .C(n_549), .D(n_555), .Y(n_614) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_582), .B(n_548), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_587), .A2(n_547), .B1(n_552), .B2(n_559), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_601), .Y(n_617) );
OAI31xp33_ASAP7_75t_L g618 ( .A1(n_581), .A2(n_556), .A3(n_549), .B(n_555), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_581), .A2(n_556), .B1(n_557), .B2(n_580), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_586), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_584), .B(n_609), .Y(n_621) );
OAI31xp33_ASAP7_75t_L g622 ( .A1(n_604), .A2(n_596), .A3(n_582), .B(n_606), .Y(n_622) );
XNOR2x1_ASAP7_75t_L g623 ( .A(n_604), .B(n_583), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_597), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_592), .A2(n_608), .B1(n_588), .B2(n_602), .C(n_590), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_591), .B(n_605), .Y(n_626) );
OAI211xp5_ASAP7_75t_SL g627 ( .A1(n_622), .A2(n_594), .B(n_585), .C(n_595), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_617), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_620), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_624), .B(n_595), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_618), .A2(n_598), .B(n_599), .C(n_603), .Y(n_631) );
CKINVDCx16_ASAP7_75t_R g632 ( .A(n_619), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_615), .B(n_599), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_625), .A2(n_589), .B1(n_598), .B2(n_626), .C(n_621), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_611), .B(n_616), .C(n_626), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_613), .A2(n_614), .B1(n_621), .B2(n_612), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_622), .A2(n_618), .B(n_625), .C(n_617), .Y(n_637) );
AO22x2_ASAP7_75t_L g638 ( .A1(n_623), .A2(n_617), .B1(n_614), .B2(n_601), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_622), .B(n_618), .C(n_619), .D(n_615), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_628), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_628), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_629), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_635), .A2(n_632), .B1(n_638), .B2(n_636), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_639), .B(n_637), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_643), .B(n_634), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_644), .B(n_627), .C(n_631), .D(n_633), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_640), .Y(n_647) );
OAI22xp5_ASAP7_75t_SL g648 ( .A1(n_645), .A2(n_644), .B1(n_641), .B2(n_630), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_646), .B(n_642), .Y(n_649) );
BUFx2_ASAP7_75t_SL g650 ( .A(n_649), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_650), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_SL g652 ( .A1(n_651), .A2(n_647), .B(n_648), .C(n_633), .Y(n_652) );
endmodule