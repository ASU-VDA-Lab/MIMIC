module fake_netlist_6_1397_n_770 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_770);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_770;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_605;
wire n_230;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_550;
wire n_487;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx5_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_31),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_49),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_38),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_98),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_48),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_63),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_66),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_69),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_39),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_86),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_43),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_52),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_119),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_62),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_85),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_95),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_42),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_47),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_8),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_20),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_23),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_25),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_57),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_34),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_4),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_46),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_128),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_116),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_41),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_136),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_0),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_0),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_173),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_1),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_3),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_4),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_5),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_6),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_208),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_6),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_152),
.B(n_7),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_173),
.B(n_7),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_8),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_177),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_152),
.B(n_9),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_161),
.B(n_21),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_163),
.B(n_9),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_10),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_209),
.B1(n_193),
.B2(n_200),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_217),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_156),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_157),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_195),
.B1(n_198),
.B2(n_187),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_160),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_232),
.A2(n_206),
.B1(n_166),
.B2(n_204),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_205),
.B1(n_182),
.B2(n_202),
.Y(n_261)
);

AOI22x1_ASAP7_75t_SL g262 ( 
.A1(n_215),
.A2(n_203),
.B1(n_199),
.B2(n_196),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_212),
.A2(n_189),
.B1(n_188),
.B2(n_185),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_223),
.B(n_159),
.Y(n_264)
);

AO22x2_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_152),
.B1(n_11),
.B2(n_12),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_152),
.B1(n_11),
.B2(n_13),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_165),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_169),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_183),
.B1(n_181),
.B2(n_178),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_239),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_246),
.A2(n_174),
.B1(n_171),
.B2(n_170),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_152),
.B1(n_13),
.B2(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_22),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_233),
.B(n_10),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_24),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_219),
.A2(n_214),
.B1(n_237),
.B2(n_225),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_26),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g286 ( 
.A1(n_237),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_221),
.A2(n_224),
.B1(n_243),
.B2(n_234),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_27),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_17),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_19),
.B1(n_29),
.B2(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_228),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_236),
.B(n_240),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_SL g301 ( 
.A(n_236),
.B(n_51),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_231),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_263),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_231),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_218),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_260),
.B(n_245),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_262),
.Y(n_320)
);

XNOR2x2_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_215),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_248),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

OR2x6_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_248),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_242),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_270),
.B(n_250),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_253),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_240),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_258),
.B(n_241),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_269),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_278),
.B(n_241),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_274),
.A2(n_244),
.B(n_218),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_278),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_242),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_242),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g352 ( 
.A(n_265),
.B(n_240),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_274),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_286),
.B(n_216),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_261),
.B(n_240),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_265),
.B(n_216),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_265),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_266),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_266),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_261),
.B(n_240),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_266),
.B(n_216),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_258),
.B(n_216),
.Y(n_363)
);

NAND2x1p5_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_216),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_249),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_303),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_244),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_244),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_249),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_348),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_244),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_295),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_316),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_249),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_344),
.A2(n_244),
.B(n_297),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_336),
.B(n_249),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_249),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_250),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_304),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_304),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_309),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_312),
.B(n_250),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_250),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_328),
.B(n_250),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_213),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_313),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_356),
.A2(n_301),
.B(n_238),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_213),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_330),
.B(n_238),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_314),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_355),
.B(n_238),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_238),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_360),
.B(n_238),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_315),
.B(n_54),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_315),
.B(n_55),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_330),
.B(n_227),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_306),
.B(n_360),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_319),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_320),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_227),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_306),
.B(n_227),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_227),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_318),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_318),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_336),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_326),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_308),
.B(n_227),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_368),
.B(n_346),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_339),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_362),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_346),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_376),
.B(n_365),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_308),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_374),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_420),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_426),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_359),
.Y(n_451)
);

BUFx8_ASAP7_75t_L g452 ( 
.A(n_434),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_326),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_426),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_326),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_343),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_374),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_383),
.B(n_318),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_383),
.B(n_316),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_379),
.B(n_385),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_378),
.Y(n_464)
);

CKINVDCx10_ASAP7_75t_R g465 ( 
.A(n_434),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_385),
.B(n_354),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_364),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_382),
.B(n_56),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_364),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_334),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_435),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_352),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_394),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_379),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_426),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_429),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_352),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_373),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_427),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_382),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

BUFx5_ASAP7_75t_L g487 ( 
.A(n_375),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_412),
.B(n_347),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_431),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_391),
.B(n_423),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_410),
.B(n_351),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

BUFx12f_ASAP7_75t_L g494 ( 
.A(n_452),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_455),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_448),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_439),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_473),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_428),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_455),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_479),
.B(n_428),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_432),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_441),
.B(n_432),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

INVx8_ASAP7_75t_L g517 ( 
.A(n_468),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_465),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_452),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

BUFx2_ASAP7_75t_SL g523 ( 
.A(n_456),
.Y(n_523)
);

BUFx4f_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_439),
.A2(n_428),
.B1(n_426),
.B2(n_416),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_491),
.Y(n_527)
);

BUFx4f_ASAP7_75t_SL g528 ( 
.A(n_452),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_440),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_456),
.Y(n_532)
);

INVx3_ASAP7_75t_SL g533 ( 
.A(n_457),
.Y(n_533)
);

CKINVDCx8_ASAP7_75t_R g534 ( 
.A(n_440),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_437),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_479),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_496),
.A2(n_463),
.B1(n_321),
.B2(n_472),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_502),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_529),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_537),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_502),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_508),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_505),
.A2(n_463),
.B1(n_426),
.B2(n_432),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

BUFx2_ASAP7_75t_SL g547 ( 
.A(n_498),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_494),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_505),
.A2(n_453),
.B1(n_451),
.B2(n_443),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_493),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_516),
.A2(n_451),
.B1(n_466),
.B2(n_430),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_537),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_527),
.B(n_474),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_531),
.A2(n_451),
.B1(n_430),
.B2(n_467),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_506),
.Y(n_559)
);

OAI22xp33_ASAP7_75t_L g560 ( 
.A1(n_534),
.A2(n_446),
.B1(n_486),
.B2(n_462),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_534),
.A2(n_469),
.B1(n_481),
.B2(n_475),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_531),
.A2(n_436),
.B1(n_417),
.B2(n_411),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_495),
.B(n_436),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_503),
.B(n_458),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_499),
.Y(n_566)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_517),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_525),
.A2(n_411),
.B1(n_459),
.B2(n_449),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_500),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_533),
.A2(n_411),
.B1(n_384),
.B2(n_490),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_517),
.A2(n_395),
.B1(n_387),
.B2(n_468),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_533),
.A2(n_411),
.B1(n_480),
.B2(n_468),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

CKINVDCx6p67_ASAP7_75t_R g574 ( 
.A(n_506),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_514),
.Y(n_575)
);

CKINVDCx11_ASAP7_75t_R g576 ( 
.A(n_520),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_517),
.A2(n_395),
.B1(n_387),
.B2(n_425),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_538),
.A2(n_499),
.B1(n_504),
.B2(n_515),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_549),
.A2(n_504),
.B1(n_507),
.B2(n_510),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_545),
.A2(n_514),
.B1(n_523),
.B2(n_535),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_560),
.A2(n_532),
.B1(n_514),
.B2(n_399),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_566),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_569),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_539),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_557),
.A2(n_471),
.B1(n_477),
.B2(n_476),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_557),
.A2(n_399),
.B1(n_404),
.B2(n_409),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_564),
.A2(n_409),
.B1(n_398),
.B2(n_460),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_571),
.A2(n_406),
.B(n_518),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_571),
.A2(n_488),
.B(n_372),
.Y(n_589)
);

AOI222xp33_ASAP7_75t_L g590 ( 
.A1(n_569),
.A2(n_528),
.B1(n_511),
.B2(n_431),
.C1(n_427),
.C2(n_423),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_566),
.A2(n_528),
.B1(n_520),
.B2(n_511),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_565),
.A2(n_447),
.B1(n_444),
.B2(n_492),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_398),
.B(n_380),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_576),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_572),
.A2(n_524),
.B1(n_522),
.B2(n_449),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_539),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_562),
.A2(n_397),
.B1(n_400),
.B2(n_380),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_542),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_542),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_540),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_540),
.B(n_427),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_544),
.Y(n_602)
);

BUFx5_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_577),
.A2(n_372),
.B(n_415),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_543),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_544),
.Y(n_606)
);

CKINVDCx6p67_ASAP7_75t_R g607 ( 
.A(n_555),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_546),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_551),
.A2(n_400),
.B1(n_397),
.B2(n_403),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_563),
.A2(n_401),
.B(n_568),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_558),
.A2(n_397),
.B1(n_403),
.B2(n_407),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_553),
.A2(n_522),
.B1(n_524),
.B2(n_509),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_567),
.A2(n_522),
.B1(n_524),
.B2(n_509),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_546),
.A2(n_407),
.B1(n_414),
.B2(n_410),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_546),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_567),
.A2(n_513),
.B1(n_537),
.B2(n_498),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_575),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_567),
.A2(n_513),
.B1(n_498),
.B2(n_415),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_574),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_567),
.A2(n_498),
.B1(n_414),
.B2(n_375),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_543),
.A2(n_526),
.B1(n_521),
.B2(n_470),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_555),
.A2(n_526),
.B1(n_461),
.B2(n_388),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_579),
.A2(n_574),
.B1(n_388),
.B2(n_548),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_579),
.A2(n_559),
.B1(n_548),
.B2(n_556),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_578),
.A2(n_388),
.B1(n_552),
.B2(n_550),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_580),
.A2(n_575),
.B1(n_559),
.B2(n_425),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_593),
.A2(n_575),
.B1(n_487),
.B2(n_552),
.Y(n_631)
);

OAI222xp33_ASAP7_75t_L g632 ( 
.A1(n_581),
.A2(n_583),
.B1(n_591),
.B2(n_586),
.C1(n_587),
.C2(n_626),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_610),
.A2(n_547),
.B1(n_541),
.B2(n_556),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_584),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_588),
.A2(n_556),
.B1(n_541),
.B2(n_547),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_586),
.A2(n_541),
.B1(n_498),
.B2(n_408),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_590),
.A2(n_575),
.B1(n_487),
.B2(n_386),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_592),
.B(n_554),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_592),
.A2(n_487),
.B1(n_396),
.B2(n_454),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_582),
.B(n_561),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_598),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_600),
.B(n_561),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_617),
.A2(n_487),
.B1(n_454),
.B2(n_482),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_611),
.Y(n_644)
);

OAI221xp5_ASAP7_75t_L g645 ( 
.A1(n_589),
.A2(n_418),
.B1(n_422),
.B2(n_370),
.C(n_377),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_591),
.A2(n_607),
.B1(n_597),
.B2(n_609),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_597),
.A2(n_487),
.B1(n_454),
.B2(n_482),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_611),
.B(n_58),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_587),
.B(n_367),
.C(n_450),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_626),
.A2(n_601),
.B1(n_612),
.B2(n_608),
.Y(n_650)
);

OAI221xp5_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_373),
.B1(n_450),
.B2(n_482),
.C(n_389),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_608),
.A2(n_618),
.B1(n_620),
.B2(n_585),
.Y(n_652)
);

OAI21xp33_ASAP7_75t_L g653 ( 
.A1(n_585),
.A2(n_373),
.B(n_372),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_608),
.A2(n_487),
.B1(n_389),
.B2(n_392),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_595),
.A2(n_536),
.B1(n_530),
.B2(n_519),
.Y(n_655)
);

OAI221xp5_ASAP7_75t_L g656 ( 
.A1(n_623),
.A2(n_389),
.B1(n_392),
.B2(n_519),
.C(n_512),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_608),
.A2(n_392),
.B1(n_372),
.B2(n_536),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_596),
.A2(n_605),
.B1(n_594),
.B2(n_599),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_622),
.A2(n_619),
.B1(n_624),
.B2(n_618),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_625),
.A2(n_536),
.B1(n_530),
.B2(n_519),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_625),
.A2(n_536),
.B1(n_530),
.B2(n_519),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_618),
.A2(n_530),
.B1(n_512),
.B2(n_497),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_618),
.A2(n_392),
.B1(n_512),
.B2(n_497),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_620),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_646),
.A2(n_613),
.B1(n_615),
.B2(n_616),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_634),
.B(n_641),
.Y(n_666)
);

OAI21xp33_ASAP7_75t_SL g667 ( 
.A1(n_627),
.A2(n_621),
.B(n_614),
.Y(n_667)
);

NAND4xp25_ASAP7_75t_L g668 ( 
.A(n_658),
.B(n_606),
.C(n_602),
.D(n_603),
.Y(n_668)
);

AOI221xp5_ASAP7_75t_L g669 ( 
.A1(n_632),
.A2(n_512),
.B1(n_497),
.B2(n_393),
.C(n_390),
.Y(n_669)
);

OAI221xp5_ASAP7_75t_L g670 ( 
.A1(n_627),
.A2(n_630),
.B1(n_658),
.B2(n_628),
.C(n_659),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_633),
.A2(n_497),
.B(n_60),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_642),
.B(n_603),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_640),
.B(n_603),
.Y(n_673)
);

AOI221xp5_ASAP7_75t_L g674 ( 
.A1(n_635),
.A2(n_393),
.B1(n_390),
.B2(n_230),
.C(n_603),
.Y(n_674)
);

NAND4xp25_ASAP7_75t_L g675 ( 
.A(n_629),
.B(n_638),
.C(n_648),
.D(n_639),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_640),
.B(n_629),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_652),
.B(n_603),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_650),
.B(n_603),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_637),
.A2(n_393),
.B1(n_390),
.B2(n_230),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_655),
.B(n_653),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_662),
.B(n_390),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_643),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_649),
.B(n_59),
.Y(n_683)
);

OA211x2_ASAP7_75t_L g684 ( 
.A1(n_663),
.A2(n_61),
.B(n_64),
.C(n_65),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_651),
.A2(n_230),
.B(n_68),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_L g686 ( 
.A1(n_647),
.A2(n_393),
.B(n_390),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_636),
.B(n_67),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_664),
.B(n_656),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_666),
.B(n_660),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_661),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_672),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_673),
.Y(n_692)
);

NOR2x1_ASAP7_75t_L g693 ( 
.A(n_668),
.B(n_645),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_670),
.B(n_657),
.C(n_654),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_677),
.B(n_678),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_676),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_675),
.B(n_70),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_671),
.A2(n_393),
.B1(n_390),
.B2(n_230),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_71),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_665),
.B(n_72),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_675),
.A2(n_393),
.B1(n_74),
.B2(n_77),
.Y(n_701)
);

XOR2x2_ASAP7_75t_L g702 ( 
.A(n_696),
.B(n_669),
.Y(n_702)
);

XOR2x2_ASAP7_75t_L g703 ( 
.A(n_697),
.B(n_680),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_691),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_692),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_700),
.B(n_681),
.Y(n_706)
);

XOR2x2_ASAP7_75t_L g707 ( 
.A(n_699),
.B(n_687),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_695),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_695),
.Y(n_709)
);

NAND4xp75_ASAP7_75t_L g710 ( 
.A(n_693),
.B(n_684),
.C(n_685),
.D(n_674),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_689),
.Y(n_711)
);

XNOR2xp5_ASAP7_75t_L g712 ( 
.A(n_703),
.B(n_694),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_704),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_709),
.B(n_688),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_708),
.B(n_690),
.Y(n_715)
);

XOR2x2_ASAP7_75t_L g716 ( 
.A(n_703),
.B(n_701),
.Y(n_716)
);

OA22x2_ASAP7_75t_L g717 ( 
.A1(n_712),
.A2(n_711),
.B1(n_705),
.B2(n_704),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_713),
.Y(n_719)
);

XNOR2xp5_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_707),
.Y(n_720)
);

OAI22x1_ASAP7_75t_L g721 ( 
.A1(n_714),
.A2(n_702),
.B1(n_706),
.B2(n_710),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_719),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_720),
.B(n_698),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_718),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_717),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_725),
.A2(n_720),
.B1(n_721),
.B2(n_706),
.Y(n_726)
);

AOI211xp5_ASAP7_75t_SL g727 ( 
.A1(n_724),
.A2(n_679),
.B(n_683),
.C(n_686),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_726),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_727),
.A2(n_723),
.B1(n_722),
.B2(n_667),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_726),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_730),
.B(n_73),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_728),
.A2(n_230),
.B1(n_79),
.B2(n_80),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_729),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_729),
.Y(n_734)
);

NOR4xp25_ASAP7_75t_L g735 ( 
.A(n_728),
.B(n_78),
.C(n_81),
.D(n_82),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_728),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_733),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_736),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_734),
.B(n_83),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_731),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_732),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_735),
.B(n_84),
.Y(n_742)
);

NOR2x1_ASAP7_75t_L g743 ( 
.A(n_731),
.B(n_87),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_737),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_738),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

NOR4xp75_ASAP7_75t_L g748 ( 
.A(n_739),
.B(n_99),
.C(n_103),
.D(n_104),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_741),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_745),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_747),
.A2(n_743),
.B1(n_110),
.B2(n_111),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_746),
.B(n_109),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_749),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_748),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_744),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_745),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_754),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_757)
);

AND4x2_ASAP7_75t_L g758 ( 
.A(n_751),
.B(n_122),
.C(n_123),
.D(n_124),
.Y(n_758)
);

OAI22x1_ASAP7_75t_L g759 ( 
.A1(n_755),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_750),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_756),
.Y(n_761)
);

INVxp67_ASAP7_75t_SL g762 ( 
.A(n_759),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_761),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_762),
.A2(n_752),
.B1(n_757),
.B2(n_753),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_763),
.A2(n_760),
.B1(n_758),
.B2(n_138),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_765),
.B1(n_137),
.B2(n_139),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_767),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_135),
.B1(n_140),
.B2(n_145),
.C(n_146),
.Y(n_769)
);

AOI211xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_148),
.B(n_149),
.C(n_151),
.Y(n_770)
);


endmodule