module fake_jpeg_21982_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_34),
.B(n_1),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_26),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_8),
.Y(n_44)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_21),
.CON(n_57),
.SN(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_53),
.Y(n_85)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_19),
.B1(n_33),
.B2(n_27),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_19),
.B1(n_33),
.B2(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_58),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_19),
.B1(n_28),
.B2(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_72),
.B1(n_23),
.B2(n_18),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_30),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_64),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_33),
.B1(n_20),
.B2(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_30),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_77),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_17),
.B(n_24),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_71),
.B(n_32),
.C(n_29),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_27),
.B1(n_20),
.B2(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_28),
.B1(n_35),
.B2(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_91),
.Y(n_127)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_87),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_88),
.B(n_90),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_35),
.B1(n_21),
.B2(n_22),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_104),
.B(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_45),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_98),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_0),
.B(n_1),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_97),
.B(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_45),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_48),
.B1(n_49),
.B2(n_22),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_56),
.B1(n_29),
.B2(n_31),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_48),
.B(n_37),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_70),
.B1(n_79),
.B2(n_58),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_38),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_65),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_111),
.Y(n_146)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_43),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_115),
.Y(n_144)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_43),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_29),
.B1(n_31),
.B2(n_10),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_131),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_145),
.B1(n_84),
.B2(n_94),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_70),
.B1(n_58),
.B2(n_52),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_107),
.B(n_106),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_133),
.B1(n_150),
.B2(n_86),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_85),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_65),
.B1(n_31),
.B2(n_59),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_140),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_93),
.B(n_43),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_139),
.C(n_114),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_38),
.C(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_88),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_97),
.B1(n_90),
.B2(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_31),
.B1(n_62),
.B2(n_59),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_103),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_169),
.B1(n_130),
.B2(n_150),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_128),
.B1(n_143),
.B2(n_137),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_95),
.Y(n_157)
);

BUFx12f_ASAP7_75t_SL g158 ( 
.A(n_141),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_182),
.B(n_179),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_175),
.C(n_119),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_95),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_83),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_170),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_83),
.B1(n_85),
.B2(n_101),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_171),
.B1(n_9),
.B2(n_13),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_83),
.B1(n_81),
.B2(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_81),
.B1(n_110),
.B2(n_107),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_180),
.B(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_99),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_106),
.C(n_82),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_80),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_99),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_182),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_0),
.B(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_62),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_87),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_185),
.B(n_154),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_198),
.C(n_206),
.Y(n_217)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_128),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_196),
.B(n_201),
.C(n_204),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_203),
.B(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_132),
.C(n_151),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_212),
.B1(n_213),
.B2(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_138),
.B(n_137),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_138),
.B(n_12),
.C(n_15),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_208),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_165),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_118),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_208),
.Y(n_220)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_118),
.B1(n_134),
.B2(n_122),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_122),
.B1(n_149),
.B2(n_123),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_2),
.B(n_3),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_155),
.B1(n_168),
.B2(n_160),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_159),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_192),
.B(n_205),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_237),
.B1(n_240),
.B2(n_215),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_175),
.C(n_163),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_222),
.C(n_230),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_177),
.C(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_177),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_235),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_213),
.B1(n_204),
.B2(n_197),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_183),
.C(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_189),
.C(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_185),
.A2(n_164),
.B1(n_156),
.B2(n_160),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_166),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_196),
.A2(n_176),
.B1(n_165),
.B2(n_181),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_211),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_248),
.B1(n_216),
.B2(n_241),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_258),
.B(n_3),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_220),
.B1(n_236),
.B2(n_228),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_256),
.B1(n_13),
.B2(n_11),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_207),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_192),
.B(n_203),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_8),
.B(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_194),
.B1(n_193),
.B2(n_226),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_190),
.B1(n_191),
.B2(n_189),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_229),
.B1(n_216),
.B2(n_227),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_210),
.B(n_195),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_10),
.B(n_14),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_217),
.C(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_217),
.C(n_222),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_235),
.C(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_270),
.Y(n_286)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_277),
.B1(n_275),
.B2(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_165),
.C(n_195),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_261),
.C(n_258),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_276),
.Y(n_283)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_246),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_259),
.B1(n_255),
.B2(n_243),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_254),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_245),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_284),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_257),
.C(n_253),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_293),
.B(n_278),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_250),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_269),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_255),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_267),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_264),
.A2(n_259),
.B(n_10),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_272),
.B1(n_271),
.B2(n_263),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_301),
.B1(n_286),
.B2(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_287),
.C(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_268),
.B1(n_266),
.B2(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_302),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_281),
.C(n_292),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

OAI211xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_312),
.B(n_307),
.C(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_281),
.C(n_290),
.Y(n_310)
);

NAND5xp2_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_4),
.C(n_5),
.D(n_6),
.E(n_7),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_296),
.A3(n_300),
.B1(n_297),
.B2(n_8),
.C1(n_3),
.C2(n_6),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_318),
.B(n_4),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_317),
.B(n_4),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_316),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_4),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_322),
.B(n_5),
.Y(n_324)
);

AO21x2_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_6),
.B(n_7),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_6),
.C(n_7),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_7),
.Y(n_328)
);


endmodule