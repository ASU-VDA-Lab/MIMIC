module fake_netlist_1_5961_n_482 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_482);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_482;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g72 ( .A(n_3), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_69), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_50), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_65), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_27), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_13), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_9), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_25), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_6), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_67), .Y(n_83) );
OR2x2_ASAP7_75t_L g84 ( .A(n_23), .B(n_11), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_35), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_31), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_10), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_56), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_7), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_42), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_53), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_6), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_60), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_7), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_15), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_41), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_55), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_23), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_19), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_4), .Y(n_101) );
BUFx2_ASAP7_75t_SL g102 ( .A(n_66), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_4), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_10), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_95), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_95), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_86), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_87), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_87), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_87), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_95), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_95), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_94), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_86), .Y(n_114) );
OAI21x1_ASAP7_75t_L g115 ( .A1(n_88), .A2(n_34), .B(n_70), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_86), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_100), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_101), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_100), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_72), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_94), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_74), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_78), .B(n_0), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_86), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_113), .B(n_78), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_113), .B(n_94), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_120), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_107), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_108), .B(n_89), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_108), .B(n_89), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_113), .B(n_94), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_124), .B(n_88), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_115), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_113), .B(n_88), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_107), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_120), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_124), .B(n_90), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_114), .B(n_90), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_114), .B(n_90), .Y(n_149) );
AO22x2_ASAP7_75t_L g150 ( .A1(n_126), .A2(n_97), .B1(n_84), .B2(n_83), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
OR2x2_ASAP7_75t_SL g152 ( .A(n_126), .B(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_147), .A2(n_80), .B(n_84), .C(n_92), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_133), .Y(n_157) );
NOR2xp33_ASAP7_75t_R g158 ( .A(n_151), .B(n_117), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_128), .B(n_109), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_150), .A2(n_110), .B1(n_109), .B2(n_80), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_128), .B(n_110), .Y(n_161) );
AND3x2_ASAP7_75t_SL g162 ( .A(n_150), .B(n_127), .C(n_116), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
NOR2xp33_ASAP7_75t_R g164 ( .A(n_151), .B(n_125), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_130), .B(n_92), .Y(n_166) );
NOR2xp33_ASAP7_75t_R g167 ( .A(n_151), .B(n_121), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_145), .B(n_74), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_150), .A2(n_127), .B1(n_114), .B2(n_116), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_145), .B(n_85), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_150), .A2(n_127), .B1(n_114), .B2(n_116), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_134), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_134), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_150), .B(n_102), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVx6_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_134), .B(n_106), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_143), .Y(n_180) );
BUFx12f_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
CKINVDCx8_ASAP7_75t_R g183 ( .A(n_143), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_150), .A2(n_82), .B1(n_96), .B2(n_104), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_163), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_183), .A2(n_152), .B1(n_135), .B2(n_143), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_135), .B1(n_72), .B2(n_121), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_183), .A2(n_152), .B1(n_135), .B2(n_143), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_158), .Y(n_191) );
BUFx12f_ASAP7_75t_L g192 ( .A(n_174), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_179), .B(n_143), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_136), .B1(n_129), .B2(n_138), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_176), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_180), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_179), .B(n_129), .Y(n_200) );
OR2x6_ASAP7_75t_L g201 ( .A(n_181), .B(n_102), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_180), .B(n_129), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_159), .B(n_137), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_167), .A2(n_93), .B1(n_83), .B2(n_136), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_178), .B(n_136), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_161), .B(n_136), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_157), .A2(n_142), .B(n_137), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_175), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
AOI21xp5_ASAP7_75t_SL g211 ( .A1(n_175), .A2(n_142), .B(n_136), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_164), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_157), .A2(n_142), .B(n_138), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_175), .A2(n_146), .B1(n_148), .B2(n_142), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_171), .A2(n_142), .B(n_148), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_181), .A2(n_147), .B1(n_85), .B2(n_149), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_171), .A2(n_149), .B(n_115), .C(n_127), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_188), .B(n_166), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_188), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_209), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_204), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_209), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_204), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_193), .B(n_166), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_189), .A2(n_174), .B1(n_175), .B2(n_173), .Y(n_225) );
OAI211xp5_ASAP7_75t_L g226 ( .A1(n_205), .A2(n_184), .B(n_154), .C(n_169), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_186), .A2(n_175), .B1(n_166), .B2(n_177), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_186), .Y(n_228) );
OAI211xp5_ASAP7_75t_SL g229 ( .A1(n_196), .A2(n_184), .B(n_170), .C(n_172), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_187), .A2(n_166), .B1(n_182), .B2(n_185), .C(n_178), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_190), .A2(n_185), .B1(n_182), .B2(n_177), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_203), .A2(n_207), .B(n_194), .C(n_217), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_193), .A2(n_177), .B1(n_176), .B2(n_165), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_191), .A2(n_162), .B1(n_177), .B2(n_104), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_200), .B(n_176), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_216), .A2(n_82), .B1(n_99), .B2(n_77), .C(n_79), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_191), .A2(n_162), .B1(n_93), .B2(n_102), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_206), .B(n_165), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_197), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_236), .A2(n_231), .B1(n_225), .B2(n_227), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_219), .B(n_206), .Y(n_246) );
OAI221xp5_ASAP7_75t_L g247 ( .A1(n_238), .A2(n_201), .B1(n_212), .B2(n_214), .C(n_103), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_228), .A2(n_201), .B1(n_192), .B2(n_212), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_229), .A2(n_192), .B1(n_201), .B2(n_202), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_232), .A2(n_208), .B(n_211), .Y(n_250) );
AOI222xp33_ASAP7_75t_L g251 ( .A1(n_233), .A2(n_224), .B1(n_230), .B2(n_226), .C1(n_219), .C2(n_218), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_224), .A2(n_201), .B1(n_202), .B2(n_206), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g253 ( .A1(n_220), .A2(n_162), .B1(n_81), .B2(n_77), .Y(n_253) );
AOI21xp33_ASAP7_75t_L g254 ( .A1(n_239), .A2(n_195), .B(n_116), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_223), .B(n_211), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_223), .B(n_202), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_237), .A2(n_199), .B1(n_195), .B2(n_142), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_231), .A2(n_218), .B1(n_222), .B2(n_220), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_233), .B(n_199), .Y(n_260) );
AOI221xp5_ASAP7_75t_SL g261 ( .A1(n_235), .A2(n_215), .B1(n_213), .B2(n_118), .C(n_111), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_81), .B1(n_99), .B2(n_96), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_244), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_244), .B(n_241), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_244), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_245), .B(n_241), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_250), .A2(n_115), .B(n_234), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_255), .B(n_242), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_245), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_255), .Y(n_270) );
OAI321xp33_ASAP7_75t_L g271 ( .A1(n_243), .A2(n_97), .A3(n_103), .B1(n_79), .B2(n_76), .C(n_73), .Y(n_271) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_261), .A2(n_97), .B(n_75), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_251), .B(n_256), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_243), .A2(n_122), .B1(n_111), .B2(n_112), .C(n_123), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_197), .B(n_198), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_256), .B(n_242), .Y(n_278) );
AOI31xp33_ASAP7_75t_SL g279 ( .A1(n_251), .A2(n_0), .A3(n_1), .B(n_2), .Y(n_279) );
OAI211xp5_ASAP7_75t_L g280 ( .A1(n_253), .A2(n_222), .B(n_220), .C(n_76), .Y(n_280) );
NAND3xp33_ASAP7_75t_L g281 ( .A(n_261), .B(n_73), .C(n_75), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_259), .B(n_220), .Y(n_282) );
OAI31xp33_ASAP7_75t_SL g283 ( .A1(n_253), .A2(n_237), .A3(n_98), .B(n_91), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_269), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_263), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_269), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_270), .B(n_263), .Y(n_288) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_276), .A2(n_246), .B(n_254), .Y(n_289) );
AOI33xp33_ASAP7_75t_L g290 ( .A1(n_274), .A2(n_262), .A3(n_248), .B1(n_249), .B2(n_252), .B3(n_91), .Y(n_290) );
OAI322xp33_ASAP7_75t_L g291 ( .A1(n_273), .A2(n_247), .A3(n_98), .B1(n_122), .B2(n_119), .C1(n_123), .C2(n_112), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_265), .B(n_258), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_273), .A2(n_247), .B1(n_254), .B2(n_222), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_270), .B(n_222), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_280), .A2(n_260), .B1(n_240), .B2(n_257), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_270), .B(n_277), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_278), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_275), .B(n_260), .Y(n_302) );
OAI31xp33_ASAP7_75t_SL g303 ( .A1(n_280), .A2(n_118), .A3(n_119), .B(n_3), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_275), .B(n_234), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
AOI322xp5_ASAP7_75t_L g306 ( .A1(n_274), .A2(n_1), .A3(n_2), .B1(n_5), .B2(n_8), .C1(n_9), .C2(n_11), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_283), .A2(n_240), .B1(n_234), .B2(n_242), .C(n_107), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_268), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_283), .B(n_242), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_288), .B(n_277), .Y(n_314) );
NOR3xp33_ASAP7_75t_L g315 ( .A(n_291), .B(n_271), .C(n_281), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_299), .B(n_277), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_SL g317 ( .A1(n_309), .A2(n_271), .B(n_276), .C(n_139), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g318 ( .A1(n_303), .A2(n_282), .B(n_281), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_301), .B(n_268), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_288), .B(n_311), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_299), .B(n_282), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_313), .B(n_268), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_285), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_305), .B(n_307), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_284), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_309), .A2(n_278), .B1(n_279), .B2(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_287), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_313), .B(n_278), .Y(n_332) );
NAND3xp33_ASAP7_75t_SL g333 ( .A(n_306), .B(n_279), .C(n_12), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_301), .B(n_5), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_300), .B(n_272), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_288), .B(n_272), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_295), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_293), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_302), .B(n_12), .Y(n_343) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_295), .B(n_292), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_308), .B(n_310), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_308), .Y(n_346) );
NOR2xp67_ASAP7_75t_SL g347 ( .A(n_303), .B(n_272), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_292), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_311), .B(n_272), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_300), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_293), .B(n_267), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_286), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_322), .B(n_294), .Y(n_355) );
OAI21xp33_ASAP7_75t_SL g356 ( .A1(n_319), .A2(n_306), .B(n_294), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_286), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_346), .B(n_304), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_335), .A2(n_334), .B1(n_318), .B2(n_343), .C(n_329), .Y(n_360) );
OAI21x1_ASAP7_75t_SL g361 ( .A1(n_344), .A2(n_297), .B(n_304), .Y(n_361) );
XOR2x2_ASAP7_75t_L g362 ( .A(n_333), .B(n_296), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_346), .B(n_297), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_348), .B(n_289), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_341), .B(n_289), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_331), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_348), .B(n_289), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_332), .A2(n_298), .B1(n_290), .B2(n_291), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_332), .A2(n_298), .B1(n_234), .B2(n_107), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_340), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_327), .B(n_13), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_317), .A2(n_289), .B(n_267), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_341), .A2(n_107), .B1(n_15), .B2(n_16), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_314), .B(n_14), .Y(n_377) );
OAI221xp5_ASAP7_75t_SL g378 ( .A1(n_316), .A2(n_14), .B1(n_16), .B2(n_17), .C(n_18), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_315), .A2(n_17), .B(n_18), .C(n_19), .Y(n_379) );
OAI32xp33_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_20), .A3(n_21), .B1(n_22), .B2(n_24), .Y(n_380) );
OAI221xp5_ASAP7_75t_SL g381 ( .A1(n_316), .A2(n_20), .B1(n_21), .B2(n_24), .C(n_25), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_345), .B(n_26), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_314), .B(n_26), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_342), .A2(n_198), .B(n_197), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_323), .B(n_144), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_347), .A2(n_198), .B(n_197), .C(n_32), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_323), .B(n_144), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_324), .B(n_28), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_341), .A2(n_198), .B1(n_156), .B2(n_155), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_351), .B(n_144), .Y(n_394) );
OAI321xp33_ASAP7_75t_L g395 ( .A1(n_338), .A2(n_140), .A3(n_139), .B1(n_131), .B2(n_132), .C(n_155), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_350), .B(n_29), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_325), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_353), .A2(n_140), .B(n_139), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_386), .B(n_354), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_357), .B(n_353), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_355), .B(n_354), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_385), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_368), .B(n_337), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_387), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_393), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_377), .B(n_337), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_373), .B(n_326), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_363), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_360), .B(n_336), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_356), .A2(n_326), .B1(n_325), .B2(n_336), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_367), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_359), .B(n_139), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_388), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_365), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_364), .B(n_131), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_362), .A2(n_131), .B1(n_156), .B2(n_132), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_371), .A2(n_156), .B1(n_131), .B2(n_132), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
AOI211xp5_ASAP7_75t_SL g421 ( .A1(n_378), .A2(n_33), .B(n_36), .C(n_37), .Y(n_421) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_381), .A2(n_38), .B(n_39), .C(n_40), .Y(n_422) );
NOR4xp25_ASAP7_75t_SL g423 ( .A(n_379), .B(n_43), .C(n_44), .D(n_45), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_383), .B(n_46), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_368), .B(n_47), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_370), .B(n_48), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_390), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_392), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_374), .B(n_49), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g434 ( .A1(n_379), .A2(n_51), .B(n_52), .C(n_54), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_411), .Y(n_435) );
XNOR2x1_ASAP7_75t_L g436 ( .A(n_410), .B(n_372), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_409), .A2(n_374), .B1(n_380), .B2(n_382), .C(n_391), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_408), .B(n_396), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_406), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_412), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_401), .B(n_394), .Y(n_441) );
OAI322xp33_ASAP7_75t_L g442 ( .A1(n_415), .A2(n_391), .A3(n_396), .B1(n_375), .B2(n_376), .C1(n_384), .C2(n_389), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_432), .A2(n_376), .B1(n_389), .B2(n_398), .Y(n_443) );
NOR3xp33_ASAP7_75t_SL g444 ( .A(n_419), .B(n_395), .C(n_58), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_421), .A2(n_57), .B(n_59), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_414), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
AOI221x1_ASAP7_75t_L g448 ( .A1(n_429), .A2(n_61), .B1(n_62), .B2(n_63), .C(n_64), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_434), .A2(n_68), .B(n_71), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_404), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_433), .A2(n_418), .B(n_424), .Y(n_451) );
NAND4xp75_ASAP7_75t_L g452 ( .A(n_428), .B(n_430), .C(n_431), .D(n_403), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_422), .A2(n_428), .B(n_405), .C(n_430), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_399), .B(n_416), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_453), .A2(n_407), .B(n_423), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_436), .A2(n_400), .B1(n_427), .B2(n_425), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_453), .A2(n_427), .B(n_402), .C(n_426), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g459 ( .A1(n_436), .A2(n_417), .B(n_413), .Y(n_459) );
NOR2xp33_ASAP7_75t_R g460 ( .A(n_446), .B(n_417), .Y(n_460) );
NAND2x1_ASAP7_75t_SL g461 ( .A(n_443), .B(n_426), .Y(n_461) );
AOI21xp33_ASAP7_75t_SL g462 ( .A1(n_445), .A2(n_402), .B(n_438), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_444), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_439), .B(n_435), .Y(n_464) );
OAI322xp33_ASAP7_75t_L g465 ( .A1(n_455), .A2(n_441), .A3(n_440), .B1(n_454), .B2(n_450), .C1(n_447), .C2(n_449), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_455), .A2(n_437), .B1(n_442), .B2(n_451), .C(n_444), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_452), .B(n_448), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_436), .A2(n_409), .B1(n_410), .B2(n_452), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_446), .B(n_415), .Y(n_469) );
OAI211xp5_ASAP7_75t_L g470 ( .A1(n_437), .A2(n_356), .B(n_410), .C(n_453), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_460), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_463), .A2(n_466), .B1(n_468), .B2(n_459), .Y(n_472) );
NAND3xp33_ASAP7_75t_SL g473 ( .A(n_463), .B(n_470), .C(n_458), .Y(n_473) );
NAND3xp33_ASAP7_75t_SL g474 ( .A(n_458), .B(n_467), .C(n_456), .Y(n_474) );
NOR4xp25_ASAP7_75t_L g475 ( .A(n_474), .B(n_473), .C(n_472), .D(n_471), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_471), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_471), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_476), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_477), .B(n_469), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_478), .B(n_464), .Y(n_480) );
AOI22xp5_ASAP7_75t_SL g481 ( .A1(n_480), .A2(n_475), .B1(n_479), .B2(n_461), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_481), .A2(n_480), .B1(n_465), .B2(n_462), .C(n_457), .Y(n_482) );
endmodule