module fake_jpeg_26791_n_219 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_42),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_17),
.B1(n_34),
.B2(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_22),
.C(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_65),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_18),
.B1(n_24),
.B2(n_57),
.Y(n_78)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_17),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_60),
.Y(n_85)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_25),
.B1(n_23),
.B2(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_26),
.B1(n_34),
.B2(n_21),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_0),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_36),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_19),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_51),
.B1(n_66),
.B2(n_62),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_31),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_89),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_36),
.B1(n_35),
.B2(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_67),
.B1(n_55),
.B2(n_54),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_27),
.C(n_19),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_14),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_98),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_3),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_21),
.B(n_20),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_18),
.B1(n_24),
.B2(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_106),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_107),
.B1(n_76),
.B2(n_70),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_61),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_86),
.B(n_91),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_120),
.B(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_77),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_27),
.C(n_29),
.Y(n_114)
);

OR2x4_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_27),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_88),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_32),
.A3(n_29),
.B1(n_27),
.B2(n_53),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_116),
.C(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_85),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_20),
.B(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_85),
.B(n_20),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_123),
.B(n_124),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_87),
.C(n_81),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_90),
.C(n_97),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_138),
.B(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_76),
.B1(n_70),
.B2(n_67),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_136),
.B1(n_140),
.B2(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_105),
.B1(n_114),
.B2(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_53),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_77),
.C(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_76),
.B1(n_96),
.B2(n_55),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_143),
.B(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_162),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_99),
.B1(n_101),
.B2(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_153),
.B1(n_129),
.B2(n_108),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_154),
.C(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_140),
.B1(n_134),
.B2(n_136),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_99),
.C(n_102),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_110),
.B(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_125),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_171),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_156),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_172),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_126),
.B1(n_128),
.B2(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_170),
.B1(n_179),
.B2(n_180),
.Y(n_188)
);

AOI321xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_122),
.A3(n_100),
.B1(n_115),
.B2(n_118),
.C(n_112),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_122),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_29),
.B(n_32),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_178),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_100),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_177),
.B(n_148),
.Y(n_185)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_152),
.B1(n_149),
.B2(n_151),
.C(n_163),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_118),
.B1(n_112),
.B2(n_115),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_96),
.B1(n_94),
.B2(n_54),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_84),
.C(n_32),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_168),
.C(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_160),
.B1(n_159),
.B2(n_16),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_180),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_6),
.B(n_7),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_12),
.B(n_13),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_15),
.C(n_7),
.Y(n_190)
);

OAI321xp33_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_12),
.A3(n_172),
.B1(n_189),
.B2(n_192),
.C(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_10),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_11),
.CI(n_12),
.CON(n_193),
.SN(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_181),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_198),
.B(n_202),
.Y(n_205)
);

OAI31xp33_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_193),
.A3(n_190),
.B(n_182),
.Y(n_203)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_185),
.B1(n_188),
.B2(n_183),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_196),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_205),
.C(n_209),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_194),
.CI(n_195),
.CON(n_211),
.SN(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_198),
.B(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_211),
.B(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_218),
.B(n_216),
.Y(n_219)
);


endmodule