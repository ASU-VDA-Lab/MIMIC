module real_jpeg_30633_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_650;
wire n_250;
wire n_254;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_686;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_0),
.Y(n_139)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_0),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_0),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g541 ( 
.A(n_0),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_1),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_1),
.A2(n_227),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_1),
.A2(n_227),
.B1(n_257),
.B2(n_261),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_1),
.A2(n_227),
.B1(n_412),
.B2(n_415),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_153),
.B1(n_155),
.B2(n_158),
.Y(n_152)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_2),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_2),
.A2(n_158),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_2),
.A2(n_158),
.B1(n_173),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_2),
.A2(n_158),
.B1(n_402),
.B2(n_404),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_112),
.B1(n_118),
.B2(n_122),
.Y(n_111)
);

INVx2_ASAP7_75t_R g122 ( 
.A(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_4),
.A2(n_122),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g303 ( 
.A1(n_4),
.A2(n_122),
.B1(n_304),
.B2(n_306),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_4),
.A2(n_122),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_5),
.A2(n_372),
.B1(n_375),
.B2(n_379),
.Y(n_371)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_5),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_5),
.A2(n_379),
.B1(n_466),
.B2(n_469),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_5),
.A2(n_379),
.B1(n_534),
.B2(n_536),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_5),
.A2(n_379),
.B1(n_609),
.B2(n_611),
.Y(n_608)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_6),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_7),
.A2(n_342),
.B1(n_343),
.B2(n_345),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_7),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_7),
.A2(n_342),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_7),
.A2(n_342),
.B1(n_527),
.B2(n_530),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_7),
.A2(n_342),
.B1(n_590),
.B2(n_591),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_8),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_8),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_8),
.A2(n_165),
.B1(n_361),
.B2(n_364),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_8),
.A2(n_165),
.B1(n_473),
.B2(n_475),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_8),
.A2(n_165),
.B1(n_404),
.B2(n_603),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_11),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_11),
.Y(n_416)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_11),
.Y(n_560)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_12),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_13),
.B(n_687),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_14),
.A2(n_348),
.B(n_350),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_14),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_14),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_14),
.A2(n_136),
.B1(n_266),
.B2(n_526),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_14),
.B(n_221),
.Y(n_605)
);

OAI32xp33_ASAP7_75t_L g622 ( 
.A1(n_14),
.A2(n_198),
.A3(n_623),
.B1(n_626),
.B2(n_627),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_14),
.A2(n_418),
.B1(n_637),
.B2(n_640),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_15),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

INVx2_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_15),
.A2(n_285),
.B1(n_381),
.B2(n_386),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_15),
.A2(n_285),
.B1(n_556),
.B2(n_561),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_15),
.A2(n_285),
.B1(n_644),
.B2(n_647),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_16),
.A2(n_68),
.B1(n_72),
.B2(n_76),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_16),
.A2(n_76),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_16),
.A2(n_76),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_16),
.A2(n_76),
.B1(n_184),
.B2(n_210),
.Y(n_311)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_17),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_17),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_17),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_18),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_18),
.A2(n_59),
.B1(n_127),
.B2(n_132),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_18),
.A2(n_59),
.B1(n_210),
.B2(n_214),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_18),
.A2(n_59),
.B1(n_146),
.B2(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_19),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_19),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_23),
.B(n_686),
.Y(n_20)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_81),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_80),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_78),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_26),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_26),
.B(n_332),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_27),
.B(n_79),
.Y(n_80)
);

NAND4xp25_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_57),
.C(n_66),
.D(n_77),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_56),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_29),
.A2(n_56),
.B(n_67),
.Y(n_79)
);

OAI22x1_ASAP7_75t_SL g279 ( 
.A1(n_29),
.A2(n_56),
.B1(n_280),
.B2(n_289),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_29),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_29),
.A2(n_56),
.B1(n_341),
.B2(n_347),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_29),
.A2(n_56),
.B1(n_280),
.B2(n_465),
.Y(n_488)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_30),
.B(n_161),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_30),
.A2(n_152),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_30),
.A2(n_238),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_32),
.Y(n_197)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_33),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_34),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_34),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_34),
.Y(n_385)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_35),
.Y(n_430)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_36),
.Y(n_427)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_37),
.Y(n_387)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_37),
.Y(n_423)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_38),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_38),
.Y(n_199)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_46),
.Y(n_164)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_46),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_46),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_50),
.Y(n_157)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_50),
.Y(n_468)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_51),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_56),
.Y(n_159)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_56),
.Y(n_238)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_56),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_56),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g417 ( 
.A(n_56),
.B(n_418),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_58),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_75),
.Y(n_344)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_75),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_333),
.B(n_679),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_313),
.C(n_331),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_290),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_246),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_85),
.B(n_246),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_222),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_167),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_87),
.B(n_293),
.C(n_295),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_135),
.B(n_148),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_88),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_135),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_89),
.A2(n_135),
.B1(n_251),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_89),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_111),
.B1(n_123),
.B2(n_126),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_90),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_90),
.A2(n_111),
.B1(n_123),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_90),
.A2(n_171),
.B1(n_356),
.B2(n_360),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_90),
.A2(n_171),
.B1(n_256),
.B2(n_356),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_90),
.A2(n_171),
.B1(n_607),
.B2(n_608),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_90),
.A2(n_660),
.B(n_661),
.Y(n_659)
);

AO21x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_99),
.B(n_103),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_96),
.Y(n_359)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_98),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_99),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_105),
.Y(n_403)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_105),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_105),
.Y(n_582)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_106),
.Y(n_414)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_115),
.Y(n_590)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_117),
.Y(n_588)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_120),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_121),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_124),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_124),
.A2(n_235),
.B1(n_643),
.B2(n_650),
.Y(n_642)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_131),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_131),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_131),
.Y(n_610)
);

BUFx6f_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_135),
.A2(n_149),
.B1(n_150),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_140),
.B(n_145),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_136),
.A2(n_145),
.B1(n_263),
.B2(n_266),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_136),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_136),
.A2(n_263),
.B1(n_438),
.B2(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_136),
.A2(n_526),
.B1(n_533),
.B2(n_540),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_136),
.A2(n_555),
.B1(n_563),
.B2(n_601),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_139),
.Y(n_548)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_144),
.Y(n_456)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_161),
.Y(n_289)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_167),
.A2(n_168),
.B1(n_237),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_180),
.B2(n_181),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_169),
.B(n_181),
.C(n_294),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_169),
.A2(n_170),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_170),
.B(n_317),
.C(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_171),
.B(n_418),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_171),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_175),
.Y(n_592)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_179),
.Y(n_629)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_179),
.Y(n_649)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_191),
.B1(n_209),
.B2(n_220),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_221),
.B1(n_226),
.B2(n_232),
.Y(n_225)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_189),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_191),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_191),
.A2(n_209),
.B1(n_220),
.B2(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_191),
.A2(n_220),
.B1(n_371),
.B2(n_380),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_191),
.A2(n_220),
.B1(n_371),
.B2(n_390),
.Y(n_389)
);

OA22x2_ASAP7_75t_L g471 ( 
.A1(n_191),
.A2(n_220),
.B1(n_380),
.B2(n_472),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_191),
.A2(n_220),
.B1(n_271),
.B2(n_472),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_191),
.A2(n_220),
.B1(n_390),
.B2(n_636),
.Y(n_635)
);

AO21x2_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_198),
.B(n_202),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_216),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_218),
.Y(n_393)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_218),
.Y(n_474)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_221),
.A2(n_226),
.B1(n_232),
.B2(n_270),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_221),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.Y(n_222)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_225),
.B(n_233),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_233),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_235),
.A2(n_585),
.B1(n_589),
.B2(n_593),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_237),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_239),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_243),
.Y(n_469)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.C(n_253),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_249),
.B(n_252),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_253),
.B(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_268),
.C(n_278),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_254),
.B(n_493),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_262),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_255),
.B(n_262),
.Y(n_510)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_269),
.B(n_279),
.Y(n_493)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_274),
.Y(n_397)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_274),
.Y(n_433)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

BUFx4f_ASAP7_75t_SL g349 ( 
.A(n_288),
.Y(n_349)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_291),
.A2(n_682),
.B(n_683),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_292),
.B(n_296),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_297),
.C(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_309),
.Y(n_298)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_309),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_303),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_304),
.A2(n_421),
.A3(n_424),
.B1(n_428),
.B2(n_434),
.Y(n_420)
);

OAI32xp33_ASAP7_75t_L g447 ( 
.A1(n_304),
.A2(n_421),
.A3(n_424),
.B1(n_428),
.B2(n_434),
.Y(n_447)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_314),
.A2(n_681),
.B(n_684),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_329),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_315),
.B(n_329),
.Y(n_684)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_320),
.C(n_328),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_323),
.B1(n_327),
.B2(n_328),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_331),
.A2(n_680),
.B(n_685),
.Y(n_679)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_518),
.B(n_674),
.Y(n_334)
);

NAND4xp25_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_479),
.C(n_499),
.D(n_512),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_449),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_337),
.B(n_449),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_388),
.C(n_419),
.Y(n_337)
);

XOR2x2_ASAP7_75t_L g670 ( 
.A(n_338),
.B(n_671),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_354),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g458 ( 
.A(n_340),
.B(n_355),
.C(n_370),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_341),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_370),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g662 ( 
.A(n_360),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_368),
.Y(n_580)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_374),
.Y(n_639)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_378),
.Y(n_641)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_388),
.B(n_419),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_398),
.C(n_417),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_389),
.B(n_666),
.Y(n_665)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_398),
.A2(n_399),
.B1(n_417),
.B2(n_667),
.Y(n_666)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_408),
.B2(n_411),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_400),
.A2(n_411),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_400),
.A2(n_553),
.B1(n_554),
.B2(n_562),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_400),
.A2(n_401),
.B1(n_602),
.B2(n_631),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_407),
.Y(n_539)
);

BUFx2_ASAP7_75t_R g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_410),
.Y(n_436)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_416),
.Y(n_572)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_417),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_418),
.B(n_547),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_418),
.B(n_579),
.Y(n_578)
);

OAI21xp33_ASAP7_75t_SL g585 ( 
.A1(n_418),
.A2(n_578),
.B(n_586),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_418),
.B(n_628),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_435),
.B1(n_446),
.B2(n_448),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_420),
.B(n_448),
.Y(n_478)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_431),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_435),
.Y(n_448)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_441),
.Y(n_603)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_459),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_458),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_451),
.B(n_459),
.C(n_501),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_457),
.Y(n_486)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_478),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_462),
.B1(n_470),
.B2(n_471),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_478),
.C(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_471),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

A2O1A1O1Ixp25_ASAP7_75t_L g674 ( 
.A1(n_479),
.A2(n_512),
.B(n_675),
.C(n_677),
.D(n_678),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_497),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_480),
.B(n_497),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_491),
.B(n_494),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_484),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_517),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_487),
.C(n_489),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_485),
.A2(n_486),
.B1(n_507),
.B2(n_511),
.Y(n_515)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_510),
.Y(n_509)
);

AO22x1_ASAP7_75t_L g507 ( 
.A1(n_487),
.A2(n_488),
.B1(n_489),
.B2(n_490),
.Y(n_507)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_496),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_500),
.B(n_502),
.C(n_676),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_514),
.C(n_515),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_508),
.B1(n_509),
.B2(n_511),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_510),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_513),
.B(n_516),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_669),
.B(n_673),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_654),
.B(n_668),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_618),
.B(n_653),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_597),
.B(n_617),
.Y(n_521)
);

AOI22x1_ASAP7_75t_SL g522 ( 
.A1(n_523),
.A2(n_551),
.B1(n_595),
.B2(n_596),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_524),
.A2(n_543),
.B(n_550),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_542),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_525),
.B(n_542),
.Y(n_550)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_533),
.Y(n_553)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_540),
.Y(n_631)
);

INVx4_ASAP7_75t_SL g540 ( 
.A(n_541),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_544),
.B(n_545),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_549),
.Y(n_545)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_566),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_552),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_567),
.A2(n_568),
.B1(n_584),
.B2(n_594),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_567),
.B(n_594),
.Y(n_598)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_569),
.A2(n_577),
.B1(n_581),
.B2(n_583),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_570),
.B(n_573),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_571),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_584),
.Y(n_594)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_588),
.Y(n_626)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_588),
.Y(n_646)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_589),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_593),
.B(n_662),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_598),
.B(n_599),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_598),
.B(n_599),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_604),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_600),
.B(n_606),
.C(n_615),
.Y(n_619)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_605),
.A2(n_606),
.B1(n_615),
.B2(n_616),
.Y(n_604)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_605),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_606),
.Y(n_616)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_608),
.Y(n_650)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_619),
.B(n_620),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_SL g653 ( 
.A(n_619),
.B(n_620),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_621),
.B(n_634),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_621),
.B(n_642),
.C(n_652),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_622),
.A2(n_630),
.B1(n_632),
.B2(n_633),
.Y(n_621)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_622),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_622),
.B(n_633),
.Y(n_664)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_630),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_635),
.A2(n_642),
.B1(n_651),
.B2(n_652),
.Y(n_634)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_635),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_638),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_642),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_643),
.Y(n_660)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_646),
.Y(n_645)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_655),
.B(n_656),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_655),
.B(n_656),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_SL g656 ( 
.A(n_657),
.B(n_665),
.Y(n_656)
);

OA22x2_ASAP7_75t_L g657 ( 
.A1(n_658),
.A2(n_659),
.B1(n_663),
.B2(n_664),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_659),
.B(n_663),
.C(n_665),
.Y(n_672)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_670),
.B(n_672),
.Y(n_669)
);

NOR2x1_ASAP7_75t_L g673 ( 
.A(n_670),
.B(n_672),
.Y(n_673)
);


endmodule