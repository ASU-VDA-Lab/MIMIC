module fake_jpeg_7357_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_47),
.Y(n_52)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_65)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_58),
.Y(n_106)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_68),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_63),
.B1(n_28),
.B2(n_19),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_70),
.B1(n_44),
.B2(n_35),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_11),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_40),
.Y(n_85)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_77),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_91),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_0),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_113),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_19),
.B1(n_28),
.B2(n_45),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_45),
.B1(n_30),
.B2(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_34),
.B1(n_27),
.B2(n_31),
.Y(n_140)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_93),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_16),
.B1(n_25),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_103),
.Y(n_120)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_16),
.B1(n_47),
.B2(n_17),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_44),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_111),
.B1(n_66),
.B2(n_74),
.Y(n_122)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_132),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_106),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_119),
.A2(n_141),
.B(n_0),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_139),
.B1(n_111),
.B2(n_97),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_137),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_42),
.B(n_39),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_51),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_42),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_42),
.C(n_39),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_66),
.B1(n_74),
.B2(n_35),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_94),
.B1(n_97),
.B2(n_75),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_109),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_151),
.B1(n_162),
.B2(n_170),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_82),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_149),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_148),
.A2(n_88),
.B1(n_128),
.B2(n_124),
.Y(n_210)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_111),
.B1(n_92),
.B2(n_79),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_87),
.B1(n_113),
.B2(n_79),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_137),
.B(n_125),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_105),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_154),
.A2(n_164),
.B(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_160),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_159),
.B(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_96),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_163),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_78),
.B1(n_61),
.B2(n_72),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_80),
.Y(n_163)
);

BUFx12f_ASAP7_75t_SL g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_132),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_165),
.A2(n_177),
.B1(n_133),
.B2(n_128),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_112),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_173),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_126),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_83),
.B1(n_77),
.B2(n_78),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_122),
.B1(n_125),
.B2(n_133),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_123),
.B(n_15),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_171),
.B(n_172),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_107),
.C(n_26),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_23),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_88),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_31),
.B1(n_26),
.B2(n_34),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_181),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_205),
.B(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_185),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_123),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_147),
.C(n_173),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_203),
.C(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_200),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_141),
.Y(n_200)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_64),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_131),
.C(n_120),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_141),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_145),
.B(n_115),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_109),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_22),
.B1(n_23),
.B2(n_4),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_226),
.C(n_180),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_170),
.B1(n_154),
.B2(n_155),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_222),
.B1(n_228),
.B2(n_195),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_217),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_114),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_114),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_223),
.A3(n_201),
.B1(n_207),
.B2(n_205),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_140),
.C(n_145),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_220),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_176),
.B1(n_161),
.B2(n_149),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_176),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_231),
.B(n_185),
.C(n_187),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_22),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_227),
.B(n_238),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_102),
.B1(n_116),
.B2(n_27),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_116),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_233),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_232),
.B1(n_209),
.B2(n_190),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_102),
.B1(n_23),
.B2(n_22),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_22),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_237),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_8),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_192),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_247),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_256),
.B1(n_184),
.B2(n_182),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_182),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_259),
.B1(n_257),
.B2(n_255),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_190),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_218),
.B(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_207),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_237),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_219),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_213),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_264),
.B(n_270),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_220),
.B1(n_178),
.B2(n_200),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_247),
.B1(n_249),
.B2(n_239),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_211),
.C(n_212),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_271),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_252),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_216),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_183),
.C(n_181),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_215),
.C(n_186),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_188),
.C(n_3),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_280),
.Y(n_295)
);

FAx1_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_1),
.CI(n_3),
.CON(n_280),
.SN(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_242),
.B1(n_254),
.B2(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_256),
.B1(n_240),
.B2(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_285),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_240),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_240),
.B(n_11),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_280),
.C(n_279),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_267),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_12),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_276),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_262),
.C(n_273),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_303),
.B(n_296),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_286),
.C(n_288),
.Y(n_303)
);

AOI221xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_280),
.B1(n_271),
.B2(n_7),
.C(n_10),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_13),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_286),
.C(n_287),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_12),
.C(n_6),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_15),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_7),
.B(n_11),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_295),
.B(n_285),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_307),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_319),
.B(n_300),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_7),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_13),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_321),
.C(n_312),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_301),
.B(n_299),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_304),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_313),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_311),
.C(n_317),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_330),
.B(n_325),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_SL g333 ( 
.A(n_331),
.B(n_332),
.C(n_328),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_324),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_14),
.B(n_5),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_5),
.Y(n_336)
);


endmodule