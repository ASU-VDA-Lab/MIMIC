module fake_jpeg_18232_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_7),
.B1(n_6),
.B2(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_18),
.Y(n_23)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_2),
.B1(n_4),
.B2(n_7),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_17),
.B(n_14),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_17),
.B(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_23),
.C(n_20),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_20),
.B(n_19),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_12),
.B(n_22),
.Y(n_31)
);

NAND4xp25_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_12),
.C(n_22),
.D(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_16),
.Y(n_33)
);


endmodule