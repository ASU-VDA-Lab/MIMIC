module fake_jpeg_22602_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx14_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_12),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_41),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_38),
.B1(n_32),
.B2(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_16),
.B1(n_33),
.B2(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_15),
.B(n_10),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_2),
.B(n_4),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_38),
.B1(n_36),
.B2(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_36),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_54),
.C(n_53),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

FAx1_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_46),
.CI(n_7),
.CON(n_68),
.SN(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_64),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_69),
.B(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_70),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_61),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_60),
.C(n_76),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_65),
.Y(n_79)
);


endmodule