module fake_jpeg_2970_n_233 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_233);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_8),
.B(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_52),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_86),
.Y(n_87)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_0),
.Y(n_86)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_66),
.B1(n_58),
.B2(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_57),
.B1(n_54),
.B2(n_67),
.Y(n_111)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_66),
.B1(n_58),
.B2(n_74),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_54),
.B(n_75),
.Y(n_112)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_71),
.B1(n_63),
.B2(n_64),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_52),
.B1(n_75),
.B2(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_85),
.B1(n_64),
.B2(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_110),
.B1(n_114),
.B2(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_56),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_112),
.C(n_60),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_132)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_2),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_96),
.B1(n_94),
.B2(n_90),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_76),
.B1(n_70),
.B2(n_68),
.Y(n_130)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_90),
.B1(n_100),
.B2(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_65),
.B1(n_73),
.B2(n_61),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_67),
.C(n_53),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_119),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_57),
.B1(n_73),
.B2(n_61),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_57),
.B1(n_60),
.B2(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_72),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_128),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_62),
.B(n_91),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_109),
.B(n_116),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_88),
.B1(n_93),
.B2(n_65),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_140),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_129),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_1),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_43),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_3),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_4),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_103),
.B1(n_120),
.B2(n_117),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_147),
.B1(n_153),
.B2(n_17),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_158),
.B(n_133),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_104),
.B1(n_116),
.B2(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_155),
.B1(n_159),
.B2(n_165),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_51),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_154),
.C(n_22),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_49),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_161),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_162),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_41),
.B(n_40),
.C(n_39),
.D(n_37),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_14),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_16),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_133),
.A3(n_139),
.B1(n_141),
.B2(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_121),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_31),
.B(n_18),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_183),
.B(n_25),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_17),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_29),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_186),
.C(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_19),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_143),
.B(n_158),
.C(n_154),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_19),
.B(n_21),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_22),
.C(n_23),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_24),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_25),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_148),
.B1(n_26),
.B2(n_27),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_176),
.B(n_183),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_26),
.C(n_27),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_178),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_184),
.C(n_211),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_177),
.B1(n_182),
.B2(n_179),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_185),
.B1(n_169),
.B2(n_187),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_210),
.B(n_199),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_182),
.B(n_171),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_213),
.B(n_192),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_189),
.B(n_168),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_193),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_186),
.C(n_203),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_219),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_192),
.B1(n_206),
.B2(n_203),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_202),
.B1(n_201),
.B2(n_200),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_213),
.B1(n_207),
.B2(n_195),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_223),
.B1(n_218),
.B2(n_215),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_214),
.B(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.C(n_224),
.Y(n_228)
);

OAI21x1_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_221),
.B(n_222),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_28),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_28),
.Y(n_233)
);


endmodule