module fake_jpeg_31531_n_26 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_26;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_9),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_7),
.Y(n_13)
);

OAI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_0),
.A2(n_7),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_0),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_1),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_11),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_12),
.B1(n_8),
.B2(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

MAJx2_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_5),
.C(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_12),
.B1(n_3),
.B2(n_5),
.Y(n_21)
);

NOR2xp67_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_20),
.B(n_22),
.Y(n_25)
);

OAI211xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_20),
.B(n_24),
.C(n_6),
.Y(n_26)
);


endmodule