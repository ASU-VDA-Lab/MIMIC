module fake_netlist_1_647_n_27 (n_3, n_1, n_2, n_0, n_27);
input n_3;
input n_1;
input n_2;
input n_0;
output n_27;
wire n_20;
wire n_5;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_4;
wire n_7;
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_0), .Y(n_5) );
CKINVDCx20_ASAP7_75t_R g6 ( .A(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_2), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_4), .B(n_0), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_5), .B(n_1), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g11 ( .A(n_4), .B(n_1), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_7), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_10), .B(n_7), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_6), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_13), .B(n_11), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_18), .B(n_14), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_14), .B1(n_6), .B2(n_8), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
NAND4xp25_ASAP7_75t_L g22 ( .A(n_20), .B(n_16), .C(n_12), .D(n_17), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_16), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_23), .B1(n_24), .B2(n_3), .Y(n_27) );
endmodule