module fake_aes_12038_n_583 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_583);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_583;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g74 ( .A(n_63), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_36), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_60), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_52), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_13), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_28), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_9), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_37), .Y(n_81) );
INVxp67_ASAP7_75t_L g82 ( .A(n_18), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_11), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_2), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_50), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_61), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_46), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_24), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_49), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_3), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_5), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_55), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_66), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_20), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_35), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_9), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_25), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_32), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_57), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_26), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_39), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_17), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_27), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_69), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_5), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_42), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_79), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_80), .B(n_92), .Y(n_122) );
BUFx8_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_79), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_91), .B(n_0), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_79), .B(n_1), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_116), .B(n_1), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_117), .B(n_3), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_76), .B(n_4), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_86), .B(n_96), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_81), .B(n_4), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_94), .B(n_6), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_110), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_110), .B(n_6), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_112), .B(n_7), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_114), .B(n_7), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_114), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g146 ( .A1(n_99), .A2(n_8), .B1(n_10), .B2(n_12), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_98), .Y(n_152) );
BUFx8_ASAP7_75t_L g153 ( .A(n_102), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_87), .B(n_8), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_84), .B(n_10), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_84), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_104), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_124), .B(n_105), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_124), .B(n_107), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_155), .Y(n_164) );
OAI22xp33_ASAP7_75t_SL g165 ( .A1(n_154), .A2(n_118), .B1(n_83), .B2(n_101), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_132), .B(n_111), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_157), .B(n_106), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_132), .B(n_108), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_142), .B(n_95), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_126), .B(n_101), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_156), .B(n_106), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_122), .A2(n_118), .B1(n_75), .B2(n_103), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_156), .B(n_100), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_122), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_149), .B(n_88), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_123), .B(n_109), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_155), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_120), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_120), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_142), .B(n_82), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_128), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_149), .B(n_113), .Y(n_188) );
BUFx4_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_156), .B(n_113), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_131), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_150), .B(n_109), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_156), .B(n_77), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_150), .A2(n_99), .B1(n_103), .B2(n_75), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
HB1xp67_ASAP7_75t_SL g202 ( .A(n_123), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_130), .B(n_77), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_152), .B(n_12), .Y(n_204) );
INVxp67_ASAP7_75t_L g205 ( .A(n_123), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
OAI22xp5_ASAP7_75t_SL g207 ( .A1(n_146), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_153), .B(n_53), .Y(n_208) );
BUFx10_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_152), .B(n_16), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_155), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_212), .B(n_153), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_172), .Y(n_216) );
BUFx12f_ASAP7_75t_L g217 ( .A(n_209), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_213), .B(n_158), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_204), .B(n_141), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_171), .A2(n_158), .B1(n_134), .B2(n_148), .Y(n_221) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_205), .B(n_151), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_209), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_172), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_167), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_204), .A2(n_136), .B1(n_148), .B2(n_151), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_193), .B(n_145), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_167), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_169), .B(n_136), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_190), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_176), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_176), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_192), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_192), .Y(n_236) );
NOR2x1p5_ASAP7_75t_L g237 ( .A(n_189), .B(n_153), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_161), .B(n_145), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_169), .B(n_136), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
INVx4_ASAP7_75t_L g241 ( .A(n_173), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_159), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_160), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_171), .B(n_145), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_203), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_170), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_181), .Y(n_247) );
INVxp33_ASAP7_75t_SL g248 ( .A(n_174), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_186), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_191), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_188), .B(n_136), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_177), .B(n_143), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_SL g255 ( .A1(n_178), .A2(n_135), .B(n_143), .C(n_136), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_180), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_187), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_180), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_187), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_202), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_188), .B(n_136), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_203), .B(n_16), .Y(n_262) );
INVxp33_ASAP7_75t_SL g263 ( .A(n_200), .Y(n_263) );
AND3x2_ASAP7_75t_SL g264 ( .A(n_200), .B(n_136), .C(n_127), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_198), .B(n_129), .Y(n_265) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_210), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
OR2x2_ASAP7_75t_SL g268 ( .A(n_202), .B(n_129), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_206), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_187), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_256), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_251), .A2(n_193), .B(n_199), .Y(n_273) );
O2A1O1Ixp5_ASAP7_75t_L g274 ( .A1(n_255), .A2(n_208), .B(n_166), .C(n_168), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_217), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g277 ( .A1(n_261), .A2(n_166), .B(n_168), .C(n_179), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_217), .Y(n_279) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_265), .A2(n_163), .B(n_162), .Y(n_280) );
BUFx10_ASAP7_75t_L g281 ( .A(n_237), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_260), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_258), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_248), .A2(n_200), .B1(n_165), .B2(n_207), .C(n_178), .Y(n_284) );
INVx3_ASAP7_75t_SL g285 ( .A(n_241), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_241), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_SL g287 ( .A1(n_231), .A2(n_162), .B(n_163), .C(n_205), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_228), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_241), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_218), .B(n_198), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_236), .Y(n_291) );
O2A1O1Ixp5_ASAP7_75t_L g292 ( .A1(n_215), .A2(n_199), .B(n_175), .C(n_184), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_220), .A2(n_173), .B1(n_175), .B2(n_184), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_232), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_254), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_254), .Y(n_298) );
BUFx6f_ASAP7_75t_SL g299 ( .A(n_225), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_254), .Y(n_301) );
AOI21xp5_ASAP7_75t_SL g302 ( .A1(n_266), .A2(n_211), .B(n_183), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_254), .B(n_218), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_232), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_230), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_230), .B(n_214), .Y(n_307) );
NOR2xp33_ASAP7_75t_SL g308 ( .A(n_260), .B(n_173), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_223), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_245), .B(n_164), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_235), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_226), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_248), .A2(n_201), .B1(n_196), .B2(n_182), .C(n_194), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_269), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_242), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_304), .B(n_244), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_316), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_304), .B(n_220), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_316), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
AND2x6_ASAP7_75t_L g323 ( .A(n_286), .B(n_252), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_288), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_284), .A2(n_263), .B1(n_173), .B2(n_253), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_312), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_283), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_312), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_272), .Y(n_335) );
INVx8_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVx4_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_272), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_290), .B(n_221), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_293), .A2(n_227), .B1(n_262), .B2(n_263), .Y(n_340) );
BUFx4f_ASAP7_75t_L g341 ( .A(n_286), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_286), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_313), .A2(n_253), .B1(n_229), .B2(n_262), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_311), .A2(n_222), .B(n_238), .C(n_229), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_343), .A2(n_238), .B1(n_229), .B2(n_292), .C(n_314), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_326), .A2(n_279), .B1(n_282), .B2(n_309), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_340), .A2(n_315), .B1(n_310), .B2(n_303), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_339), .A2(n_315), .B1(n_310), .B2(n_303), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_302), .B1(n_315), .B2(n_309), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_335), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g353 ( .A1(n_344), .A2(n_273), .B(n_302), .C(n_297), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_320), .A2(n_287), .B(n_277), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_337), .B(n_304), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_320), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_318), .A2(n_308), .B1(n_264), .B2(n_304), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_325), .A2(n_306), .B1(n_275), .B2(n_299), .C(n_307), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_320), .A2(n_304), .B1(n_303), .B2(n_223), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_345), .A2(n_304), .B1(n_268), .B2(n_306), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_345), .A2(n_268), .B1(n_280), .B2(n_289), .Y(n_362) );
AOI21x1_ASAP7_75t_L g363 ( .A1(n_325), .A2(n_280), .B(n_243), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_345), .A2(n_289), .B1(n_242), .B2(n_243), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_338), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_321), .A2(n_246), .B1(n_249), .B2(n_250), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_327), .A2(n_246), .B1(n_249), .B2(n_250), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_327), .A2(n_267), .B1(n_307), .B2(n_276), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_337), .B(n_300), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_338), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_319), .A2(n_275), .B(n_264), .C(n_185), .Y(n_371) );
NAND3xp33_ASAP7_75t_L g372 ( .A(n_348), .B(n_274), .C(n_125), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_357), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_363), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_347), .A2(n_331), .B1(n_329), .B2(n_299), .C(n_307), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_351), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_359), .A2(n_319), .B1(n_329), .B2(n_331), .C(n_317), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_350), .A2(n_317), .B1(n_337), .B2(n_333), .C(n_334), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_350), .A2(n_337), .B1(n_333), .B2(n_334), .C(n_322), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_353), .B(n_119), .C(n_121), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_349), .A2(n_336), .B1(n_307), .B2(n_323), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_321), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_356), .B(n_328), .Y(n_386) );
OAI322xp33_ASAP7_75t_L g387 ( .A1(n_352), .A2(n_264), .A3(n_119), .B1(n_125), .B2(n_129), .C1(n_121), .C2(n_324), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_369), .B(n_328), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_370), .B(n_332), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_367), .B(n_332), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_358), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_369), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_360), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_358), .A2(n_336), .B1(n_323), .B2(n_334), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_361), .A2(n_299), .B1(n_324), .B2(n_332), .C(n_267), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_368), .A2(n_336), .B1(n_276), .B2(n_291), .C(n_278), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_371), .B(n_129), .C(n_125), .Y(n_397) );
OAI31xp33_ASAP7_75t_L g398 ( .A1(n_362), .A2(n_322), .A3(n_239), .B(n_291), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_367), .B(n_336), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_322), .B1(n_336), .B2(n_341), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_355), .A2(n_125), .B(n_129), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_366), .B(n_281), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_364), .A2(n_278), .B(n_281), .C(n_342), .Y(n_403) );
OAI31xp33_ASAP7_75t_SL g404 ( .A1(n_400), .A2(n_323), .A3(n_281), .B(n_341), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_385), .B(n_342), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_323), .B1(n_281), .B2(n_341), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_399), .A2(n_323), .B1(n_341), .B2(n_286), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_390), .B(n_323), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_379), .A2(n_323), .B1(n_286), .B2(n_298), .Y(n_409) );
AOI211xp5_ASAP7_75t_SL g410 ( .A1(n_382), .A2(n_298), .B(n_296), .C(n_23), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_389), .B(n_121), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_393), .A2(n_298), .B1(n_296), .B2(n_300), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_389), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_376), .B(n_121), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_386), .B(n_121), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_390), .A2(n_384), .B1(n_381), .B2(n_392), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_378), .B(n_21), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_374), .B(n_119), .Y(n_419) );
OAI33xp33_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_119), .A3(n_30), .B1(n_31), .B2(n_33), .B3(n_38), .Y(n_420) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_380), .A2(n_119), .A3(n_195), .B1(n_296), .B2(n_44), .C1(n_45), .C2(n_47), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_378), .B(n_22), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_375), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_376), .B(n_41), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_392), .B(n_300), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_388), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_388), .B(n_43), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_388), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_391), .B(n_54), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_401), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_394), .B(n_56), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_398), .B(n_58), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_402), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_372), .B(n_195), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_395), .B(n_62), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_396), .B(n_64), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_65), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_385), .B(n_67), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_389), .B(n_68), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_373), .B(n_70), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_375), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_385), .B(n_71), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_385), .B(n_72), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_413), .B(n_73), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_446), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_446), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_427), .Y(n_454) );
NAND5xp2_ASAP7_75t_L g455 ( .A(n_404), .B(n_301), .C(n_219), .D(n_224), .E(n_216), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_430), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_430), .B(n_247), .Y(n_460) );
AND2x4_ASAP7_75t_SL g461 ( .A(n_405), .B(n_301), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_404), .B(n_247), .C(n_271), .D(n_270), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_437), .A2(n_301), .B1(n_219), .B2(n_224), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_408), .B(n_240), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_437), .B(n_216), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_429), .B(n_240), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_428), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
NAND2x2_ASAP7_75t_L g471 ( .A(n_429), .B(n_216), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_405), .B(n_270), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_415), .B(n_233), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_411), .B(n_233), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_411), .B(n_257), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_428), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_425), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_416), .B(n_257), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_418), .B(n_216), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_416), .B(n_259), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_415), .B(n_259), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_419), .B(n_216), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_419), .B(n_219), .Y(n_486) );
AND3x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_219), .C(n_224), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_418), .B(n_224), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_451), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_481), .B(n_423), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_476), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_458), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_485), .B(n_423), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_459), .B(n_423), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_455), .B(n_410), .C(n_406), .D(n_409), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_450), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_469), .B(n_421), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_461), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_480), .A2(n_406), .B1(n_407), .B2(n_434), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_456), .B(n_410), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_457), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_470), .B(n_448), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_458), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_466), .B(n_447), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_479), .A2(n_421), .B(n_442), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_468), .B(n_434), .C(n_440), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_461), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_488), .B(n_432), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_477), .B(n_443), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_478), .B(n_433), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_481), .B(n_442), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_482), .A2(n_440), .B1(n_441), .B2(n_426), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_464), .B(n_412), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_464), .B(n_432), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_472), .B(n_438), .Y(n_519) );
AOI211xp5_ASAP7_75t_L g520 ( .A1(n_462), .A2(n_441), .B(n_420), .C(n_435), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_490), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_499), .Y(n_522) );
OAI21xp5_ASAP7_75t_SL g523 ( .A1(n_498), .A2(n_487), .B(n_463), .Y(n_523) );
XOR2x2_ASAP7_75t_L g524 ( .A(n_494), .B(n_510), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_502), .Y(n_525) );
NAND2xp33_ASAP7_75t_SL g526 ( .A(n_511), .B(n_489), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_498), .A2(n_420), .B(n_465), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_491), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_501), .B(n_449), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_520), .B(n_463), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_493), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_503), .B(n_460), .Y(n_532) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_492), .B(n_471), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_512), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_500), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_503), .B(n_467), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_505), .Y(n_537) );
XOR2x2_ASAP7_75t_L g538 ( .A(n_492), .B(n_474), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_507), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_509), .A2(n_439), .B(n_474), .C(n_473), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_509), .A2(n_473), .B1(n_483), .B2(n_484), .C1(n_486), .C2(n_475), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_518), .Y(n_542) );
AOI21x1_ASAP7_75t_L g543 ( .A1(n_515), .A2(n_484), .B(n_486), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_504), .B(n_234), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_516), .A2(n_234), .B1(n_514), .B2(n_496), .Y(n_545) );
AOI211xp5_ASAP7_75t_SL g546 ( .A1(n_504), .A2(n_234), .B(n_496), .C(n_519), .Y(n_546) );
OAI31xp33_ASAP7_75t_L g547 ( .A1(n_517), .A2(n_234), .A3(n_497), .B(n_506), .Y(n_547) );
XNOR2xp5_ASAP7_75t_L g548 ( .A(n_513), .B(n_508), .Y(n_548) );
OAI211xp5_ASAP7_75t_L g549 ( .A1(n_495), .A2(n_501), .B(n_404), .C(n_498), .Y(n_549) );
OAI22x1_ASAP7_75t_L g550 ( .A1(n_492), .A2(n_494), .B1(n_502), .B2(n_490), .Y(n_550) );
OAI22xp33_ASAP7_75t_SL g551 ( .A1(n_494), .A2(n_476), .B1(n_471), .B2(n_501), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_499), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_499), .A2(n_485), .B1(n_501), .B2(n_263), .C(n_503), .Y(n_553) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_498), .B(n_455), .Y(n_554) );
AO22x2_ASAP7_75t_L g555 ( .A1(n_521), .A2(n_549), .B1(n_525), .B2(n_552), .Y(n_555) );
AOI221x1_ASAP7_75t_L g556 ( .A1(n_551), .A2(n_550), .B1(n_529), .B2(n_527), .C(n_540), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_522), .Y(n_557) );
OAI21xp33_ASAP7_75t_L g558 ( .A1(n_524), .A2(n_554), .B(n_529), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_542), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_539), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_528), .Y(n_561) );
INVxp33_ASAP7_75t_SL g562 ( .A(n_548), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_534), .B(n_541), .Y(n_563) );
AND3x1_ASAP7_75t_L g564 ( .A(n_553), .B(n_524), .C(n_523), .Y(n_564) );
OAI221xp5_ASAP7_75t_R g565 ( .A1(n_564), .A2(n_545), .B1(n_538), .B2(n_532), .C(n_530), .Y(n_565) );
AOI221xp5_ASAP7_75t_SL g566 ( .A1(n_558), .A2(n_530), .B1(n_540), .B2(n_533), .C(n_532), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_556), .A2(n_546), .B(n_533), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_560), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_563), .B(n_544), .C(n_536), .Y(n_569) );
AO22x2_ASAP7_75t_L g570 ( .A1(n_557), .A2(n_531), .B1(n_535), .B2(n_537), .Y(n_570) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_555), .A2(n_536), .B(n_547), .C(n_526), .Y(n_571) );
NAND4xp25_ASAP7_75t_SL g572 ( .A(n_566), .B(n_571), .C(n_567), .D(n_565), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_568), .A2(n_555), .B1(n_562), .B2(n_560), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_569), .B(n_561), .Y(n_574) );
NAND3x1_ASAP7_75t_L g575 ( .A(n_570), .B(n_555), .C(n_543), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_574), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_575), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_576), .B(n_573), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_577), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_578), .B(n_579), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_580), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_581), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_577), .B1(n_572), .B2(n_559), .Y(n_583) );
endmodule