module fake_ariane_59_n_4411 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_478, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_4411);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_478;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_4411;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4030;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_589;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_4342;
wire n_691;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_610;
wire n_4403;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_690;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_4178;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_3765;
wire n_2006;
wire n_4090;
wire n_952;
wire n_864;
wire n_4058;
wire n_2446;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_4363;
wire n_524;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_634;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_4103;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_2873;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_568;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_520;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_945;
wire n_958;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4106;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_500;
wire n_665;
wire n_754;
wire n_4260;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_829;
wire n_1761;
wire n_4148;
wire n_1062;
wire n_3679;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_4038;
wire n_4132;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_953;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_2634;
wire n_3451;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_645;
wire n_2663;
wire n_495;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_821;
wire n_561;
wire n_770;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_507;
wire n_901;
wire n_2782;
wire n_3879;
wire n_569;
wire n_4136;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_787;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_4176;
wire n_1207;
wire n_4124;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_3948;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4147;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3828;
wire n_3975;
wire n_3073;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_4018;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_661;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_3003;
wire n_2874;
wire n_4117;
wire n_533;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_3739;
wire n_3962;
wire n_512;
wire n_1597;
wire n_4082;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_579;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_2956;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_1021;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_570;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_2909;
wire n_1416;
wire n_3554;
wire n_4276;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_575;
wire n_546;
wire n_3472;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_4109;
wire n_3777;
wire n_4108;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_3588;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_3280;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_2216;
wire n_4115;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_652;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_1260;
wire n_930;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_1179;
wire n_4311;
wire n_3284;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_696;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_4378;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_2398;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2930;
wire n_2871;
wire n_3000;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_619;
wire n_967;
wire n_1083;
wire n_3937;
wire n_4130;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_746;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_615;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_3891;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_4410;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_3257;
wire n_650;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3727;
wire n_3700;
wire n_712;
wire n_976;
wire n_3567;
wire n_909;
wire n_4003;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2795;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_799;
wire n_3884;
wire n_1147;
wire n_2829;
wire n_4367;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_965;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_646;
wire n_4254;
wire n_2507;
wire n_4219;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_3661;
wire n_2223;
wire n_836;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_564;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_3179;
wire n_2262;
wire n_2565;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_927;
wire n_1095;
wire n_2980;
wire n_3699;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3971;
wire n_4315;
wire n_2120;
wire n_706;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_4201;
wire n_3711;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_3994;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_4263;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3876;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4089;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_1198;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_4138;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_855;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_1609;
wire n_1053;
wire n_600;
wire n_3118;
wire n_4072;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_4323;
wire n_1899;
wire n_529;
wire n_3039;
wire n_2195;
wire n_3922;
wire n_502;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_3599;
wire n_3618;
wire n_604;
wire n_677;
wire n_3705;
wire n_3983;
wire n_3022;
wire n_703;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_681;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_707;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_3788;
wire n_3939;
wire n_590;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_3542;
wire n_3569;
wire n_2523;
wire n_1945;
wire n_3835;
wire n_3837;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_3819;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_4348;
wire n_688;
wire n_3139;
wire n_636;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_2802;
wire n_1104;
wire n_1963;
wire n_986;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_887;
wire n_729;
wire n_3403;
wire n_4261;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_627;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_957;
wire n_1402;
wire n_1242;
wire n_3957;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_877;
wire n_3995;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_527;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_3896;
wire n_4049;
wire n_4067;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_551;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_4387;
wire n_1919;
wire n_710;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_560;
wire n_890;
wire n_4324;
wire n_842;
wire n_3626;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_742;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_4396;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_3064;
wire n_2904;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_4114;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_837;
wire n_812;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_509;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4351;
wire n_3340;
wire n_4192;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_3836;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_624;
wire n_3507;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_3864;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_4050;
wire n_3173;
wire n_3732;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_4306;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_602;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_805;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_695;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_730;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_4289;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1524;
wire n_1856;
wire n_1733;
wire n_2016;
wire n_1476;
wire n_2667;
wire n_2725;
wire n_3925;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_651;
wire n_3167;
wire n_1874;
wire n_1293;
wire n_2850;
wire n_3746;
wire n_961;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_726;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_771;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_649;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_586;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_686;
wire n_4279;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_4330;
wire n_1130;
wire n_1450;
wire n_4152;
wire n_3718;
wire n_756;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_3140;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_2986;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2890;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2813;
wire n_515;
wire n_3455;
wire n_807;
wire n_3736;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3605;
wire n_3345;
wire n_2170;
wire n_3560;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4404;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_4377;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2477;
wire n_2314;
wire n_2279;
wire n_3169;
wire n_594;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4301;
wire n_3573;
wire n_2203;
wire n_2076;
wire n_2133;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_3291;
wire n_3654;
wire n_4188;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_4140;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_3982;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_2771;
wire n_3755;
wire n_1090;
wire n_2403;
wire n_3842;
wire n_2947;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_928;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_3769;
wire n_4078;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_562;
wire n_4070;
wire n_2020;
wire n_748;
wire n_3987;
wire n_2310;
wire n_510;
wire n_4249;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_4139;
wire n_914;
wire n_689;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_644;
wire n_3462;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_588;
wire n_3358;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4370;
wire n_3444;
wire n_4368;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_4091;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_667;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_4184;
wire n_846;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_2935;
wire n_4246;
wire n_715;
wire n_889;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1066;
wire n_1549;
wire n_4355;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_685;
wire n_911;
wire n_4061;
wire n_2658;
wire n_623;
wire n_3587;
wire n_3509;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_4155;
wire n_810;
wire n_3376;
wire n_3381;
wire n_4278;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_617;
wire n_3770;
wire n_4375;
wire n_2396;
wire n_3243;
wire n_543;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_3927;
wire n_628;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_743;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_3790;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_4241;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_639;
wire n_673;
wire n_3288;
wire n_3251;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_571;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3904;
wire n_3887;
wire n_593;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_526;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_4366;
wire n_1157;
wire n_1584;
wire n_4384;
wire n_848;
wire n_1664;
wire n_3481;
wire n_629;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_4210;
wire n_532;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_540;
wire n_2624;
wire n_692;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_3926;
wire n_4209;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_4004;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_621;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_697;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_622;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_3751;
wire n_2299;
wire n_4388;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_4110;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_4217;
wire n_530;
wire n_1785;
wire n_1262;
wire n_792;
wire n_4271;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_580;
wire n_3664;
wire n_1579;
wire n_494;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_3873;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_508;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_558;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3576;
wire n_3558;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_4053;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_581;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_4105;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_679;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_663;
wire n_2409;
wire n_3163;
wire n_2966;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_3360;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_765;
wire n_2787;
wire n_4092;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_4057;
wire n_2770;
wire n_631;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_4144;
wire n_4335;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_2012;
wire n_1937;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_633;
wire n_900;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_761;
wire n_2212;
wire n_733;
wire n_3838;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_2897;
wire n_4339;
wire n_1322;
wire n_3273;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_4300;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_1865;
wire n_1710;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2699;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_1792;
wire n_4064;
wire n_504;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_3970;
wire n_4371;
wire n_778;
wire n_1619;
wire n_2351;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_4080;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_3898;
wire n_2541;
wire n_694;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3232;
wire n_3001;
wire n_3188;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_4295;
wire n_3932;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_671;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_4087;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_4238;
wire n_904;
wire n_505;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_498;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_4397;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_539;
wire n_1150;
wire n_4266;
wire n_977;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_4373;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_4407;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_4165;
wire n_4154;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_4380;
wire n_4361;
wire n_3941;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4258;
wire n_2846;
wire n_4298;
wire n_3371;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_4250;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_881;
wire n_1019;
wire n_1777;
wire n_1477;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_4211;
wire n_3094;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_4408;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_4036;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_3918;
wire n_716;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_3244;
wire n_4383;
wire n_3499;
wire n_4391;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_4095;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_656;
wire n_574;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_3361;
wire n_2995;
wire n_3293;
wire n_4287;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3327;
wire n_3228;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3779;
wire n_3895;
wire n_3149;
wire n_1063;
wire n_537;
wire n_3934;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_4338;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_4224;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_583;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_626;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_946;
wire n_3058;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_3986;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_3399;
wire n_1702;
wire n_3894;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_4120;
wire n_4149;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2880;
wire n_2819;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4222;
wire n_1871;
wire n_803;
wire n_2514;
wire n_718;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_548;
wire n_3427;
wire n_2336;
wire n_523;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_4046;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_3041;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_268),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_170),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_381),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_126),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_198),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_241),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_276),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_145),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_92),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_126),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_188),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_51),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_414),
.Y(n_506)
);

BUFx2_ASAP7_75t_SL g507 ( 
.A(n_201),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_134),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_416),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_206),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_338),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_367),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_166),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_234),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_129),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_318),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_76),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_476),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_20),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_368),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_398),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_102),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_234),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_14),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_159),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_29),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_417),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_384),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_54),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_288),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_17),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_94),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_197),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_330),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_151),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_469),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_144),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_278),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_71),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_85),
.Y(n_541)
);

BUFx5_ASAP7_75t_L g542 ( 
.A(n_430),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_463),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_325),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_324),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_57),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_479),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_256),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_22),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_333),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_166),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_314),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_36),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_340),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_83),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_292),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_404),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_204),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_262),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_491),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_150),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_310),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_215),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_48),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_164),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_222),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_431),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_118),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_169),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_314),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_320),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_160),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_349),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_73),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_316),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_327),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_318),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_79),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_278),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_424),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_231),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_219),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_113),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_409),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_4),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_493),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_351),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_350),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_328),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_109),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_184),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_331),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_172),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_326),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_113),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_306),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_62),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_311),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_482),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_104),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_331),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_313),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_455),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_51),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_291),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_196),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_270),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_141),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_108),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_434),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_226),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_484),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_403),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_224),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_193),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_442),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_466),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_447),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_219),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_413),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_248),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_481),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_254),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_39),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_348),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_229),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_112),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_344),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_220),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_353),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_308),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_181),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_334),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_47),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_154),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_423),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_60),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_52),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_138),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_136),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_221),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_432),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_123),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_14),
.Y(n_647)
);

CKINVDCx16_ASAP7_75t_R g648 ( 
.A(n_316),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_429),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_375),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_12),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_483),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_112),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_304),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_12),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_96),
.Y(n_656)
);

CKINVDCx16_ASAP7_75t_R g657 ( 
.A(n_152),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_170),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_313),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_168),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_388),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_212),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_437),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_103),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_232),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_1),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_322),
.Y(n_667)
);

CKINVDCx14_ASAP7_75t_R g668 ( 
.A(n_322),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_488),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_317),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_244),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_365),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_465),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_263),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_224),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_419),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_449),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_144),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_327),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_473),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_1),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_188),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_61),
.Y(n_683)
);

BUFx2_ASAP7_75t_SL g684 ( 
.A(n_20),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_450),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_43),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_61),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_397),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_29),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_110),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_173),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_422),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_244),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_124),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_262),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_141),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_13),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_66),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_492),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_370),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_6),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_206),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_288),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_383),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_342),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_46),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_406),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_196),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_176),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_328),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_150),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_54),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_7),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_269),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_18),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_62),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_204),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_85),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_199),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_81),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_435),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_336),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_232),
.Y(n_723)
);

CKINVDCx16_ASAP7_75t_R g724 ( 
.A(n_390),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_151),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_104),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_348),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_84),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_364),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_174),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_108),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_2),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_474),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_75),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_129),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_148),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_140),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_452),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_70),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_342),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_190),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_380),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_223),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_373),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_22),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_179),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_68),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_237),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_40),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_309),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_378),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_338),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_428),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_410),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_286),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_444),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_19),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_462),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_307),
.Y(n_759)
);

BUFx5_ASAP7_75t_L g760 ( 
.A(n_160),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_356),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_279),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_73),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_49),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_24),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_179),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_111),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_123),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_361),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_402),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_5),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_377),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_77),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_47),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_251),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_19),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_48),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_443),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_52),
.Y(n_779)
);

BUFx5_ASAP7_75t_L g780 ( 
.A(n_227),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_128),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_116),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_5),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_9),
.Y(n_784)
);

CKINVDCx14_ASAP7_75t_R g785 ( 
.A(n_69),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_247),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_9),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_46),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_420),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_326),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_287),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_237),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_400),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_242),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_284),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_88),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_190),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_180),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_454),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_161),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_10),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_323),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_153),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_114),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_241),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_63),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_199),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_438),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_271),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_705),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_536),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_705),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_705),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_705),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_705),
.Y(n_816)
);

INVxp33_ASAP7_75t_SL g817 ( 
.A(n_497),
.Y(n_817)
);

INVxp33_ASAP7_75t_SL g818 ( 
.A(n_612),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_705),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_507),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_705),
.Y(n_821)
);

INVxp33_ASAP7_75t_SL g822 ( 
.A(n_507),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_705),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_705),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_760),
.Y(n_826)
);

INVxp33_ASAP7_75t_SL g827 ( 
.A(n_684),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_760),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_760),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_760),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_760),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_760),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_760),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_760),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_536),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_780),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

INVxp33_ASAP7_75t_SL g838 ( 
.A(n_684),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_780),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_780),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_780),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_780),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_780),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_780),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_661),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_648),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_780),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_536),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_522),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_522),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_543),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_657),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_576),
.Y(n_853)
);

INVxp67_ASAP7_75t_SL g854 ( 
.A(n_530),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_494),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_543),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_508),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_557),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_557),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_577),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_508),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_577),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_772),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_508),
.Y(n_864)
);

CKINVDCx14_ASAP7_75t_R g865 ( 
.A(n_668),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_785),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_588),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_588),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_589),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_589),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_590),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_772),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_590),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_528),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_621),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_508),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_621),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_669),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_720),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_669),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_495),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_676),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_676),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_530),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_680),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_580),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_580),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_642),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_642),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_499),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_502),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_651),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_508),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_808),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_651),
.Y(n_895)
);

CKINVDCx14_ASAP7_75t_R g896 ( 
.A(n_633),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_495),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_499),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_505),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_505),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_791),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_680),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_573),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_699),
.Y(n_904)
);

INVxp33_ASAP7_75t_L g905 ( 
.A(n_510),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_685),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_699),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_721),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_791),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_721),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_744),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_744),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_799),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_791),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_571),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_791),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_704),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_793),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_799),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_571),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_791),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_510),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_513),
.Y(n_923)
);

INVxp67_ASAP7_75t_SL g924 ( 
.A(n_513),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_498),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_808),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_514),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_514),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_515),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_515),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_501),
.Y(n_931)
);

INVxp33_ASAP7_75t_L g932 ( 
.A(n_516),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_516),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_524),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_524),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_532),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_532),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_503),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_724),
.Y(n_939)
);

BUFx5_ASAP7_75t_L g940 ( 
.A(n_633),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_527),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_567),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_567),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_540),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_549),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_533),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_533),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_538),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_554),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_538),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_539),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_539),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_548),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_548),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_552),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_504),
.Y(n_956)
);

INVxp33_ASAP7_75t_L g957 ( 
.A(n_552),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_579),
.B(n_0),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_579),
.Y(n_959)
);

INVxp67_ASAP7_75t_SL g960 ( 
.A(n_565),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_863),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_863),
.B(n_584),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_917),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_814),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_814),
.Y(n_965)
);

AND2x6_ASAP7_75t_L g966 ( 
.A(n_825),
.B(n_585),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_915),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_872),
.B(n_584),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_814),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_872),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_921),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_915),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_817),
.A2(n_724),
.B1(n_570),
.B2(n_575),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_814),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_814),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_845),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_940),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_894),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_920),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_921),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_894),
.B(n_605),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_905),
.B(n_753),
.Y(n_982)
);

BUFx12f_ASAP7_75t_L g983 ( 
.A(n_846),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_845),
.Y(n_984)
);

OA21x2_ASAP7_75t_L g985 ( 
.A1(n_810),
.A2(n_700),
.B(n_585),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_845),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_845),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_810),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_852),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_941),
.Y(n_990)
);

AOI22x1_ASAP7_75t_SL g991 ( 
.A1(n_944),
.A2(n_611),
.B1(n_626),
.B2(n_555),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_845),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_879),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_812),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_825),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_857),
.Y(n_996)
);

CKINVDCx11_ASAP7_75t_R g997 ( 
.A(n_949),
.Y(n_997)
);

OA21x2_ASAP7_75t_L g998 ( 
.A1(n_812),
.A2(n_761),
.B(n_700),
.Y(n_998)
);

OAI22x1_ASAP7_75t_L g999 ( 
.A1(n_881),
.A2(n_500),
.B1(n_641),
.B2(n_556),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_925),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_811),
.B(n_605),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_834),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_835),
.B(n_662),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_834),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_932),
.B(n_544),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_857),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_837),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_849),
.B(n_662),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_837),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_813),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_813),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_L g1012 ( 
.A(n_940),
.B(n_956),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_849),
.B(n_702),
.Y(n_1013)
);

CKINVDCx11_ASAP7_75t_R g1014 ( 
.A(n_874),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_842),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_818),
.A2(n_698),
.B1(n_762),
.B2(n_718),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_926),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_842),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_861),
.Y(n_1019)
);

OAI22x1_ASAP7_75t_SL g1020 ( 
.A1(n_903),
.A2(n_764),
.B1(n_750),
.B2(n_670),
.Y(n_1020)
);

XNOR2x2_ASAP7_75t_L g1021 ( 
.A(n_855),
.B(n_565),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_815),
.A2(n_761),
.B(n_756),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_957),
.B(n_544),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_884),
.B(n_544),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_896),
.B(n_560),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_942),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_939),
.A2(n_702),
.B1(n_511),
.B2(n_519),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_940),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_897),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_861),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_931),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_866),
.B(n_633),
.Y(n_1032)
);

AOI22x1_ASAP7_75t_SL g1033 ( 
.A1(n_906),
.A2(n_523),
.B1(n_525),
.B2(n_517),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_815),
.Y(n_1034)
);

INVxp33_ASAP7_75t_SL g1035 ( 
.A(n_918),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_816),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_891),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_884),
.B(n_604),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_864),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_942),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_864),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_876),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_876),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_822),
.A2(n_569),
.B1(n_583),
.B2(n_566),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_945),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_893),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_893),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_816),
.A2(n_509),
.B(n_550),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_850),
.B(n_550),
.Y(n_1049)
);

INVx5_ASAP7_75t_L g1050 ( 
.A(n_943),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_914),
.Y(n_1051)
);

INVx6_ASAP7_75t_L g1052 ( 
.A(n_940),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_926),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_819),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_854),
.B(n_544),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_914),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_916),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_819),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_916),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_887),
.B(n_603),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_821),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_940),
.B(n_560),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_821),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_823),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_943),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_853),
.A2(n_827),
.B1(n_838),
.B2(n_958),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_938),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_823),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_940),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_824),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_892),
.B(n_679),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_850),
.B(n_661),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_895),
.B(n_679),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_824),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_826),
.A2(n_614),
.B(n_572),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_826),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_959),
.A2(n_804),
.B1(n_806),
.B2(n_802),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_890),
.A2(n_569),
.B1(n_583),
.B2(n_566),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_940),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_940),
.B(n_496),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_828),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_828),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_940),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_959),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_829),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_829),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1002),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1002),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_967),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1002),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_990),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1017),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1000),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1000),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1045),
.B(n_820),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1017),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1054),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1000),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_963),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1004),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1014),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_997),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_982),
.B(n_851),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_983),
.B(n_865),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1017),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1035),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1053),
.Y(n_1107)
);

CKINVDCx16_ASAP7_75t_R g1108 ( 
.A(n_983),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1037),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_983),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1053),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_961),
.B(n_901),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_989),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1004),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1053),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1004),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1072),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_982),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1072),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_1016),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_989),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1085),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_989),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1054),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1054),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1081),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1081),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_971),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_970),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1005),
.B(n_851),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_993),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1007),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1085),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_971),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_967),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_980),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_980),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_993),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_961),
.B(n_909),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_993),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_978),
.B(n_856),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_L g1142 ( 
.A(n_1025),
.B(n_862),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1007),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_979),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1005),
.B(n_924),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_979),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1023),
.B(n_950),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1016),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1023),
.B(n_954),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_995),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_995),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1085),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_972),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1084),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1084),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1084),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_995),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_995),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1081),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1077),
.A2(n_775),
.B1(n_779),
.B2(n_675),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1009),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1009),
.Y(n_1162)
);

BUFx8_ASAP7_75t_L g1163 ( 
.A(n_972),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_R g1164 ( 
.A(n_1012),
.B(n_856),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1007),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1015),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1015),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1015),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1009),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_978),
.B(n_858),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_973),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1063),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1001),
.B(n_858),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1085),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1085),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1009),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1063),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1031),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1063),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_991),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1064),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1064),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1049),
.B(n_960),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1064),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1068),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1049),
.B(n_922),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1001),
.B(n_859),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1068),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_991),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_970),
.B(n_859),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1068),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_L g1192 ( 
.A(n_1048),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1031),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1070),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1001),
.B(n_860),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_970),
.B(n_947),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1001),
.B(n_860),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1033),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1033),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1070),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1085),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_SL g1203 ( 
.A(n_1003),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1082),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1082),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1020),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1075),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1003),
.B(n_862),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1020),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1032),
.B(n_877),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1067),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1086),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1029),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1086),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_L g1216 ( 
.A(n_1028),
.B(n_542),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1086),
.Y(n_1217)
);

CKINVDCx16_ASAP7_75t_R g1218 ( 
.A(n_1066),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1075),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_988),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_988),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1066),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1081),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_994),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1062),
.A2(n_831),
.B(n_830),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1049),
.B(n_922),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_994),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1021),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1049),
.B(n_923),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1010),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_996),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_1003),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1077),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1003),
.B(n_948),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1021),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1027),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1010),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1011),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1011),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1034),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_996),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1024),
.B(n_923),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1034),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1024),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1036),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1036),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1044),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1058),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1038),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_996),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1008),
.B(n_951),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1058),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1038),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1044),
.B(n_868),
.C(n_867),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1061),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1061),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_996),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1055),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1055),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1060),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1074),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1060),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1074),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1071),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1071),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1076),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1076),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1073),
.B(n_867),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1073),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_962),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_R g1271 ( 
.A(n_1050),
.B(n_868),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_962),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1019),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_999),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1078),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_962),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_962),
.B(n_869),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_999),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1019),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_968),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_968),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_968),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_996),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_968),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_981),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1078),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1008),
.B(n_953),
.Y(n_1287)
);

BUFx8_ASAP7_75t_L g1288 ( 
.A(n_981),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_981),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_996),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_981),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_966),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1019),
.Y(n_1293)
);

AND2x2_ASAP7_75t_SL g1294 ( 
.A(n_1048),
.B(n_572),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_966),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1039),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1008),
.B(n_955),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1008),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_966),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1039),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1039),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_966),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1047),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1047),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1006),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1047),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1059),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1059),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1013),
.B(n_927),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1013),
.B(n_955),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1059),
.Y(n_1311)
);

XOR2xp5_ASAP7_75t_L g1312 ( 
.A(n_1013),
.B(n_886),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1013),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1048),
.Y(n_1314)
);

BUFx10_ASAP7_75t_L g1315 ( 
.A(n_1099),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1234),
.B(n_1028),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1178),
.B(n_888),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1232),
.B(n_977),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1220),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1259),
.A2(n_869),
.B1(n_871),
.B2(n_870),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1087),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1095),
.B(n_889),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1221),
.Y(n_1323)
);

INVxp33_ASAP7_75t_L g1324 ( 
.A(n_1193),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1224),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1227),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1269),
.B(n_977),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1234),
.B(n_1069),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1230),
.Y(n_1329)
);

BUFx8_ASAP7_75t_SL g1330 ( 
.A(n_1101),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1087),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1238),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1118),
.B(n_977),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1088),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1239),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1234),
.B(n_1069),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1240),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1243),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1088),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1258),
.B(n_977),
.Y(n_1340)
);

AND2x6_ASAP7_75t_L g1341 ( 
.A(n_1314),
.B(n_870),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1265),
.B(n_1083),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1203),
.A2(n_1048),
.B1(n_1022),
.B2(n_966),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1090),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_SL g1345 ( 
.A(n_1093),
.B(n_633),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1245),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1246),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1207),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1268),
.B(n_1083),
.Y(n_1349)
);

BUFx4f_ASAP7_75t_L g1350 ( 
.A(n_1145),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1248),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1252),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1090),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1251),
.B(n_871),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1255),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1190),
.B(n_1083),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1256),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1129),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1203),
.A2(n_1022),
.B1(n_966),
.B2(n_782),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1251),
.B(n_1310),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1097),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1266),
.Y(n_1362)
);

AND3x1_ASAP7_75t_L g1363 ( 
.A(n_1089),
.B(n_596),
.C(n_593),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1292),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1135),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1267),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1097),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1128),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1134),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1292),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1251),
.B(n_927),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1288),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1136),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1207),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1232),
.B(n_1083),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1100),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1137),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1259),
.B(n_531),
.C(n_526),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1173),
.B(n_1022),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1097),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1126),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1203),
.A2(n_1022),
.B1(n_966),
.B2(n_875),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1100),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1126),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1153),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1114),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1126),
.Y(n_1387)
);

INVx5_ASAP7_75t_L g1388 ( 
.A(n_1207),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1294),
.A2(n_985),
.B1(n_998),
.B2(n_966),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1232),
.B(n_1079),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1127),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1287),
.B(n_928),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1114),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1127),
.B(n_1079),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1294),
.A2(n_998),
.B1(n_985),
.B2(n_875),
.Y(n_1395)
);

INVx4_ASAP7_75t_SL g1396 ( 
.A(n_1207),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1127),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1212),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1159),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1116),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1228),
.A2(n_535),
.B1(n_541),
.B2(n_534),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1159),
.B(n_1079),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1159),
.B(n_1079),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1212),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1237),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1295),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1187),
.B(n_1080),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1116),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1198),
.B(n_1052),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1237),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1261),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1132),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1261),
.Y(n_1413)
);

AO22x2_ASAP7_75t_L g1414 ( 
.A1(n_1228),
.A2(n_877),
.B1(n_878),
.B2(n_873),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1132),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1170),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1219),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_L g1418 ( 
.A(n_1219),
.B(n_1079),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1287),
.B(n_1297),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1263),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1264),
.B(n_1052),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1145),
.B(n_1052),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1219),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1143),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1164),
.B(n_1079),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1260),
.B(n_546),
.C(n_545),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1219),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1143),
.Y(n_1428)
);

INVx4_ASAP7_75t_SL g1429 ( 
.A(n_1219),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1091),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1099),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1263),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1165),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1208),
.B(n_1052),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1165),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1166),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1313),
.B(n_1052),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1260),
.B(n_553),
.C(n_551),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1147),
.B(n_928),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1214),
.B(n_929),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1262),
.A2(n_558),
.B1(n_561),
.B2(n_559),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_SL g1442 ( 
.A(n_1106),
.B(n_873),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1286),
.A2(n_998),
.B1(n_985),
.B2(n_880),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1091),
.Y(n_1444)
);

CKINVDCx6p67_ASAP7_75t_R g1445 ( 
.A(n_1108),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1287),
.B(n_929),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1192),
.B(n_1079),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1297),
.B(n_930),
.Y(n_1448)
);

BUFx10_ASAP7_75t_L g1449 ( 
.A(n_1106),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1192),
.B(n_1018),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1150),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1147),
.B(n_1149),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1295),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1149),
.B(n_1050),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1270),
.B(n_1050),
.Y(n_1455)
);

BUFx10_ASAP7_75t_L g1456 ( 
.A(n_1093),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1151),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1122),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1242),
.B(n_1050),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1157),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1166),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1242),
.B(n_1050),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1130),
.B(n_1050),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1223),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1262),
.B(n_1286),
.C(n_1171),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1167),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1192),
.B(n_1018),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1158),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1129),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1297),
.B(n_1310),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1299),
.Y(n_1471)
);

BUFx10_ASAP7_75t_L g1472 ( 
.A(n_1094),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1144),
.B(n_930),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1167),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1168),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1168),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1172),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1288),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1196),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1122),
.Y(n_1480)
);

INVxp33_ASAP7_75t_L g1481 ( 
.A(n_1312),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1223),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1172),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1122),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1161),
.Y(n_1485)
);

CKINVDCx6p67_ASAP7_75t_R g1486 ( 
.A(n_1109),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1310),
.B(n_1050),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1162),
.Y(n_1488)
);

NAND2x1p5_ASAP7_75t_L g1489 ( 
.A(n_1186),
.B(n_1065),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1122),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1288),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1247),
.A2(n_998),
.B1(n_985),
.B2(n_880),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1247),
.A2(n_882),
.B1(n_883),
.B2(n_878),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1181),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1133),
.B(n_1018),
.Y(n_1495)
);

BUFx10_ASAP7_75t_L g1496 ( 
.A(n_1094),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1133),
.B(n_1018),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1169),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1144),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1275),
.A2(n_883),
.B1(n_885),
.B2(n_882),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1181),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1186),
.B(n_933),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1275),
.A2(n_902),
.B1(n_904),
.B2(n_885),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1146),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1176),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1142),
.A2(n_904),
.B1(n_907),
.B2(n_902),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1092),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1103),
.B(n_1065),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1146),
.B(n_933),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1133),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1191),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1109),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1191),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1195),
.A2(n_908),
.B1(n_910),
.B2(n_907),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1096),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1309),
.B(n_934),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1194),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1177),
.A2(n_910),
.B(n_908),
.Y(n_1518)
);

INVx8_ASAP7_75t_L g1519 ( 
.A(n_1299),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1105),
.Y(n_1520)
);

INVx4_ASAP7_75t_L g1521 ( 
.A(n_1302),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1194),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1215),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1281),
.B(n_1065),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1272),
.B(n_1065),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1110),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1110),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1107),
.Y(n_1528)
);

CKINVDCx8_ASAP7_75t_R g1529 ( 
.A(n_1101),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1179),
.A2(n_912),
.B(n_911),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1133),
.B(n_1018),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1215),
.Y(n_1532)
);

BUFx10_ASAP7_75t_L g1533 ( 
.A(n_1098),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1273),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1141),
.B(n_1065),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1111),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1273),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1115),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1279),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1309),
.B(n_1065),
.Y(n_1540)
);

AND2x6_ASAP7_75t_L g1541 ( 
.A(n_1211),
.B(n_911),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1280),
.B(n_1065),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1226),
.B(n_934),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1124),
.Y(n_1544)
);

NOR2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1098),
.B(n_898),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1298),
.B(n_912),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1125),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1279),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1231),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1152),
.B(n_1018),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1182),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1235),
.A2(n_919),
.B1(n_913),
.B2(n_673),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1113),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1163),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1276),
.B(n_1282),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1152),
.B(n_1018),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1184),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1196),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1244),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1196),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1113),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1473),
.B(n_1171),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1519),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1371),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1350),
.B(n_1152),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1419),
.B(n_1226),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1321),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1452),
.B(n_1244),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1358),
.B(n_1469),
.Y(n_1569)
);

INVx4_ASAP7_75t_L g1570 ( 
.A(n_1360),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1419),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1439),
.B(n_1183),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1350),
.B(n_1222),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1348),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1360),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1371),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1419),
.B(n_1446),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1470),
.A2(n_1253),
.B1(n_1249),
.B2(n_1236),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1509),
.B(n_1398),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1419),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1446),
.B(n_1229),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1404),
.B(n_1249),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1446),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1446),
.B(n_1229),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1478),
.B(n_1491),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1465),
.B(n_1222),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1430),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1479),
.Y(n_1588)
);

NAND2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1358),
.B(n_1231),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1371),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1502),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1392),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1478),
.B(n_1183),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1392),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1431),
.A2(n_1233),
.B1(n_1236),
.B2(n_1120),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1392),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1491),
.B(n_1284),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1448),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1448),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1448),
.B(n_1285),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1502),
.A2(n_1235),
.B1(n_1254),
.B2(n_1289),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1321),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1319),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1331),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1479),
.B(n_1218),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1558),
.B(n_1253),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1323),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1464),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1422),
.B(n_1291),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1348),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1325),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1331),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1348),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1422),
.B(n_1421),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1558),
.B(n_1233),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1326),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1431),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1329),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1330),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1332),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1502),
.B(n_1543),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1388),
.B(n_1152),
.Y(n_1622)
);

CKINVDCx11_ASAP7_75t_R g1623 ( 
.A(n_1529),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1335),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1502),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1360),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1334),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1348),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1543),
.B(n_1277),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1444),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1374),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1334),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1322),
.B(n_1154),
.Y(n_1633)
);

NAND3x1_ASAP7_75t_L g1634 ( 
.A(n_1330),
.B(n_1102),
.C(n_1163),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1543),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1374),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1559),
.B(n_1154),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1543),
.B(n_1121),
.Y(n_1638)
);

AND2x2_ASAP7_75t_SL g1639 ( 
.A(n_1418),
.B(n_1216),
.Y(n_1639)
);

INVx4_ASAP7_75t_L g1640 ( 
.A(n_1360),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1445),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1464),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1337),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1338),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1464),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1499),
.B(n_1155),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1360),
.A2(n_1160),
.B1(n_1121),
.B2(n_1131),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1421),
.B(n_1112),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1516),
.B(n_1139),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1320),
.B(n_1117),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1516),
.B(n_1123),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1442),
.A2(n_1138),
.B1(n_1140),
.B2(n_1131),
.C(n_1123),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1346),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1347),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1354),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1351),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1352),
.Y(n_1657)
);

NOR2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1486),
.B(n_1102),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1504),
.B(n_1155),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1355),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1357),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1339),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1385),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1442),
.A2(n_1140),
.B1(n_1138),
.B2(n_1156),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1362),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1374),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1482),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1516),
.B(n_1156),
.Y(n_1668)
);

INVx8_ASAP7_75t_L g1669 ( 
.A(n_1354),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1366),
.Y(n_1670)
);

INVx5_ASAP7_75t_L g1671 ( 
.A(n_1519),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1440),
.B(n_1104),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1512),
.B(n_1274),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1354),
.A2(n_1120),
.B1(n_1148),
.B2(n_1216),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1482),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1368),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1369),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1482),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1493),
.B(n_1185),
.Y(n_1679)
);

INVx5_ASAP7_75t_L g1680 ( 
.A(n_1519),
.Y(n_1680)
);

AND2x6_ASAP7_75t_L g1681 ( 
.A(n_1343),
.B(n_1119),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1500),
.A2(n_1278),
.B1(n_1274),
.B2(n_564),
.C(n_568),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1372),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1373),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1374),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1377),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1339),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1344),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1414),
.B(n_1148),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1354),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1405),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1316),
.A2(n_1197),
.B1(n_1201),
.B2(n_1188),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1344),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1410),
.Y(n_1694)
);

CKINVDCx20_ASAP7_75t_R g1695 ( 
.A(n_1486),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1411),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1353),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1413),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1469),
.B(n_1231),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1353),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1381),
.B(n_1204),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1340),
.B(n_1205),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1340),
.B(n_1342),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1372),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1376),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1545),
.B(n_1302),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1372),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1503),
.A2(n_1278),
.B1(n_574),
.B2(n_578),
.C(n_563),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1364),
.B(n_1250),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1388),
.B(n_1423),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1345),
.A2(n_1210),
.B1(n_1206),
.B2(n_1200),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1526),
.B(n_935),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1420),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1519),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1388),
.B(n_1174),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1376),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1526),
.B(n_935),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1432),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1365),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1383),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1423),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1342),
.B(n_1209),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1364),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1354),
.A2(n_1163),
.B1(n_1217),
.B2(n_1213),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1544),
.Y(n_1725)
);

OAI21xp33_ASAP7_75t_L g1726 ( 
.A1(n_1441),
.A2(n_646),
.B(n_636),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1317),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1416),
.B(n_1293),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1383),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1315),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1423),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1381),
.B(n_1225),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1328),
.A2(n_1175),
.B1(n_1202),
.B2(n_1174),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1416),
.B(n_1296),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1364),
.B(n_1250),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1414),
.A2(n_919),
.B1(n_913),
.B2(n_1301),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1445),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1546),
.B(n_1304),
.Y(n_1738)
);

OR2x2_ASAP7_75t_SL g1739 ( 
.A(n_1378),
.B(n_1199),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1388),
.B(n_1174),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1333),
.B(n_1306),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1315),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1547),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1386),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1370),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1423),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1324),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1386),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1333),
.B(n_1307),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1381),
.B(n_1391),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1327),
.B(n_659),
.C(n_637),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1327),
.B(n_1308),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1414),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1527),
.B(n_936),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1507),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1515),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1324),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1520),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1391),
.B(n_1225),
.Y(n_1759)
);

AND2x6_ASAP7_75t_L g1760 ( 
.A(n_1427),
.B(n_1174),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1393),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1336),
.A2(n_1202),
.B1(n_1175),
.B2(n_1225),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1315),
.B(n_1206),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1527),
.B(n_1210),
.Y(n_1764)
);

NAND3x1_ASAP7_75t_L g1765 ( 
.A(n_1529),
.B(n_1200),
.C(n_1199),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1391),
.B(n_1250),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1528),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1536),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1489),
.Y(n_1769)
);

AND2x6_ASAP7_75t_L g1770 ( 
.A(n_1427),
.B(n_1175),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1538),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1551),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1481),
.B(n_936),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1557),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1553),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1449),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1553),
.B(n_937),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1449),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1427),
.B(n_1175),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1451),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1393),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1481),
.B(n_937),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1457),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1506),
.B(n_1454),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1561),
.B(n_946),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1427),
.Y(n_1786)
);

CKINVDCx14_ASAP7_75t_R g1787 ( 
.A(n_1449),
.Y(n_1787)
);

BUFx10_ASAP7_75t_L g1788 ( 
.A(n_1541),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1458),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1400),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1458),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1396),
.Y(n_1792)
);

CKINVDCx14_ASAP7_75t_R g1793 ( 
.A(n_1456),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1426),
.B(n_1290),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1460),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1561),
.B(n_1554),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1396),
.B(n_1202),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1370),
.B(n_946),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1400),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1468),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1456),
.Y(n_1801)
);

BUFx4f_ASAP7_75t_L g1802 ( 
.A(n_1541),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1438),
.B(n_1290),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1370),
.B(n_948),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1552),
.B(n_951),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1485),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1488),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1408),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1498),
.Y(n_1809)
);

NAND2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1406),
.B(n_1290),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1572),
.B(n_1514),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1562),
.A2(n_1363),
.B1(n_1541),
.B2(n_1472),
.Y(n_1812)
);

AO22x1_ASAP7_75t_L g1813 ( 
.A1(n_1573),
.A2(n_1189),
.B1(n_1180),
.B2(n_1541),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1641),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1568),
.B(n_1456),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1578),
.B(n_1472),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1736),
.A2(n_1401),
.B1(n_1454),
.B2(n_1341),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_SL g1818 ( 
.A(n_1617),
.B(n_582),
.C(n_562),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1606),
.B(n_1472),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1603),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1639),
.B(n_1614),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1650),
.B(n_1541),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1719),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1579),
.B(n_1496),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1607),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1737),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1567),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1606),
.B(n_1496),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1639),
.B(n_1396),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1683),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1802),
.B(n_1429),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1650),
.B(n_1555),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1573),
.B(n_1341),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1600),
.B(n_1341),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1623),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1792),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1611),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1581),
.B(n_1341),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1584),
.B(n_1341),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1584),
.B(n_1455),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1792),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1777),
.B(n_1455),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1785),
.B(n_1407),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1633),
.A2(n_1533),
.B1(n_1496),
.B2(n_1524),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1727),
.B(n_1505),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1582),
.A2(n_1533),
.B1(n_1524),
.B2(n_1406),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1802),
.B(n_1429),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1567),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1616),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1727),
.B(n_1180),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_SL g1852 ( 
.A1(n_1689),
.A2(n_1189),
.B1(n_1533),
.B2(n_1453),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1564),
.B(n_1361),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1602),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1618),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1576),
.B(n_1361),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1747),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1663),
.B(n_1586),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1590),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1672),
.A2(n_1406),
.B1(n_1471),
.B2(n_1453),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1602),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1592),
.B(n_1594),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1669),
.B(n_1453),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1683),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1577),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1585),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1595),
.A2(n_1521),
.B1(n_1471),
.B2(n_604),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1570),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1736),
.A2(n_1518),
.B1(n_1530),
.B2(n_1477),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1663),
.B(n_1384),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1586),
.A2(n_586),
.B1(n_594),
.B2(n_592),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1620),
.Y(n_1872)
);

OR2x6_ASAP7_75t_L g1873 ( 
.A(n_1669),
.B(n_1471),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1703),
.B(n_1429),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1621),
.A2(n_1521),
.B1(n_1437),
.B2(n_1525),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1721),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1596),
.B(n_1361),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1598),
.B(n_1367),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1599),
.B(n_1367),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1624),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1577),
.B(n_1521),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1588),
.B(n_1367),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1707),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1604),
.Y(n_1884)
);

INVx8_ASAP7_75t_L g1885 ( 
.A(n_1669),
.Y(n_1885)
);

NAND2x1p5_ASAP7_75t_L g1886 ( 
.A(n_1570),
.B(n_1458),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1588),
.B(n_1380),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1604),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1784),
.B(n_1458),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1615),
.B(n_952),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1615),
.B(n_952),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1671),
.B(n_1680),
.Y(n_1892)
);

BUFx8_ASAP7_75t_SL g1893 ( 
.A(n_1619),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1575),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1747),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1707),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1630),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1621),
.A2(n_1609),
.B1(n_1722),
.B2(n_1702),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1601),
.B(n_1380),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1612),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1601),
.B(n_1380),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1585),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1704),
.B(n_1480),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1741),
.A2(n_1356),
.B1(n_1417),
.B2(n_1349),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1643),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1612),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1668),
.B(n_1605),
.Y(n_1907)
);

A2O1A1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1732),
.A2(n_1387),
.B(n_1399),
.C(n_1397),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1644),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1653),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1593),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1749),
.A2(n_1417),
.B1(n_1434),
.B2(n_1409),
.Y(n_1912)
);

AND3x1_ASAP7_75t_L g1913 ( 
.A(n_1664),
.B(n_596),
.C(n_593),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1753),
.A2(n_1805),
.B1(n_1674),
.B2(n_1682),
.Y(n_1914)
);

INVx8_ASAP7_75t_L g1915 ( 
.A(n_1566),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1566),
.B(n_1712),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1671),
.B(n_1480),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1654),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1773),
.B(n_1530),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1593),
.B(n_1549),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1627),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1753),
.A2(n_1518),
.B1(n_1477),
.B2(n_1494),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1712),
.B(n_1717),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1717),
.B(n_1754),
.Y(n_1924)
);

OAI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1583),
.A2(n_665),
.B1(n_714),
.B2(n_614),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1656),
.Y(n_1926)
);

AND2x6_ASAP7_75t_SL g1927 ( 
.A(n_1763),
.B(n_598),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1668),
.A2(n_1525),
.B1(n_1542),
.B2(n_1508),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1671),
.B(n_1480),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1627),
.Y(n_1930)
);

O2A1O1Ixp5_ASAP7_75t_L g1931 ( 
.A1(n_1779),
.A2(n_1467),
.B(n_1450),
.C(n_1417),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1754),
.B(n_1379),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1657),
.Y(n_1933)
);

INVx5_ASAP7_75t_L g1934 ( 
.A(n_1575),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1649),
.B(n_1492),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1623),
.Y(n_1936)
);

INVxp67_ASAP7_75t_SL g1937 ( 
.A(n_1583),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1671),
.B(n_1480),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1651),
.A2(n_1542),
.B1(n_1508),
.B2(n_1463),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1752),
.A2(n_1418),
.B(n_1375),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1660),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1730),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1591),
.B(n_1443),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1591),
.B(n_1483),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1661),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1730),
.Y(n_1946)
);

NOR2x1p5_ASAP7_75t_L g1947 ( 
.A(n_1742),
.B(n_1549),
.Y(n_1947)
);

AND2x2_ASAP7_75t_SL g1948 ( 
.A(n_1626),
.B(n_1382),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1625),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_SL g1950 ( 
.A1(n_1695),
.A2(n_595),
.B1(n_599),
.B2(n_597),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1679),
.A2(n_1494),
.B1(n_1501),
.B2(n_1483),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1704),
.B(n_1484),
.Y(n_1952)
);

NOR3xp33_ASAP7_75t_L g1953 ( 
.A(n_1652),
.B(n_600),
.C(n_598),
.Y(n_1953)
);

NOR2x1p5_ASAP7_75t_L g1954 ( 
.A(n_1742),
.B(n_1549),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1625),
.B(n_1635),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1680),
.B(n_1484),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1680),
.B(n_1484),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1605),
.B(n_1459),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1619),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1635),
.B(n_1501),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1665),
.B(n_1511),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1721),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1680),
.B(n_1484),
.Y(n_1963)
);

INVxp67_ASAP7_75t_L g1964 ( 
.A(n_1782),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1670),
.A2(n_1513),
.B1(n_1517),
.B2(n_1511),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1676),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1677),
.B(n_1513),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1684),
.B(n_1517),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1686),
.B(n_1522),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1775),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1632),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1725),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1629),
.B(n_1798),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1629),
.B(n_1522),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1798),
.B(n_1523),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1789),
.B(n_1490),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1632),
.Y(n_1977)
);

CKINVDCx16_ASAP7_75t_R g1978 ( 
.A(n_1695),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1804),
.B(n_1523),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1789),
.B(n_1490),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1732),
.A2(n_1462),
.B(n_1375),
.Y(n_1981)
);

INVx4_ASAP7_75t_L g1982 ( 
.A(n_1626),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1743),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1755),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_SL g1985 ( 
.A1(n_1647),
.A2(n_608),
.B1(n_609),
.B2(n_601),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1804),
.B(n_1532),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1662),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1569),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1789),
.B(n_1490),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1651),
.A2(n_1463),
.B1(n_1390),
.B2(n_1318),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1756),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1571),
.B(n_1580),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1757),
.B(n_1540),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1638),
.B(n_953),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1789),
.B(n_1490),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1758),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1662),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1791),
.B(n_1510),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1791),
.B(n_1510),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1638),
.A2(n_1390),
.B1(n_1318),
.B2(n_1359),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1687),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1580),
.B(n_1395),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1640),
.B(n_1450),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1687),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1708),
.A2(n_1681),
.B1(n_1774),
.B2(n_1772),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1791),
.B(n_1510),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1791),
.B(n_1510),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1681),
.A2(n_1412),
.B1(n_1415),
.B2(n_1408),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1574),
.B(n_1467),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1646),
.A2(n_1487),
.B1(n_1489),
.B2(n_1447),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1688),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1767),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1574),
.B(n_1202),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1597),
.B(n_1412),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1787),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1688),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1693),
.Y(n_2018)
);

NAND2x1p5_ASAP7_75t_L g2019 ( 
.A(n_1640),
.B(n_1495),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1764),
.B(n_899),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1597),
.B(n_1415),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1658),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_SL g2023 ( 
.A1(n_1711),
.A2(n_603),
.B1(n_679),
.B2(n_604),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1780),
.B(n_1783),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1796),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1795),
.B(n_1424),
.Y(n_2026)
);

A2O1A1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1832),
.A2(n_1701),
.B(n_1648),
.C(n_1759),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1949),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1844),
.B(n_1659),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1827),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1820),
.Y(n_2031)
);

OR2x6_ASAP7_75t_L g2032 ( 
.A(n_1885),
.B(n_1915),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1914),
.A2(n_1673),
.B1(n_1681),
.B2(n_1768),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1825),
.Y(n_2034)
);

OR2x6_ASAP7_75t_L g2035 ( 
.A(n_1885),
.B(n_1655),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1865),
.B(n_1706),
.Y(n_2036)
);

OR2x6_ASAP7_75t_L g2037 ( 
.A(n_1885),
.B(n_1915),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1837),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1865),
.B(n_1706),
.Y(n_2039)
);

BUFx8_ASAP7_75t_L g2040 ( 
.A(n_1897),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1850),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_R g2042 ( 
.A(n_1835),
.B(n_1787),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_1830),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1858),
.B(n_1587),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1855),
.Y(n_2045)
);

NAND2xp33_ASAP7_75t_SL g2046 ( 
.A(n_1947),
.B(n_1721),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1830),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1849),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1898),
.B(n_1724),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1872),
.Y(n_2050)
);

CKINVDCx20_ASAP7_75t_R g2051 ( 
.A(n_1893),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1949),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1970),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1994),
.B(n_1793),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1858),
.A2(n_1796),
.B1(n_1637),
.B2(n_1793),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1880),
.Y(n_2056)
);

INVx4_ASAP7_75t_L g2057 ( 
.A(n_1915),
.Y(n_2057)
);

AND3x1_ASAP7_75t_SL g2058 ( 
.A(n_1954),
.B(n_607),
.C(n_600),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1881),
.B(n_1769),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1890),
.B(n_1771),
.Y(n_2060)
);

AOI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_1816),
.A2(n_1726),
.B1(n_1765),
.B2(n_1655),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_SL g2062 ( 
.A(n_1959),
.B(n_1751),
.C(n_629),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1881),
.B(n_1769),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_1836),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_SL g2065 ( 
.A(n_1936),
.B(n_630),
.C(n_622),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1836),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1843),
.B(n_1728),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1905),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1864),
.B(n_1776),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1864),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2020),
.B(n_603),
.Y(n_2071)
);

INVx5_ASAP7_75t_L g2072 ( 
.A(n_1863),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1909),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_2016),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1883),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1910),
.Y(n_2076)
);

NAND2x1p5_ASAP7_75t_L g2077 ( 
.A(n_1934),
.B(n_1797),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1836),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1854),
.Y(n_2079)
);

BUFx2_ASAP7_75t_L g2080 ( 
.A(n_1970),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1884),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1918),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1926),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1933),
.Y(n_2084)
);

NOR3xp33_ASAP7_75t_SL g2085 ( 
.A(n_1978),
.B(n_632),
.C(n_631),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_R g2086 ( 
.A(n_1934),
.B(n_1778),
.Y(n_2086)
);

INVx4_ASAP7_75t_L g2087 ( 
.A(n_1836),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_1955),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1842),
.Y(n_2089)
);

BUFx2_ASAP7_75t_SL g2090 ( 
.A(n_1883),
.Y(n_2090)
);

BUFx3_ASAP7_75t_L g2091 ( 
.A(n_1896),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1941),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1842),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1841),
.B(n_1734),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1822),
.B(n_1721),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1958),
.B(n_1731),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1958),
.B(n_1731),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1888),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_R g2099 ( 
.A(n_1934),
.B(n_1801),
.Y(n_2099)
);

CKINVDCx6p67_ASAP7_75t_R g2100 ( 
.A(n_1896),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1875),
.B(n_1731),
.Y(n_2101)
);

INVx5_ASAP7_75t_L g2102 ( 
.A(n_1863),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_R g2103 ( 
.A(n_1934),
.B(n_1563),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1923),
.B(n_1690),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1891),
.B(n_1800),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_1924),
.B(n_1690),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1900),
.Y(n_2107)
);

NAND3xp33_ASAP7_75t_SL g2108 ( 
.A(n_1816),
.B(n_635),
.C(n_634),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_1842),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1964),
.B(n_1806),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1866),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1842),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1911),
.Y(n_2113)
);

NOR3xp33_ASAP7_75t_SL g2114 ( 
.A(n_1818),
.B(n_640),
.C(n_638),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1819),
.B(n_1807),
.Y(n_2115)
);

OR2x2_ASAP7_75t_SL g2116 ( 
.A(n_1851),
.B(n_1634),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1945),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1876),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1906),
.Y(n_2119)
);

NAND3xp33_ASAP7_75t_L g2120 ( 
.A(n_2006),
.B(n_1794),
.C(n_1803),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1876),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1921),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1966),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_1823),
.Y(n_2124)
);

INVx1_ASAP7_75t_SL g2125 ( 
.A(n_1824),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1907),
.B(n_603),
.Y(n_2126)
);

NAND2xp33_ASAP7_75t_SL g2127 ( 
.A(n_1821),
.B(n_1731),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1819),
.B(n_1809),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1972),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1815),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1983),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1876),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1984),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1916),
.B(n_1857),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1828),
.B(n_1691),
.Y(n_2135)
);

BUFx12f_ASAP7_75t_L g2136 ( 
.A(n_1814),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1991),
.Y(n_2137)
);

BUFx3_ASAP7_75t_L g2138 ( 
.A(n_1902),
.Y(n_2138)
);

INVx4_ASAP7_75t_L g2139 ( 
.A(n_1903),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1930),
.Y(n_2140)
);

BUFx4f_ASAP7_75t_SL g2141 ( 
.A(n_1826),
.Y(n_2141)
);

INVx5_ASAP7_75t_L g2142 ( 
.A(n_1863),
.Y(n_2142)
);

OAI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_1828),
.A2(n_1750),
.B1(n_1701),
.B2(n_1738),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1996),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2013),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1971),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_1838),
.B(n_1565),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_2025),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1977),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2024),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1987),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1993),
.B(n_1694),
.Y(n_2152)
);

BUFx12f_ASAP7_75t_L g2153 ( 
.A(n_1927),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1982),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1993),
.B(n_1696),
.Y(n_2155)
);

INVx4_ASAP7_75t_L g2156 ( 
.A(n_1903),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_R g2157 ( 
.A(n_1868),
.B(n_1563),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1939),
.B(n_1746),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1997),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1988),
.B(n_1565),
.Y(n_2160)
);

NOR3xp33_ASAP7_75t_SL g2161 ( 
.A(n_1950),
.B(n_644),
.C(n_643),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1846),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_1973),
.B(n_1739),
.Y(n_2163)
);

AOI211xp5_ASAP7_75t_L g2164 ( 
.A1(n_1871),
.A2(n_607),
.B(n_617),
.C(n_610),
.Y(n_2164)
);

AND2x6_ASAP7_75t_SL g2165 ( 
.A(n_1920),
.B(n_610),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1895),
.B(n_1698),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2026),
.Y(n_2167)
);

INVx6_ASAP7_75t_L g2168 ( 
.A(n_1952),
.Y(n_2168)
);

NOR2xp67_ASAP7_75t_L g2169 ( 
.A(n_1942),
.B(n_1794),
.Y(n_2169)
);

NOR3xp33_ASAP7_75t_SL g2170 ( 
.A(n_1870),
.B(n_654),
.C(n_653),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1859),
.B(n_1713),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_1914),
.A2(n_1681),
.B1(n_1718),
.B2(n_1716),
.Y(n_2172)
);

BUFx10_ASAP7_75t_L g2173 ( 
.A(n_2022),
.Y(n_2173)
);

CKINVDCx14_ASAP7_75t_R g2174 ( 
.A(n_1985),
.Y(n_2174)
);

NOR3xp33_ASAP7_75t_SL g2175 ( 
.A(n_1870),
.B(n_660),
.C(n_658),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_1946),
.Y(n_2176)
);

CKINVDCx11_ASAP7_75t_R g2177 ( 
.A(n_1876),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_1988),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2002),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1913),
.A2(n_1812),
.B1(n_2006),
.B2(n_1833),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_1919),
.B(n_1569),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1859),
.B(n_1681),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_1920),
.A2(n_1803),
.B1(n_1750),
.B2(n_1759),
.Y(n_2183)
);

AOI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1904),
.A2(n_1779),
.B(n_1710),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2005),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_1952),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1932),
.B(n_1693),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1961),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2012),
.Y(n_2189)
);

OAI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1940),
.A2(n_1766),
.B(n_1692),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_1852),
.B(n_604),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1821),
.B(n_1608),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_1982),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1928),
.B(n_1746),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_R g2195 ( 
.A(n_1868),
.B(n_1714),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_1937),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_1894),
.B(n_1714),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2017),
.Y(n_2198)
);

NOR3xp33_ASAP7_75t_SL g2199 ( 
.A(n_1874),
.B(n_666),
.C(n_664),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1967),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1813),
.B(n_1925),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1925),
.B(n_1697),
.Y(n_2202)
);

BUFx4f_ASAP7_75t_SL g2203 ( 
.A(n_1962),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1992),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2015),
.B(n_1697),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2021),
.B(n_1700),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1899),
.B(n_1746),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_2023),
.Y(n_2208)
);

INVx5_ASAP7_75t_L g2209 ( 
.A(n_1873),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1968),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2018),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1969),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1845),
.B(n_1700),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1962),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_1873),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1861),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1861),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_1962),
.Y(n_2218)
);

AND2x6_ASAP7_75t_L g2219 ( 
.A(n_2004),
.B(n_1746),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1862),
.B(n_1705),
.Y(n_2220)
);

CKINVDCx14_ASAP7_75t_R g2221 ( 
.A(n_1962),
.Y(n_2221)
);

NOR3xp33_ASAP7_75t_SL g2222 ( 
.A(n_1874),
.B(n_674),
.C(n_667),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1944),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1960),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1953),
.B(n_679),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1901),
.B(n_1786),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_1974),
.B(n_1744),
.Y(n_2227)
);

BUFx4f_ASAP7_75t_L g2228 ( 
.A(n_1873),
.Y(n_2228)
);

AOI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_1912),
.A2(n_1710),
.B(n_1786),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_1894),
.B(n_1797),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1999),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1975),
.Y(n_2232)
);

AOI21x1_ASAP7_75t_L g2233 ( 
.A1(n_1889),
.A2(n_1762),
.B(n_1715),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1979),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1811),
.B(n_1705),
.Y(n_2235)
);

INVx1_ASAP7_75t_SL g2236 ( 
.A(n_1839),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1986),
.Y(n_2237)
);

BUFx3_ASAP7_75t_L g2238 ( 
.A(n_1886),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1867),
.B(n_1720),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1886),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_1840),
.B(n_1574),
.Y(n_2241)
);

OR2x6_ASAP7_75t_SL g2242 ( 
.A(n_1834),
.B(n_682),
.Y(n_2242)
);

BUFx4f_ASAP7_75t_SL g2243 ( 
.A(n_1892),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_R g2244 ( 
.A(n_1948),
.B(n_1574),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1817),
.B(n_1720),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_2019),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1892),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1853),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1817),
.B(n_1729),
.Y(n_2249)
);

NOR3xp33_ASAP7_75t_SL g2250 ( 
.A(n_1908),
.B(n_687),
.C(n_683),
.Y(n_2250)
);

BUFx2_ASAP7_75t_L g2251 ( 
.A(n_2019),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1847),
.B(n_900),
.Y(n_2252)
);

BUFx6f_ASAP7_75t_L g2253 ( 
.A(n_1831),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_1948),
.Y(n_2254)
);

AOI21x1_ASAP7_75t_L g2255 ( 
.A1(n_1889),
.A2(n_1715),
.B(n_1622),
.Y(n_2255)
);

BUFx3_ASAP7_75t_L g2256 ( 
.A(n_1856),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1877),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_1831),
.Y(n_2258)
);

BUFx2_ASAP7_75t_L g2259 ( 
.A(n_2001),
.Y(n_2259)
);

CKINVDCx20_ASAP7_75t_R g2260 ( 
.A(n_1917),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1878),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2044),
.B(n_2071),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_SL g2263 ( 
.A1(n_2027),
.A2(n_1860),
.B(n_1848),
.Y(n_2263)
);

OA22x2_ASAP7_75t_L g2264 ( 
.A1(n_2180),
.A2(n_1990),
.B1(n_2011),
.B2(n_1829),
.Y(n_2264)
);

AOI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2049),
.A2(n_1829),
.B(n_2014),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2259),
.B(n_1943),
.Y(n_2266)
);

OAI21x1_ASAP7_75t_L g2267 ( 
.A1(n_2233),
.A2(n_1931),
.B(n_1981),
.Y(n_2267)
);

AOI21xp5_ASAP7_75t_L g2268 ( 
.A1(n_2190),
.A2(n_1786),
.B(n_1740),
.Y(n_2268)
);

OAI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_2120),
.A2(n_1908),
.B(n_1887),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_2059),
.B(n_1848),
.Y(n_2270)
);

OAI21x1_ASAP7_75t_SL g2271 ( 
.A1(n_2135),
.A2(n_1882),
.B(n_1879),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2030),
.Y(n_2272)
);

O2A1O1Ixp5_ASAP7_75t_L g2273 ( 
.A1(n_2049),
.A2(n_2010),
.B(n_1980),
.C(n_1989),
.Y(n_2273)
);

NAND2x1_ASAP7_75t_L g2274 ( 
.A(n_2219),
.B(n_1760),
.Y(n_2274)
);

OAI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2027),
.A2(n_2004),
.B(n_2009),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2067),
.B(n_1935),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2184),
.A2(n_1786),
.B(n_1740),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_2177),
.Y(n_2278)
);

AOI21xp5_ASAP7_75t_L g2279 ( 
.A1(n_2184),
.A2(n_1622),
.B(n_1613),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2229),
.A2(n_2010),
.B(n_2009),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2143),
.A2(n_1613),
.B(n_1610),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2229),
.A2(n_1922),
.B(n_1976),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2067),
.B(n_2044),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2094),
.B(n_2003),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2096),
.A2(n_2097),
.B(n_2194),
.Y(n_2285)
);

AOI21x1_ASAP7_75t_L g2286 ( 
.A1(n_2255),
.A2(n_2095),
.B(n_2096),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2059),
.B(n_1938),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_SL g2288 ( 
.A(n_2228),
.B(n_1788),
.Y(n_2288)
);

OAI21x1_ASAP7_75t_L g2289 ( 
.A1(n_2095),
.A2(n_1922),
.B(n_1976),
.Y(n_2289)
);

A2O1A1Ixp33_ASAP7_75t_L g2290 ( 
.A1(n_2250),
.A2(n_1869),
.B(n_1745),
.C(n_1723),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_2053),
.Y(n_2291)
);

AO31x2_ASAP7_75t_L g2292 ( 
.A1(n_2245),
.A2(n_2249),
.A3(n_2217),
.B(n_2216),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2031),
.Y(n_2293)
);

BUFx6f_ASAP7_75t_L g2294 ( 
.A(n_2177),
.Y(n_2294)
);

BUFx2_ASAP7_75t_L g2295 ( 
.A(n_2040),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2115),
.A2(n_1733),
.B(n_1869),
.Y(n_2296)
);

AOI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2097),
.A2(n_1613),
.B(n_1610),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2223),
.B(n_1965),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2231),
.B(n_1965),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2194),
.A2(n_1613),
.B(n_1610),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2224),
.B(n_1951),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2158),
.A2(n_1628),
.B(n_1610),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2034),
.Y(n_2303)
);

AOI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2158),
.A2(n_2128),
.B(n_2207),
.Y(n_2304)
);

OAI21x1_ASAP7_75t_SL g2305 ( 
.A1(n_2183),
.A2(n_1645),
.B(n_1642),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2150),
.B(n_1951),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2207),
.A2(n_1631),
.B(n_1628),
.Y(n_2307)
);

OA21x2_ASAP7_75t_L g2308 ( 
.A1(n_2226),
.A2(n_2014),
.B(n_1989),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2028),
.B(n_2000),
.Y(n_2309)
);

AOI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2226),
.A2(n_1631),
.B(n_1628),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2048),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2038),
.Y(n_2312)
);

NAND2x1p5_ASAP7_75t_L g2313 ( 
.A(n_2228),
.B(n_1929),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2174),
.B(n_689),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2127),
.A2(n_1631),
.B(n_1628),
.Y(n_2315)
);

NAND2x1p5_ASAP7_75t_L g2316 ( 
.A(n_2072),
.B(n_1956),
.Y(n_2316)
);

AO31x2_ASAP7_75t_L g2317 ( 
.A1(n_2235),
.A2(n_1761),
.A3(n_1781),
.B(n_1729),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_2040),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2063),
.B(n_1917),
.Y(n_2319)
);

OAI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2101),
.A2(n_1995),
.B(n_1980),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2032),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2033),
.A2(n_618),
.B1(n_624),
.B2(n_617),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2094),
.B(n_1761),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2127),
.A2(n_1636),
.B(n_1631),
.Y(n_2324)
);

AOI21xp33_ASAP7_75t_L g2325 ( 
.A1(n_2172),
.A2(n_1766),
.B(n_1995),
.Y(n_2325)
);

O2A1O1Ixp33_ASAP7_75t_L g2326 ( 
.A1(n_2108),
.A2(n_624),
.B(n_627),
.C(n_618),
.Y(n_2326)
);

BUFx4_ASAP7_75t_R g2327 ( 
.A(n_2058),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2041),
.Y(n_2328)
);

OAI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2108),
.A2(n_2000),
.B(n_1998),
.Y(n_2329)
);

OAI21x1_ASAP7_75t_L g2330 ( 
.A1(n_2101),
.A2(n_2007),
.B(n_1998),
.Y(n_2330)
);

OAI21x1_ASAP7_75t_L g2331 ( 
.A1(n_2215),
.A2(n_2008),
.B(n_2007),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_2174),
.B(n_690),
.Y(n_2332)
);

AOI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_2046),
.A2(n_1666),
.B(n_1636),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2070),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2125),
.B(n_691),
.Y(n_2335)
);

OAI21x1_ASAP7_75t_L g2336 ( 
.A1(n_2215),
.A2(n_2008),
.B(n_1938),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2046),
.A2(n_1666),
.B(n_1636),
.Y(n_2337)
);

INVx2_ASAP7_75t_SL g2338 ( 
.A(n_2173),
.Y(n_2338)
);

INVx4_ASAP7_75t_L g2339 ( 
.A(n_2203),
.Y(n_2339)
);

AO31x2_ASAP7_75t_L g2340 ( 
.A1(n_2192),
.A2(n_1781),
.A3(n_1808),
.B(n_1790),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2213),
.A2(n_1666),
.B(n_1636),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2079),
.Y(n_2342)
);

OAI21x1_ASAP7_75t_L g2343 ( 
.A1(n_2077),
.A2(n_1956),
.B(n_1929),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_L g2344 ( 
.A(n_2164),
.B(n_628),
.C(n_627),
.Y(n_2344)
);

INVx3_ASAP7_75t_L g2345 ( 
.A(n_2032),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2045),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2167),
.B(n_1790),
.Y(n_2347)
);

BUFx2_ASAP7_75t_L g2348 ( 
.A(n_2070),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2063),
.B(n_1957),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2126),
.B(n_628),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2050),
.Y(n_2351)
);

NAND3xp33_ASAP7_75t_L g2352 ( 
.A(n_2250),
.B(n_655),
.C(n_647),
.Y(n_2352)
);

NAND2x1p5_ASAP7_75t_L g2353 ( 
.A(n_2072),
.B(n_1963),
.Y(n_2353)
);

BUFx6f_ASAP7_75t_L g2354 ( 
.A(n_2032),
.Y(n_2354)
);

OAI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2077),
.A2(n_1963),
.B(n_1957),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2240),
.A2(n_1735),
.B(n_1709),
.Y(n_2356)
);

AOI21x1_ASAP7_75t_L g2357 ( 
.A1(n_2169),
.A2(n_1497),
.B(n_1495),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2054),
.B(n_2134),
.Y(n_2358)
);

OAI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_2252),
.A2(n_1447),
.B(n_1667),
.Y(n_2359)
);

AOI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2182),
.A2(n_1685),
.B(n_1666),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2060),
.A2(n_1685),
.B(n_1723),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2188),
.B(n_1808),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2200),
.B(n_1748),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2130),
.B(n_647),
.Y(n_2364)
);

INVxp67_ASAP7_75t_L g2365 ( 
.A(n_2124),
.Y(n_2365)
);

A2O1A1Ixp33_ASAP7_75t_L g2366 ( 
.A1(n_2033),
.A2(n_1745),
.B(n_656),
.C(n_671),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2081),
.Y(n_2367)
);

OAI21x1_ASAP7_75t_L g2368 ( 
.A1(n_2240),
.A2(n_2192),
.B(n_2248),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2210),
.B(n_1799),
.Y(n_2369)
);

OAI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2257),
.A2(n_1735),
.B(n_1709),
.Y(n_2370)
);

OAI21x1_ASAP7_75t_L g2371 ( 
.A1(n_2187),
.A2(n_1810),
.B(n_1428),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2056),
.Y(n_2372)
);

NOR2x1_ASAP7_75t_L g2373 ( 
.A(n_2091),
.B(n_1675),
.Y(n_2373)
);

BUFx2_ASAP7_75t_L g2374 ( 
.A(n_2091),
.Y(n_2374)
);

OAI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2172),
.A2(n_1678),
.B(n_1810),
.Y(n_2375)
);

AOI21x1_ASAP7_75t_L g2376 ( 
.A1(n_2239),
.A2(n_1531),
.B(n_1497),
.Y(n_2376)
);

OAI21x1_ASAP7_75t_L g2377 ( 
.A1(n_2261),
.A2(n_1428),
.B(n_1424),
.Y(n_2377)
);

AOI21xp33_ASAP7_75t_L g2378 ( 
.A1(n_2201),
.A2(n_1389),
.B(n_1433),
.Y(n_2378)
);

OAI21x1_ASAP7_75t_L g2379 ( 
.A1(n_2220),
.A2(n_1435),
.B(n_1433),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2068),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2212),
.B(n_1685),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_2061),
.B(n_1685),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2105),
.A2(n_1425),
.B(n_1760),
.Y(n_2383)
);

OAI21x1_ASAP7_75t_L g2384 ( 
.A1(n_2205),
.A2(n_1436),
.B(n_1435),
.Y(n_2384)
);

OAI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2029),
.A2(n_1770),
.B(n_1760),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2202),
.A2(n_1425),
.B(n_1760),
.Y(n_2386)
);

O2A1O1Ixp5_ASAP7_75t_L g2387 ( 
.A1(n_2230),
.A2(n_1550),
.B(n_1556),
.C(n_1531),
.Y(n_2387)
);

OAI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2206),
.A2(n_1461),
.B(n_1436),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2208),
.A2(n_697),
.B1(n_706),
.B2(n_696),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_SL g2390 ( 
.A1(n_2171),
.A2(n_714),
.B(n_665),
.Y(n_2390)
);

AOI21x1_ASAP7_75t_L g2391 ( 
.A1(n_2251),
.A2(n_1556),
.B(n_1550),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2152),
.A2(n_1770),
.B(n_1760),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2088),
.B(n_1589),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2088),
.B(n_1589),
.Y(n_2394)
);

OAI21x1_ASAP7_75t_L g2395 ( 
.A1(n_2078),
.A2(n_1466),
.B(n_1461),
.Y(n_2395)
);

NAND2x1_ASAP7_75t_L g2396 ( 
.A(n_2219),
.B(n_1770),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2155),
.A2(n_1770),
.B(n_1699),
.Y(n_2397)
);

OAI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2225),
.A2(n_1770),
.B(n_1699),
.Y(n_2398)
);

AOI21xp33_ASAP7_75t_L g2399 ( 
.A1(n_2196),
.A2(n_1474),
.B(n_1466),
.Y(n_2399)
);

AOI21xp33_ASAP7_75t_L g2400 ( 
.A1(n_2196),
.A2(n_1475),
.B(n_1474),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2037),
.Y(n_2401)
);

AND2x6_ASAP7_75t_L g2402 ( 
.A(n_2254),
.B(n_1788),
.Y(n_2402)
);

OAI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2170),
.A2(n_1535),
.B(n_1476),
.Y(n_2403)
);

NAND2x1p5_ASAP7_75t_L g2404 ( 
.A(n_2072),
.B(n_1475),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2073),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2037),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2098),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2107),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2055),
.A2(n_656),
.B1(n_671),
.B2(n_655),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2080),
.B(n_701),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2162),
.B(n_678),
.Y(n_2411)
);

OAI21x1_ASAP7_75t_L g2412 ( 
.A1(n_2078),
.A2(n_1534),
.B(n_1476),
.Y(n_2412)
);

OAI21x1_ASAP7_75t_L g2413 ( 
.A1(n_2109),
.A2(n_1537),
.B(n_1534),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2104),
.A2(n_710),
.B1(n_713),
.B2(n_709),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2109),
.A2(n_1539),
.B(n_1537),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2035),
.A2(n_1402),
.B(n_1394),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2204),
.B(n_678),
.Y(n_2417)
);

BUFx12f_ASAP7_75t_L g2418 ( 
.A(n_2074),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2139),
.B(n_1539),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2028),
.A2(n_2052),
.B1(n_2175),
.B2(n_2170),
.Y(n_2420)
);

A2O1A1Ixp33_ASAP7_75t_L g2421 ( 
.A1(n_2175),
.A2(n_686),
.B(n_693),
.C(n_681),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2113),
.B(n_681),
.Y(n_2422)
);

OAI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2052),
.A2(n_1548),
.B(n_1402),
.Y(n_2423)
);

CKINVDCx20_ASAP7_75t_R g2424 ( 
.A(n_2051),
.Y(n_2424)
);

AOI21xp33_ASAP7_75t_L g2425 ( 
.A1(n_2191),
.A2(n_1548),
.B(n_693),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2035),
.A2(n_1403),
.B(n_1394),
.Y(n_2426)
);

NAND2x1_ASAP7_75t_L g2427 ( 
.A(n_2219),
.B(n_1305),
.Y(n_2427)
);

INVx2_ASAP7_75t_SL g2428 ( 
.A(n_2173),
.Y(n_2428)
);

OAI21xp5_ASAP7_75t_L g2429 ( 
.A1(n_2104),
.A2(n_1403),
.B(n_694),
.Y(n_2429)
);

NOR2xp67_ASAP7_75t_L g2430 ( 
.A(n_2043),
.B(n_1305),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2204),
.B(n_1300),
.Y(n_2431)
);

OAI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2106),
.A2(n_694),
.B(n_686),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_2037),
.Y(n_2433)
);

INVx2_ASAP7_75t_SL g2434 ( 
.A(n_2100),
.Y(n_2434)
);

OAI21x1_ASAP7_75t_L g2435 ( 
.A1(n_2254),
.A2(n_1305),
.B(n_1303),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2076),
.Y(n_2436)
);

OAI21x1_ASAP7_75t_L g2437 ( 
.A1(n_2154),
.A2(n_1303),
.B(n_1300),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2106),
.A2(n_703),
.B(n_695),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2035),
.A2(n_1241),
.B(n_1257),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2234),
.B(n_1311),
.Y(n_2440)
);

AOI21xp5_ASAP7_75t_L g2441 ( 
.A1(n_2072),
.A2(n_1241),
.B(n_1257),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2256),
.B(n_1311),
.Y(n_2442)
);

OAI21x1_ASAP7_75t_L g2443 ( 
.A1(n_2154),
.A2(n_965),
.B(n_964),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_2244),
.B(n_1257),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2102),
.A2(n_1241),
.B(n_1257),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2256),
.B(n_848),
.Y(n_2446)
);

OAI21x1_ASAP7_75t_L g2447 ( 
.A1(n_2193),
.A2(n_965),
.B(n_964),
.Y(n_2447)
);

AO21x1_ASAP7_75t_L g2448 ( 
.A1(n_2147),
.A2(n_703),
.B(n_695),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2193),
.A2(n_965),
.B(n_964),
.Y(n_2449)
);

OAI21x1_ASAP7_75t_L g2450 ( 
.A1(n_2082),
.A2(n_992),
.B(n_975),
.Y(n_2450)
);

OAI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2199),
.A2(n_711),
.B(n_708),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2244),
.B(n_1283),
.Y(n_2452)
);

BUFx12f_ASAP7_75t_L g2453 ( 
.A(n_2136),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2083),
.Y(n_2454)
);

OAI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2199),
.A2(n_711),
.B(n_708),
.Y(n_2455)
);

INVx5_ASAP7_75t_L g2456 ( 
.A(n_2102),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2110),
.A2(n_712),
.B1(n_722),
.B2(n_715),
.Y(n_2457)
);

OAI21x1_ASAP7_75t_L g2458 ( 
.A1(n_2084),
.A2(n_992),
.B(n_975),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2113),
.B(n_712),
.Y(n_2459)
);

OAI21x1_ASAP7_75t_L g2460 ( 
.A1(n_2092),
.A2(n_992),
.B(n_975),
.Y(n_2460)
);

OAI21x1_ASAP7_75t_L g2461 ( 
.A1(n_2117),
.A2(n_848),
.B(n_831),
.Y(n_2461)
);

OAI22x1_ASAP7_75t_L g2462 ( 
.A1(n_2163),
.A2(n_722),
.B1(n_723),
.B2(n_715),
.Y(n_2462)
);

OAI21x1_ASAP7_75t_L g2463 ( 
.A1(n_2123),
.A2(n_832),
.B(n_830),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2161),
.B(n_723),
.Y(n_2464)
);

OAI21x1_ASAP7_75t_L g2465 ( 
.A1(n_2129),
.A2(n_833),
.B(n_832),
.Y(n_2465)
);

AOI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2102),
.A2(n_1241),
.B(n_1283),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2243),
.B(n_1283),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2232),
.B(n_740),
.Y(n_2468)
);

OAI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2222),
.A2(n_755),
.B(n_740),
.Y(n_2469)
);

O2A1O1Ixp5_ASAP7_75t_L g2470 ( 
.A1(n_2230),
.A2(n_759),
.B(n_765),
.C(n_755),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2237),
.B(n_759),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2102),
.A2(n_2209),
.B(n_2142),
.Y(n_2472)
);

OAI21x1_ASAP7_75t_L g2473 ( 
.A1(n_2131),
.A2(n_836),
.B(n_833),
.Y(n_2473)
);

OAI21x1_ASAP7_75t_L g2474 ( 
.A1(n_2133),
.A2(n_839),
.B(n_836),
.Y(n_2474)
);

OAI21x1_ASAP7_75t_L g2475 ( 
.A1(n_2137),
.A2(n_840),
.B(n_839),
.Y(n_2475)
);

OAI21xp33_ASAP7_75t_L g2476 ( 
.A1(n_2161),
.A2(n_2114),
.B(n_2222),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2036),
.Y(n_2477)
);

AOI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2142),
.A2(n_1241),
.B(n_1283),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2166),
.B(n_765),
.Y(n_2479)
);

O2A1O1Ixp5_ASAP7_75t_L g2480 ( 
.A1(n_2064),
.A2(n_773),
.B(n_787),
.C(n_771),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2144),
.B(n_2145),
.Y(n_2481)
);

AOI21x1_ASAP7_75t_L g2482 ( 
.A1(n_2160),
.A2(n_773),
.B(n_771),
.Y(n_2482)
);

OAI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2219),
.A2(n_794),
.B(n_787),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2243),
.B(n_1006),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2036),
.Y(n_2485)
);

AND3x4_ASAP7_75t_L g2486 ( 
.A(n_2085),
.B(n_736),
.C(n_735),
.Y(n_2486)
);

AOI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2058),
.A2(n_717),
.B1(n_719),
.B2(n_716),
.Y(n_2487)
);

AOI21x1_ASAP7_75t_L g2488 ( 
.A1(n_2160),
.A2(n_795),
.B(n_794),
.Y(n_2488)
);

AOI22xp33_ASAP7_75t_L g2489 ( 
.A1(n_2153),
.A2(n_2236),
.B1(n_2181),
.B2(n_2119),
.Y(n_2489)
);

INVx3_ASAP7_75t_L g2490 ( 
.A(n_2066),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2219),
.B(n_2147),
.Y(n_2491)
);

OA21x2_ASAP7_75t_L g2492 ( 
.A1(n_2122),
.A2(n_2146),
.B(n_2140),
.Y(n_2492)
);

OR2x6_ASAP7_75t_L g2493 ( 
.A(n_2253),
.B(n_2258),
.Y(n_2493)
);

AOI21x1_ASAP7_75t_L g2494 ( 
.A1(n_2246),
.A2(n_798),
.B(n_795),
.Y(n_2494)
);

AND3x4_ASAP7_75t_L g2495 ( 
.A(n_2085),
.B(n_2065),
.C(n_2062),
.Y(n_2495)
);

AOI21xp5_ASAP7_75t_L g2496 ( 
.A1(n_2142),
.A2(n_2209),
.B(n_2197),
.Y(n_2496)
);

A2O1A1Ixp33_ASAP7_75t_L g2497 ( 
.A1(n_2114),
.A2(n_801),
.B(n_803),
.C(n_798),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2142),
.A2(n_736),
.B(n_735),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2149),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2209),
.A2(n_739),
.B(n_801),
.Y(n_2500)
);

NAND2xp33_ASAP7_75t_L g2501 ( 
.A(n_2042),
.B(n_725),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2062),
.B(n_803),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2227),
.B(n_805),
.Y(n_2503)
);

HB1xp67_ASAP7_75t_L g2504 ( 
.A(n_2221),
.Y(n_2504)
);

OAI21x1_ASAP7_75t_L g2505 ( 
.A1(n_2151),
.A2(n_841),
.B(n_840),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2042),
.Y(n_2506)
);

AOI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2241),
.A2(n_805),
.B(n_841),
.Y(n_2507)
);

OAI21x1_ASAP7_75t_L g2508 ( 
.A1(n_2159),
.A2(n_844),
.B(n_843),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2209),
.A2(n_2197),
.B(n_2221),
.Y(n_2509)
);

A2O1A1Ixp33_ASAP7_75t_L g2510 ( 
.A1(n_2039),
.A2(n_739),
.B(n_727),
.C(n_728),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2179),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2139),
.B(n_1006),
.Y(n_2512)
);

OAI21xp33_ASAP7_75t_L g2513 ( 
.A1(n_2065),
.A2(n_730),
.B(n_726),
.Y(n_2513)
);

OAI21xp5_ASAP7_75t_L g2514 ( 
.A1(n_2241),
.A2(n_844),
.B(n_843),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2039),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2118),
.A2(n_778),
.B(n_661),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2141),
.B(n_731),
.Y(n_2517)
);

AOI21xp5_ASAP7_75t_L g2518 ( 
.A1(n_2118),
.A2(n_778),
.B(n_661),
.Y(n_2518)
);

AO31x2_ASAP7_75t_L g2519 ( 
.A1(n_2185),
.A2(n_847),
.A3(n_1040),
.B(n_1026),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2189),
.Y(n_2520)
);

OAI21x1_ASAP7_75t_L g2521 ( 
.A1(n_2198),
.A2(n_847),
.B(n_1006),
.Y(n_2521)
);

OA21x2_ASAP7_75t_L g2522 ( 
.A1(n_2211),
.A2(n_512),
.B(n_506),
.Y(n_2522)
);

OAI21xp33_ASAP7_75t_L g2523 ( 
.A1(n_2086),
.A2(n_734),
.B(n_732),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2090),
.B(n_737),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2047),
.A2(n_743),
.B(n_745),
.C(n_741),
.Y(n_2525)
);

OAI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2260),
.A2(n_747),
.B1(n_748),
.B2(n_746),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_L g2527 ( 
.A1(n_2118),
.A2(n_778),
.B(n_1006),
.Y(n_2527)
);

INVxp67_ASAP7_75t_L g2528 ( 
.A(n_2176),
.Y(n_2528)
);

AO31x2_ASAP7_75t_L g2529 ( 
.A1(n_2064),
.A2(n_1040),
.A3(n_1026),
.B(n_663),
.Y(n_2529)
);

AOI21xp33_ASAP7_75t_L g2530 ( 
.A1(n_2253),
.A2(n_752),
.B(n_749),
.Y(n_2530)
);

BUFx12f_ASAP7_75t_L g2531 ( 
.A(n_2453),
.Y(n_2531)
);

INVx3_ASAP7_75t_SL g2532 ( 
.A(n_2506),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2277),
.A2(n_2279),
.B(n_2268),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2283),
.B(n_2075),
.Y(n_2534)
);

INVx1_ASAP7_75t_SL g2535 ( 
.A(n_2334),
.Y(n_2535)
);

AOI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2392),
.A2(n_2121),
.B(n_2118),
.Y(n_2536)
);

AOI22xp33_ASAP7_75t_L g2537 ( 
.A1(n_2322),
.A2(n_2148),
.B1(n_663),
.B2(n_673),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2477),
.Y(n_2538)
);

BUFx6f_ASAP7_75t_L g2539 ( 
.A(n_2477),
.Y(n_2539)
);

BUFx10_ASAP7_75t_L g2540 ( 
.A(n_2517),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2276),
.B(n_2247),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2314),
.B(n_2141),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2293),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2321),
.B(n_2247),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2358),
.B(n_2069),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2278),
.B(n_2218),
.Y(n_2546)
);

BUFx6f_ASAP7_75t_L g2547 ( 
.A(n_2477),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2272),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2309),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2303),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2312),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2278),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2278),
.B(n_2294),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2348),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2321),
.Y(n_2555)
);

AOI21xp33_ASAP7_75t_SL g2556 ( 
.A1(n_2495),
.A2(n_2434),
.B(n_2420),
.Y(n_2556)
);

OAI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_2264),
.A2(n_2242),
.B1(n_2156),
.B2(n_2138),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2281),
.A2(n_2263),
.B(n_2385),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2374),
.Y(n_2559)
);

INVx1_ASAP7_75t_SL g2560 ( 
.A(n_2291),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2291),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2328),
.Y(n_2562)
);

OR2x6_ASAP7_75t_L g2563 ( 
.A(n_2274),
.B(n_2253),
.Y(n_2563)
);

BUFx6f_ASAP7_75t_L g2564 ( 
.A(n_2485),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2284),
.B(n_2247),
.Y(n_2565)
);

INVx5_ASAP7_75t_L g2566 ( 
.A(n_2456),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2294),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2346),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2321),
.B(n_2247),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2485),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2354),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2294),
.Y(n_2572)
);

BUFx6f_ASAP7_75t_L g2573 ( 
.A(n_2485),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2311),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2351),
.Y(n_2575)
);

OR2x6_ASAP7_75t_L g2576 ( 
.A(n_2396),
.B(n_2253),
.Y(n_2576)
);

OAI22xp33_ASAP7_75t_SL g2577 ( 
.A1(n_2322),
.A2(n_2178),
.B1(n_2168),
.B2(n_2165),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_SL g2578 ( 
.A(n_2456),
.B(n_2156),
.Y(n_2578)
);

BUFx2_ASAP7_75t_L g2579 ( 
.A(n_2504),
.Y(n_2579)
);

INVx5_ASAP7_75t_L g2580 ( 
.A(n_2456),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2264),
.A2(n_663),
.B1(n_673),
.B2(n_2111),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_2515),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2342),
.Y(n_2583)
);

AOI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2332),
.A2(n_2168),
.B1(n_2138),
.B2(n_2069),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2367),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2372),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2266),
.B(n_2214),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2266),
.B(n_2218),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2262),
.B(n_2121),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2407),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2408),
.Y(n_2591)
);

AOI22xp33_ASAP7_75t_SL g2592 ( 
.A1(n_2409),
.A2(n_2258),
.B1(n_2168),
.B2(n_763),
.Y(n_2592)
);

BUFx3_ASAP7_75t_L g2593 ( 
.A(n_2318),
.Y(n_2593)
);

INVx4_ASAP7_75t_L g2594 ( 
.A(n_2339),
.Y(n_2594)
);

AOI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2385),
.A2(n_2132),
.B(n_2121),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2515),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2481),
.B(n_2116),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2491),
.B(n_2258),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2476),
.A2(n_2186),
.B1(n_2258),
.B2(n_2057),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2380),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2354),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2405),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2304),
.B(n_2323),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2511),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2354),
.B(n_2066),
.Y(n_2605)
);

CKINVDCx20_ASAP7_75t_R g2606 ( 
.A(n_2424),
.Y(n_2606)
);

BUFx3_ASAP7_75t_L g2607 ( 
.A(n_2418),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2436),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2454),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2422),
.B(n_2121),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2499),
.Y(n_2611)
);

NAND2x1p5_ASAP7_75t_L g2612 ( 
.A(n_2456),
.B(n_2057),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2491),
.B(n_2066),
.Y(n_2613)
);

BUFx6f_ASAP7_75t_L g2614 ( 
.A(n_2515),
.Y(n_2614)
);

AND2x4_ASAP7_75t_L g2615 ( 
.A(n_2493),
.B(n_2066),
.Y(n_2615)
);

INVx4_ASAP7_75t_SL g2616 ( 
.A(n_2402),
.Y(n_2616)
);

NOR2xp67_ASAP7_75t_L g2617 ( 
.A(n_2338),
.B(n_2087),
.Y(n_2617)
);

BUFx2_ASAP7_75t_L g2618 ( 
.A(n_2365),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2520),
.Y(n_2619)
);

INVx2_ASAP7_75t_SL g2620 ( 
.A(n_2295),
.Y(n_2620)
);

AOI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2425),
.A2(n_663),
.B1(n_673),
.B2(n_2238),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2428),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2292),
.Y(n_2623)
);

CKINVDCx11_ASAP7_75t_R g2624 ( 
.A(n_2406),
.Y(n_2624)
);

CKINVDCx20_ASAP7_75t_R g2625 ( 
.A(n_2528),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2285),
.B(n_2132),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2306),
.B(n_2132),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2389),
.A2(n_766),
.B1(n_767),
.B2(n_757),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2292),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2492),
.Y(n_2630)
);

OAI21x1_ASAP7_75t_L g2631 ( 
.A1(n_2267),
.A2(n_2103),
.B(n_2203),
.Y(n_2631)
);

BUFx3_ASAP7_75t_L g2632 ( 
.A(n_2459),
.Y(n_2632)
);

BUFx12f_ASAP7_75t_L g2633 ( 
.A(n_2339),
.Y(n_2633)
);

NAND2x1p5_ASAP7_75t_L g2634 ( 
.A(n_2444),
.B(n_2089),
.Y(n_2634)
);

BUFx3_ASAP7_75t_L g2635 ( 
.A(n_2406),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2493),
.B(n_2089),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2292),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2406),
.Y(n_2638)
);

INVxp67_ASAP7_75t_L g2639 ( 
.A(n_2308),
.Y(n_2639)
);

OAI21x1_ASAP7_75t_L g2640 ( 
.A1(n_2376),
.A2(n_2103),
.B(n_2132),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2433),
.Y(n_2641)
);

NAND2xp33_ASAP7_75t_L g2642 ( 
.A(n_2290),
.B(n_2157),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2493),
.B(n_2089),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_2410),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2431),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2433),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_L g2647 ( 
.A1(n_2425),
.A2(n_1030),
.B1(n_1041),
.B2(n_1006),
.Y(n_2647)
);

OAI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2275),
.A2(n_2087),
.B(n_774),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2306),
.B(n_2089),
.Y(n_2649)
);

BUFx4_ASAP7_75t_SL g2650 ( 
.A(n_2344),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2393),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2431),
.Y(n_2652)
);

INVx1_ASAP7_75t_SL g2653 ( 
.A(n_2393),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2394),
.Y(n_2654)
);

BUFx5_ASAP7_75t_L g2655 ( 
.A(n_2402),
.Y(n_2655)
);

CKINVDCx16_ASAP7_75t_R g2656 ( 
.A(n_2524),
.Y(n_2656)
);

INVx5_ASAP7_75t_L g2657 ( 
.A(n_2402),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2433),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2335),
.Y(n_2659)
);

O2A1O1Ixp33_ASAP7_75t_L g2660 ( 
.A1(n_2366),
.A2(n_776),
.B(n_777),
.C(n_768),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2301),
.B(n_2093),
.Y(n_2661)
);

AND2x2_ASAP7_75t_SL g2662 ( 
.A(n_2288),
.B(n_2093),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2409),
.A2(n_783),
.B1(n_784),
.B2(n_781),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2394),
.Y(n_2664)
);

AO21x2_ASAP7_75t_L g2665 ( 
.A1(n_2296),
.A2(n_2099),
.B(n_2086),
.Y(n_2665)
);

OR2x6_ASAP7_75t_L g2666 ( 
.A(n_2472),
.B(n_2093),
.Y(n_2666)
);

INVxp67_ASAP7_75t_L g2667 ( 
.A(n_2308),
.Y(n_2667)
);

AOI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2275),
.A2(n_2112),
.B(n_2093),
.Y(n_2668)
);

INVx4_ASAP7_75t_L g2669 ( 
.A(n_2327),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2492),
.Y(n_2670)
);

BUFx6f_ASAP7_75t_L g2671 ( 
.A(n_2287),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2490),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_L g2673 ( 
.A1(n_2502),
.A2(n_1030),
.B1(n_1042),
.B2(n_1041),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2317),
.Y(n_2674)
);

BUFx6f_ASAP7_75t_L g2675 ( 
.A(n_2287),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2364),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2319),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2350),
.B(n_2112),
.Y(n_2678)
);

AOI221x1_ASAP7_75t_L g2679 ( 
.A1(n_2420),
.A2(n_2112),
.B1(n_778),
.B2(n_1041),
.C(n_1042),
.Y(n_2679)
);

INVx5_ASAP7_75t_L g2680 ( 
.A(n_2402),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2301),
.B(n_2112),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_R g2682 ( 
.A(n_2501),
.B(n_518),
.Y(n_2682)
);

BUFx10_ASAP7_75t_L g2683 ( 
.A(n_2512),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2486),
.A2(n_788),
.B1(n_790),
.B2(n_786),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2368),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2317),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2483),
.A2(n_796),
.B1(n_797),
.B2(n_792),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2269),
.B(n_2099),
.Y(n_2688)
);

INVxp67_ASAP7_75t_SL g2689 ( 
.A(n_2381),
.Y(n_2689)
);

INVx5_ASAP7_75t_L g2690 ( 
.A(n_2345),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2317),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2345),
.B(n_1030),
.Y(n_2692)
);

BUFx3_ASAP7_75t_L g2693 ( 
.A(n_2319),
.Y(n_2693)
);

INVx2_ASAP7_75t_SL g2694 ( 
.A(n_2490),
.Y(n_2694)
);

INVx3_ASAP7_75t_SL g2695 ( 
.A(n_2349),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2401),
.B(n_1030),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2464),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2349),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2432),
.B(n_0),
.Y(n_2699)
);

INVx3_ASAP7_75t_L g2700 ( 
.A(n_2401),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2432),
.B(n_2),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2269),
.B(n_2157),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2438),
.A2(n_800),
.B1(n_809),
.B2(n_807),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2438),
.B(n_3),
.Y(n_2704)
);

BUFx6f_ASAP7_75t_L g2705 ( 
.A(n_2270),
.Y(n_2705)
);

AND2x4_ASAP7_75t_L g2706 ( 
.A(n_2270),
.B(n_1030),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2417),
.B(n_3),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_SL g2708 ( 
.A(n_2483),
.B(n_2195),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2347),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2347),
.Y(n_2710)
);

BUFx12f_ASAP7_75t_L g2711 ( 
.A(n_2512),
.Y(n_2711)
);

BUFx2_ASAP7_75t_L g2712 ( 
.A(n_2398),
.Y(n_2712)
);

INVx1_ASAP7_75t_SL g2713 ( 
.A(n_2373),
.Y(n_2713)
);

BUFx5_ASAP7_75t_L g2714 ( 
.A(n_2419),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2398),
.B(n_4),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_2526),
.B(n_6),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2362),
.Y(n_2717)
);

NOR3xp33_ASAP7_75t_L g2718 ( 
.A(n_2421),
.B(n_521),
.C(n_520),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2381),
.Y(n_2719)
);

OAI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2414),
.A2(n_2195),
.B1(n_778),
.B2(n_10),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2362),
.Y(n_2721)
);

INVxp67_ASAP7_75t_SL g2722 ( 
.A(n_2442),
.Y(n_2722)
);

CKINVDCx16_ASAP7_75t_R g2723 ( 
.A(n_2288),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2363),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2363),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2369),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2489),
.Y(n_2727)
);

BUFx10_ASAP7_75t_L g2728 ( 
.A(n_2419),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2296),
.B(n_1030),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2462),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2369),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2340),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2313),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2522),
.A2(n_1042),
.B1(n_1043),
.B2(n_1041),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2340),
.Y(n_2735)
);

AOI22xp33_ASAP7_75t_L g2736 ( 
.A1(n_2522),
.A2(n_1042),
.B1(n_1043),
.B2(n_1041),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2340),
.Y(n_2737)
);

AND2x4_ASAP7_75t_L g2738 ( 
.A(n_2509),
.B(n_1041),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2446),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2427),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2446),
.Y(n_2741)
);

A2O1A1Ixp33_ASAP7_75t_SL g2742 ( 
.A1(n_2451),
.A2(n_11),
.B(n_7),
.C(n_8),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2298),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2442),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2379),
.Y(n_2745)
);

INVx3_ASAP7_75t_L g2746 ( 
.A(n_2336),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2429),
.B(n_8),
.Y(n_2747)
);

HB1xp67_ASAP7_75t_L g2748 ( 
.A(n_2265),
.Y(n_2748)
);

AOI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2386),
.A2(n_1043),
.B(n_1042),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2298),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2448),
.A2(n_1043),
.B1(n_1046),
.B2(n_1042),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2299),
.Y(n_2752)
);

AOI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_2382),
.A2(n_537),
.B1(n_547),
.B2(n_529),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2299),
.Y(n_2754)
);

BUFx3_ASAP7_75t_L g2755 ( 
.A(n_2313),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2343),
.Y(n_2756)
);

BUFx2_ASAP7_75t_SL g2757 ( 
.A(n_2430),
.Y(n_2757)
);

OAI21x1_ASAP7_75t_L g2758 ( 
.A1(n_2384),
.A2(n_1046),
.B(n_1043),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2388),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2320),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_2316),
.Y(n_2761)
);

INVx8_ASAP7_75t_L g2762 ( 
.A(n_2496),
.Y(n_2762)
);

OR2x2_ASAP7_75t_L g2763 ( 
.A(n_2503),
.B(n_1043),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2355),
.B(n_1046),
.Y(n_2764)
);

INVx8_ASAP7_75t_L g2765 ( 
.A(n_2467),
.Y(n_2765)
);

BUFx5_ASAP7_75t_L g2766 ( 
.A(n_2273),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2440),
.Y(n_2767)
);

A2O1A1Ixp33_ASAP7_75t_L g2768 ( 
.A1(n_2510),
.A2(n_2497),
.B(n_2523),
.C(n_2326),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2397),
.A2(n_1051),
.B(n_1046),
.Y(n_2769)
);

AOI221xp5_ASAP7_75t_L g2770 ( 
.A1(n_2457),
.A2(n_591),
.B1(n_602),
.B2(n_587),
.C(n_581),
.Y(n_2770)
);

NAND3xp33_ASAP7_75t_L g2771 ( 
.A(n_2352),
.B(n_1051),
.C(n_1046),
.Y(n_2771)
);

BUFx4f_ASAP7_75t_SL g2772 ( 
.A(n_2484),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2503),
.B(n_1046),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2468),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2383),
.A2(n_1056),
.B(n_1051),
.Y(n_2775)
);

INVx4_ASAP7_75t_L g2776 ( 
.A(n_2316),
.Y(n_2776)
);

BUFx2_ASAP7_75t_L g2777 ( 
.A(n_2353),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2330),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2429),
.B(n_11),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2353),
.Y(n_2780)
);

BUFx2_ASAP7_75t_L g2781 ( 
.A(n_2329),
.Y(n_2781)
);

BUFx2_ASAP7_75t_L g2782 ( 
.A(n_2329),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_2479),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2440),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2526),
.A2(n_606),
.B1(n_615),
.B2(n_613),
.Y(n_2785)
);

NOR3xp33_ASAP7_75t_L g2786 ( 
.A(n_2451),
.B(n_619),
.C(n_616),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2271),
.B(n_1051),
.Y(n_2787)
);

INVx3_ASAP7_75t_L g2788 ( 
.A(n_2331),
.Y(n_2788)
);

INVx1_ASAP7_75t_SL g2789 ( 
.A(n_2452),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2423),
.B(n_1051),
.Y(n_2790)
);

BUFx3_ASAP7_75t_L g2791 ( 
.A(n_2606),
.Y(n_2791)
);

OAI21x1_ASAP7_75t_L g2792 ( 
.A1(n_2749),
.A2(n_2286),
.B(n_2282),
.Y(n_2792)
);

OAI21x1_ASAP7_75t_L g2793 ( 
.A1(n_2749),
.A2(n_2280),
.B(n_2289),
.Y(n_2793)
);

HB1xp67_ASAP7_75t_L g2794 ( 
.A(n_2639),
.Y(n_2794)
);

OAI21x1_ASAP7_75t_L g2795 ( 
.A1(n_2775),
.A2(n_2371),
.B(n_2435),
.Y(n_2795)
);

OA21x2_ASAP7_75t_L g2796 ( 
.A1(n_2639),
.A2(n_2667),
.B(n_2629),
.Y(n_2796)
);

OAI21x1_ASAP7_75t_L g2797 ( 
.A1(n_2775),
.A2(n_2769),
.B(n_2758),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2543),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2611),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2662),
.Y(n_2800)
);

OAI21x1_ASAP7_75t_L g2801 ( 
.A1(n_2769),
.A2(n_2310),
.B(n_2307),
.Y(n_2801)
);

AOI21xp33_ASAP7_75t_SL g2802 ( 
.A1(n_2532),
.A2(n_2469),
.B(n_2455),
.Y(n_2802)
);

OAI22xp5_ASAP7_75t_SL g2803 ( 
.A1(n_2669),
.A2(n_2469),
.B1(n_2455),
.B2(n_2457),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2550),
.Y(n_2804)
);

CKINVDCx6p67_ASAP7_75t_R g2805 ( 
.A(n_2531),
.Y(n_2805)
);

BUFx12f_ASAP7_75t_L g2806 ( 
.A(n_2540),
.Y(n_2806)
);

AO32x2_ASAP7_75t_L g2807 ( 
.A1(n_2694),
.A2(n_2390),
.A3(n_2423),
.B1(n_2325),
.B2(n_2387),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2603),
.B(n_2411),
.Y(n_2808)
);

O2A1O1Ixp33_ASAP7_75t_L g2809 ( 
.A1(n_2768),
.A2(n_2525),
.B(n_2530),
.C(n_2470),
.Y(n_2809)
);

O2A1O1Ixp33_ASAP7_75t_SL g2810 ( 
.A1(n_2742),
.A2(n_2530),
.B(n_2325),
.C(n_2361),
.Y(n_2810)
);

OAI21x1_ASAP7_75t_L g2811 ( 
.A1(n_2533),
.A2(n_2302),
.B(n_2300),
.Y(n_2811)
);

O2A1O1Ixp5_ASAP7_75t_L g2812 ( 
.A1(n_2720),
.A2(n_2403),
.B(n_2518),
.C(n_2516),
.Y(n_2812)
);

AO21x2_ASAP7_75t_L g2813 ( 
.A1(n_2674),
.A2(n_2400),
.B(n_2399),
.Y(n_2813)
);

OAI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2648),
.A2(n_2480),
.B(n_2500),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2747),
.A2(n_2487),
.B1(n_2359),
.B2(n_2375),
.Y(n_2815)
);

AOI21x1_ASAP7_75t_L g2816 ( 
.A1(n_2787),
.A2(n_2498),
.B(n_2494),
.Y(n_2816)
);

OAI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2779),
.A2(n_2359),
.B1(n_2375),
.B2(n_2416),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2619),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2603),
.B(n_2468),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2689),
.B(n_2341),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2548),
.Y(n_2821)
);

O2A1O1Ixp33_ASAP7_75t_L g2822 ( 
.A1(n_2720),
.A2(n_2513),
.B(n_2305),
.C(n_2403),
.Y(n_2822)
);

BUFx3_ASAP7_75t_L g2823 ( 
.A(n_2593),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2589),
.B(n_2535),
.Y(n_2824)
);

OAI21x1_ASAP7_75t_L g2825 ( 
.A1(n_2533),
.A2(n_2324),
.B(n_2315),
.Y(n_2825)
);

OR2x6_ASAP7_75t_L g2826 ( 
.A(n_2762),
.B(n_2360),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2719),
.B(n_2471),
.Y(n_2827)
);

OR2x6_ASAP7_75t_L g2828 ( 
.A(n_2762),
.B(n_2404),
.Y(n_2828)
);

A2O1A1Ixp33_ASAP7_75t_L g2829 ( 
.A1(n_2648),
.A2(n_2426),
.B(n_2378),
.C(n_2514),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2558),
.A2(n_2439),
.B(n_2297),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2574),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2583),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2585),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2558),
.A2(n_2642),
.B(n_2708),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2654),
.B(n_2399),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2551),
.Y(n_2836)
);

NOR2x1_ASAP7_75t_L g2837 ( 
.A(n_2552),
.B(n_2333),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2562),
.Y(n_2838)
);

BUFx2_ASAP7_75t_L g2839 ( 
.A(n_2561),
.Y(n_2839)
);

AOI221x1_ASAP7_75t_L g2840 ( 
.A1(n_2556),
.A2(n_2527),
.B1(n_2378),
.B2(n_2400),
.C(n_2337),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_2716),
.A2(n_2514),
.B1(n_2377),
.B2(n_542),
.Y(n_2841)
);

OA21x2_ASAP7_75t_L g2842 ( 
.A1(n_2667),
.A2(n_2458),
.B(n_2450),
.Y(n_2842)
);

BUFx6f_ASAP7_75t_L g2843 ( 
.A(n_2711),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2590),
.Y(n_2844)
);

OR2x6_ASAP7_75t_L g2845 ( 
.A(n_2762),
.B(n_2404),
.Y(n_2845)
);

OAI21x1_ASAP7_75t_L g2846 ( 
.A1(n_2631),
.A2(n_2357),
.B(n_2391),
.Y(n_2846)
);

OR2x6_ASAP7_75t_L g2847 ( 
.A(n_2712),
.B(n_2370),
.Y(n_2847)
);

NOR2x1_ASAP7_75t_SL g2848 ( 
.A(n_2665),
.B(n_2482),
.Y(n_2848)
);

OAI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2786),
.A2(n_2488),
.B(n_2461),
.Y(n_2849)
);

OA21x2_ASAP7_75t_L g2850 ( 
.A1(n_2623),
.A2(n_2460),
.B(n_2447),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_2553),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2568),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2699),
.A2(n_2507),
.B1(n_2445),
.B2(n_2466),
.Y(n_2853)
);

OR2x6_ASAP7_75t_L g2854 ( 
.A(n_2668),
.B(n_2356),
.Y(n_2854)
);

OAI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2786),
.A2(n_2465),
.B(n_2463),
.Y(n_2855)
);

BUFx4f_ASAP7_75t_SL g2856 ( 
.A(n_2633),
.Y(n_2856)
);

BUFx6f_ASAP7_75t_L g2857 ( 
.A(n_2538),
.Y(n_2857)
);

OAI21x1_ASAP7_75t_L g2858 ( 
.A1(n_2640),
.A2(n_2521),
.B(n_2449),
.Y(n_2858)
);

AOI221xp5_ASAP7_75t_L g2859 ( 
.A1(n_2703),
.A2(n_625),
.B1(n_639),
.B2(n_623),
.C(n_620),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2591),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2575),
.Y(n_2861)
);

AOI22xp33_ASAP7_75t_SL g2862 ( 
.A1(n_2708),
.A2(n_542),
.B1(n_2474),
.B2(n_2473),
.Y(n_2862)
);

OAI21x1_ASAP7_75t_L g2863 ( 
.A1(n_2536),
.A2(n_2443),
.B(n_2437),
.Y(n_2863)
);

INVxp67_ASAP7_75t_L g2864 ( 
.A(n_2748),
.Y(n_2864)
);

OAI21x1_ASAP7_75t_SL g2865 ( 
.A1(n_2669),
.A2(n_2478),
.B(n_2441),
.Y(n_2865)
);

AOI21xp33_ASAP7_75t_SL g2866 ( 
.A1(n_2542),
.A2(n_13),
.B(n_15),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2535),
.B(n_2529),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2604),
.Y(n_2868)
);

OAI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2536),
.A2(n_2412),
.B(n_2395),
.Y(n_2869)
);

OAI21x1_ASAP7_75t_L g2870 ( 
.A1(n_2679),
.A2(n_2415),
.B(n_2413),
.Y(n_2870)
);

OAI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2787),
.A2(n_2475),
.B(n_2505),
.Y(n_2871)
);

OAI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2701),
.A2(n_2704),
.B1(n_2581),
.B2(n_2702),
.Y(n_2872)
);

CKINVDCx5p33_ASAP7_75t_R g2873 ( 
.A(n_2607),
.Y(n_2873)
);

OAI21x1_ASAP7_75t_L g2874 ( 
.A1(n_2668),
.A2(n_2508),
.B(n_2529),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2586),
.Y(n_2875)
);

OAI21x1_ASAP7_75t_L g2876 ( 
.A1(n_2745),
.A2(n_2529),
.B(n_2519),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2702),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2877)
);

AO21x2_ASAP7_75t_L g2878 ( 
.A1(n_2686),
.A2(n_2519),
.B(n_1271),
.Y(n_2878)
);

INVx2_ASAP7_75t_SL g2879 ( 
.A(n_2553),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2600),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2783),
.A2(n_542),
.B1(n_1056),
.B2(n_1051),
.Y(n_2881)
);

OA21x2_ASAP7_75t_L g2882 ( 
.A1(n_2637),
.A2(n_649),
.B(n_645),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2602),
.Y(n_2883)
);

NAND2x1p5_ASAP7_75t_L g2884 ( 
.A(n_2657),
.B(n_1056),
.Y(n_2884)
);

INVx2_ASAP7_75t_SL g2885 ( 
.A(n_2567),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2592),
.A2(n_21),
.B1(n_16),
.B2(n_18),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2608),
.Y(n_2887)
);

OAI211xp5_ASAP7_75t_L g2888 ( 
.A1(n_2663),
.A2(n_24),
.B(n_21),
.C(n_23),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2577),
.A2(n_542),
.B1(n_1057),
.B2(n_1056),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2577),
.A2(n_542),
.B1(n_1057),
.B2(n_1056),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2609),
.Y(n_2891)
);

NAND2x1p5_ASAP7_75t_L g2892 ( 
.A(n_2657),
.B(n_1056),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2725),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_SL g2894 ( 
.A(n_2781),
.B(n_542),
.Y(n_2894)
);

BUFx12f_ASAP7_75t_L g2895 ( 
.A(n_2540),
.Y(n_2895)
);

NOR3xp33_ASAP7_75t_L g2896 ( 
.A(n_2557),
.B(n_2718),
.C(n_2703),
.Y(n_2896)
);

OAI21x1_ASAP7_75t_L g2897 ( 
.A1(n_2759),
.A2(n_2519),
.B(n_1057),
.Y(n_2897)
);

A2O1A1Ixp33_ASAP7_75t_L g2898 ( 
.A1(n_2660),
.A2(n_652),
.B(n_672),
.C(n_650),
.Y(n_2898)
);

NOR2xp67_ASAP7_75t_L g2899 ( 
.A(n_2552),
.B(n_23),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2549),
.Y(n_2900)
);

NAND3xp33_ASAP7_75t_SL g2901 ( 
.A(n_2592),
.B(n_688),
.C(n_677),
.Y(n_2901)
);

NAND2x1p5_ASAP7_75t_L g2902 ( 
.A(n_2657),
.B(n_1057),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_2659),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2718),
.A2(n_542),
.B1(n_1057),
.B2(n_1040),
.Y(n_2904)
);

A2O1A1Ixp33_ASAP7_75t_L g2905 ( 
.A1(n_2660),
.A2(n_707),
.B(n_729),
.C(n_692),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2726),
.Y(n_2906)
);

OAI21x1_ASAP7_75t_L g2907 ( 
.A1(n_2729),
.A2(n_1057),
.B(n_542),
.Y(n_2907)
);

NAND2x1_ASAP7_75t_L g2908 ( 
.A(n_2740),
.B(n_969),
.Y(n_2908)
);

AO21x2_ASAP7_75t_L g2909 ( 
.A1(n_2691),
.A2(n_1040),
.B(n_1026),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2651),
.Y(n_2910)
);

INVxp67_ASAP7_75t_L g2911 ( 
.A(n_2760),
.Y(n_2911)
);

BUFx3_ASAP7_75t_L g2912 ( 
.A(n_2625),
.Y(n_2912)
);

AO31x2_ASAP7_75t_L g2913 ( 
.A1(n_2737),
.A2(n_1040),
.A3(n_1026),
.B(n_27),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2664),
.Y(n_2914)
);

OAI21x1_ASAP7_75t_L g2915 ( 
.A1(n_2729),
.A2(n_1040),
.B(n_1026),
.Y(n_2915)
);

AOI21x1_ASAP7_75t_L g2916 ( 
.A1(n_2782),
.A2(n_738),
.B(n_733),
.Y(n_2916)
);

OAI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2687),
.A2(n_751),
.B(n_742),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2653),
.B(n_25),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2554),
.B(n_25),
.Y(n_2919)
);

AOI22xp33_ASAP7_75t_L g2920 ( 
.A1(n_2730),
.A2(n_1040),
.B1(n_1026),
.B2(n_758),
.Y(n_2920)
);

OA21x2_ASAP7_75t_L g2921 ( 
.A1(n_2732),
.A2(n_769),
.B(n_754),
.Y(n_2921)
);

AOI22xp33_ASAP7_75t_SL g2922 ( 
.A1(n_2715),
.A2(n_789),
.B1(n_770),
.B2(n_28),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2588),
.Y(n_2923)
);

OAI21x1_ASAP7_75t_L g2924 ( 
.A1(n_2756),
.A2(n_1026),
.B(n_354),
.Y(n_2924)
);

OR2x2_ASAP7_75t_L g2925 ( 
.A(n_2653),
.B(n_26),
.Y(n_2925)
);

OAI21x1_ASAP7_75t_L g2926 ( 
.A1(n_2756),
.A2(n_355),
.B(n_352),
.Y(n_2926)
);

INVx5_ASAP7_75t_L g2927 ( 
.A(n_2566),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2588),
.Y(n_2928)
);

OA21x2_ASAP7_75t_L g2929 ( 
.A1(n_2735),
.A2(n_2688),
.B(n_2626),
.Y(n_2929)
);

BUFx12f_ASAP7_75t_L g2930 ( 
.A(n_2644),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2683),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2717),
.Y(n_2932)
);

NAND2x1p5_ASAP7_75t_L g2933 ( 
.A(n_2657),
.B(n_969),
.Y(n_2933)
);

OA21x2_ASAP7_75t_L g2934 ( 
.A1(n_2688),
.A2(n_26),
.B(n_27),
.Y(n_2934)
);

NOR2xp67_ASAP7_75t_SL g2935 ( 
.A(n_2680),
.B(n_969),
.Y(n_2935)
);

BUFx2_ASAP7_75t_R g2936 ( 
.A(n_2632),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2744),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_L g2938 ( 
.A(n_2538),
.Y(n_2938)
);

INVx3_ASAP7_75t_L g2939 ( 
.A(n_2700),
.Y(n_2939)
);

AND2x4_ASAP7_75t_L g2940 ( 
.A(n_2554),
.B(n_28),
.Y(n_2940)
);

BUFx2_ASAP7_75t_L g2941 ( 
.A(n_2579),
.Y(n_2941)
);

O2A1O1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2770),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_2942)
);

OR2x2_ASAP7_75t_L g2943 ( 
.A(n_2560),
.B(n_30),
.Y(n_2943)
);

OAI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2771),
.A2(n_31),
.B(n_32),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2630),
.Y(n_2945)
);

BUFx3_ASAP7_75t_L g2946 ( 
.A(n_2618),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2697),
.A2(n_974),
.B1(n_976),
.B2(n_969),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2724),
.Y(n_2948)
);

CKINVDCx5p33_ASAP7_75t_R g2949 ( 
.A(n_2656),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2731),
.Y(n_2950)
);

AO21x2_ASAP7_75t_L g2951 ( 
.A1(n_2685),
.A2(n_974),
.B(n_969),
.Y(n_2951)
);

AOI22xp33_ASAP7_75t_SL g2952 ( 
.A1(n_2665),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2559),
.B(n_2560),
.Y(n_2953)
);

AO31x2_ASAP7_75t_L g2954 ( 
.A1(n_2670),
.A2(n_35),
.A3(n_33),
.B(n_34),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2676),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_2955)
);

BUFx6f_ASAP7_75t_L g2956 ( 
.A(n_2538),
.Y(n_2956)
);

OR2x2_ASAP7_75t_L g2957 ( 
.A(n_2559),
.B(n_37),
.Y(n_2957)
);

AO21x2_ASAP7_75t_L g2958 ( 
.A1(n_2790),
.A2(n_974),
.B(n_969),
.Y(n_2958)
);

AO31x2_ASAP7_75t_L g2959 ( 
.A1(n_2767),
.A2(n_40),
.A3(n_38),
.B(n_39),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2537),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2722),
.Y(n_2961)
);

OAI21x1_ASAP7_75t_L g2962 ( 
.A1(n_2788),
.A2(n_358),
.B(n_357),
.Y(n_2962)
);

AOI21x1_ASAP7_75t_L g2963 ( 
.A1(n_2778),
.A2(n_41),
.B(n_42),
.Y(n_2963)
);

AOI221xp5_ASAP7_75t_L g2964 ( 
.A1(n_2770),
.A2(n_49),
.B1(n_44),
.B2(n_45),
.C(n_50),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2709),
.Y(n_2965)
);

AOI22xp5_ASAP7_75t_L g2966 ( 
.A1(n_2723),
.A2(n_987),
.B1(n_976),
.B2(n_984),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2534),
.A2(n_50),
.B1(n_44),
.B2(n_45),
.Y(n_2967)
);

INVx3_ASAP7_75t_L g2968 ( 
.A(n_2700),
.Y(n_2968)
);

CKINVDCx5p33_ASAP7_75t_R g2969 ( 
.A(n_2624),
.Y(n_2969)
);

NOR2xp67_ASAP7_75t_L g2970 ( 
.A(n_2594),
.B(n_53),
.Y(n_2970)
);

OR2x6_ASAP7_75t_L g2971 ( 
.A(n_2595),
.B(n_974),
.Y(n_2971)
);

CKINVDCx5p33_ASAP7_75t_R g2972 ( 
.A(n_2572),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2649),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2710),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2721),
.Y(n_2975)
);

OA21x2_ASAP7_75t_L g2976 ( 
.A1(n_2626),
.A2(n_53),
.B(n_55),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2649),
.Y(n_2977)
);

AO21x2_ASAP7_75t_L g2978 ( 
.A1(n_2790),
.A2(n_976),
.B(n_974),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_SL g2979 ( 
.A1(n_2727),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2979)
);

OAI21x1_ASAP7_75t_L g2980 ( 
.A1(n_2788),
.A2(n_360),
.B(n_359),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2784),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2661),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2661),
.Y(n_2983)
);

HB1xp67_ASAP7_75t_L g2984 ( 
.A(n_2746),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2645),
.B(n_56),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_L g2986 ( 
.A1(n_2746),
.A2(n_363),
.B(n_362),
.Y(n_2986)
);

CKINVDCx11_ASAP7_75t_R g2987 ( 
.A(n_2728),
.Y(n_2987)
);

INVx1_ASAP7_75t_SL g2988 ( 
.A(n_2545),
.Y(n_2988)
);

OA21x2_ASAP7_75t_L g2989 ( 
.A1(n_2595),
.A2(n_58),
.B(n_59),
.Y(n_2989)
);

CKINVDCx11_ASAP7_75t_R g2990 ( 
.A(n_2728),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2707),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2681),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2621),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2681),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2627),
.Y(n_2995)
);

AND2x6_ASAP7_75t_L g2996 ( 
.A(n_2598),
.B(n_974),
.Y(n_2996)
);

BUFx2_ASAP7_75t_L g2997 ( 
.A(n_2546),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2587),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2998)
);

OAI21x1_ASAP7_75t_L g2999 ( 
.A1(n_2634),
.A2(n_369),
.B(n_366),
.Y(n_2999)
);

OAI21x1_ASAP7_75t_L g3000 ( 
.A1(n_2634),
.A2(n_372),
.B(n_371),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2627),
.Y(n_3001)
);

BUFx3_ASAP7_75t_L g3002 ( 
.A(n_2620),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2652),
.B(n_67),
.Y(n_3003)
);

OAI21x1_ASAP7_75t_L g3004 ( 
.A1(n_2740),
.A2(n_376),
.B(n_374),
.Y(n_3004)
);

INVx6_ASAP7_75t_L g3005 ( 
.A(n_2539),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2743),
.Y(n_3006)
);

BUFx6f_ASAP7_75t_L g3007 ( 
.A(n_2539),
.Y(n_3007)
);

OA21x2_ASAP7_75t_L g3008 ( 
.A1(n_2750),
.A2(n_2754),
.B(n_2752),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2587),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_2622),
.Y(n_3010)
);

NOR2xp67_ASAP7_75t_L g3011 ( 
.A(n_2594),
.B(n_70),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2953),
.B(n_2616),
.Y(n_3012)
);

INVx6_ASAP7_75t_L g3013 ( 
.A(n_2930),
.Y(n_3013)
);

CKINVDCx6p67_ASAP7_75t_R g3014 ( 
.A(n_2805),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2923),
.B(n_2766),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2910),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2824),
.B(n_2546),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_2953),
.B(n_2616),
.Y(n_3018)
);

INVx4_ASAP7_75t_L g3019 ( 
.A(n_2806),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2896),
.A2(n_2599),
.B1(n_2598),
.B2(n_2584),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2896),
.A2(n_2872),
.B1(n_2803),
.B2(n_2815),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2798),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2804),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2839),
.B(n_2610),
.Y(n_3024)
);

OAI221xp5_ASAP7_75t_L g3025 ( 
.A1(n_2979),
.A2(n_2785),
.B1(n_2628),
.B2(n_2684),
.C(n_2597),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2991),
.A2(n_2772),
.B1(n_2541),
.B2(n_2565),
.Y(n_3026)
);

INVxp33_ASAP7_75t_SL g3027 ( 
.A(n_2903),
.Y(n_3027)
);

OAI22xp5_ASAP7_75t_L g3028 ( 
.A1(n_2991),
.A2(n_2541),
.B1(n_2565),
.B2(n_2739),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2928),
.B(n_2766),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2836),
.Y(n_3030)
);

AO21x2_ASAP7_75t_L g3031 ( 
.A1(n_2894),
.A2(n_2741),
.B(n_2774),
.Y(n_3031)
);

INVx2_ASAP7_75t_SL g3032 ( 
.A(n_2823),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2955),
.A2(n_2695),
.B1(n_2680),
.B2(n_2678),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2838),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2875),
.Y(n_3035)
);

OAI222xp33_ASAP7_75t_L g3036 ( 
.A1(n_2872),
.A2(n_2713),
.B1(n_2789),
.B2(n_2736),
.C1(n_2734),
.C2(n_2693),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_2941),
.B(n_2613),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2852),
.Y(n_3038)
);

INVx3_ASAP7_75t_L g3039 ( 
.A(n_2946),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2973),
.B(n_2977),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2887),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2799),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2818),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_2873),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2815),
.A2(n_2671),
.B1(n_2677),
.B2(n_2675),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2895),
.Y(n_3046)
);

NAND3xp33_ASAP7_75t_L g3047 ( 
.A(n_2952),
.B(n_2753),
.C(n_2771),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2965),
.Y(n_3048)
);

AOI21xp33_ASAP7_75t_L g3049 ( 
.A1(n_2877),
.A2(n_2713),
.B(n_2763),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2834),
.A2(n_2578),
.B(n_2765),
.Y(n_3050)
);

OAI21x1_ASAP7_75t_L g3051 ( 
.A1(n_2834),
.A2(n_2825),
.B(n_2811),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2830),
.A2(n_2578),
.B(n_2765),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2901),
.A2(n_2671),
.B1(n_2677),
.B2(n_2675),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2791),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_2997),
.B(n_2616),
.Y(n_3055)
);

AOI221xp5_ASAP7_75t_L g3056 ( 
.A1(n_2886),
.A2(n_2682),
.B1(n_2773),
.B2(n_2757),
.C(n_2650),
.Y(n_3056)
);

OAI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_2955),
.A2(n_2680),
.B1(n_2765),
.B2(n_2755),
.Y(n_3057)
);

OAI22xp33_ASAP7_75t_SL g3058 ( 
.A1(n_2918),
.A2(n_2544),
.B1(n_2569),
.B2(n_2789),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2982),
.B(n_2983),
.Y(n_3059)
);

AO32x2_ASAP7_75t_L g3060 ( 
.A1(n_2817),
.A2(n_2776),
.A3(n_2672),
.B1(n_2658),
.B2(n_2766),
.Y(n_3060)
);

AOI22xp33_ASAP7_75t_L g3061 ( 
.A1(n_2901),
.A2(n_2671),
.B1(n_2677),
.B2(n_2675),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_SL g3062 ( 
.A1(n_2882),
.A2(n_2766),
.B1(n_2680),
.B2(n_2655),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2974),
.Y(n_3063)
);

NAND2x1_ASAP7_75t_L g3064 ( 
.A(n_2939),
.B(n_2672),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2975),
.Y(n_3065)
);

INVx3_ASAP7_75t_L g3066 ( 
.A(n_2939),
.Y(n_3066)
);

AND2x4_ASAP7_75t_L g3067 ( 
.A(n_2968),
.B(n_2900),
.Y(n_3067)
);

OAI22xp33_ASAP7_75t_SL g3068 ( 
.A1(n_2925),
.A2(n_2635),
.B1(n_2571),
.B2(n_2601),
.Y(n_3068)
);

OR2x2_ASAP7_75t_L g3069 ( 
.A(n_2992),
.B(n_2613),
.Y(n_3069)
);

AOI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2830),
.A2(n_2829),
.B(n_2822),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2861),
.Y(n_3071)
);

HB1xp67_ASAP7_75t_L g3072 ( 
.A(n_2864),
.Y(n_3072)
);

AND2x4_ASAP7_75t_L g3073 ( 
.A(n_2968),
.B(n_2690),
.Y(n_3073)
);

OAI221xp5_ASAP7_75t_L g3074 ( 
.A1(n_2979),
.A2(n_2751),
.B1(n_2673),
.B2(n_2773),
.C(n_2647),
.Y(n_3074)
);

O2A1O1Ixp33_ASAP7_75t_SL g3075 ( 
.A1(n_2998),
.A2(n_2605),
.B(n_74),
.C(n_71),
.Y(n_3075)
);

OAI21x1_ASAP7_75t_L g3076 ( 
.A1(n_2846),
.A2(n_2571),
.B(n_2555),
.Y(n_3076)
);

OAI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_2817),
.A2(n_2705),
.B1(n_2698),
.B2(n_2733),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2994),
.B(n_2995),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2880),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_2921),
.A2(n_2698),
.B1(n_2705),
.B2(n_2766),
.Y(n_3080)
);

AND2x2_ASAP7_75t_SL g3081 ( 
.A(n_2800),
.B(n_2919),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2883),
.Y(n_3082)
);

AOI222xp33_ASAP7_75t_L g3083 ( 
.A1(n_2964),
.A2(n_2705),
.B1(n_2698),
.B2(n_2761),
.C1(n_2777),
.C2(n_2706),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_2921),
.A2(n_2952),
.B1(n_2882),
.B2(n_2886),
.Y(n_3084)
);

CKINVDCx5p33_ASAP7_75t_R g3085 ( 
.A(n_2969),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_L g3086 ( 
.A1(n_2922),
.A2(n_2617),
.B1(n_2612),
.B2(n_2776),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2891),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2922),
.A2(n_2612),
.B1(n_2563),
.B2(n_2576),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_SL g3089 ( 
.A(n_2800),
.B(n_2655),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_2988),
.B(n_2714),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2914),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_2964),
.A2(n_2890),
.B1(n_2889),
.B2(n_2881),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2889),
.A2(n_2706),
.B1(n_2733),
.B2(n_2601),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_SL g3094 ( 
.A1(n_2934),
.A2(n_2655),
.B1(n_2733),
.B2(n_2714),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2948),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3001),
.B(n_2690),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2961),
.B(n_2690),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_SL g3098 ( 
.A1(n_2934),
.A2(n_2655),
.B1(n_2714),
.B2(n_2780),
.Y(n_3098)
);

AND2x4_ASAP7_75t_L g3099 ( 
.A(n_2867),
.B(n_2690),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_2927),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2950),
.Y(n_3101)
);

INVx4_ASAP7_75t_L g3102 ( 
.A(n_2843),
.Y(n_3102)
);

NAND2xp33_ASAP7_75t_L g3103 ( 
.A(n_2949),
.B(n_2655),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2864),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2821),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2927),
.Y(n_3106)
);

NAND2x1p5_ASAP7_75t_L g3107 ( 
.A(n_2927),
.B(n_2566),
.Y(n_3107)
);

AND2x4_ASAP7_75t_L g3108 ( 
.A(n_2851),
.B(n_2615),
.Y(n_3108)
);

OR2x6_ASAP7_75t_L g3109 ( 
.A(n_2800),
.B(n_2828),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3006),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_2890),
.A2(n_2638),
.B1(n_2641),
.B2(n_2555),
.Y(n_3111)
);

INVxp67_ASAP7_75t_L g3112 ( 
.A(n_2936),
.Y(n_3112)
);

AOI22xp33_ASAP7_75t_L g3113 ( 
.A1(n_2881),
.A2(n_2641),
.B1(n_2646),
.B2(n_2638),
.Y(n_3113)
);

BUFx12f_ASAP7_75t_L g3114 ( 
.A(n_2919),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_2912),
.Y(n_3115)
);

NAND2xp33_ASAP7_75t_SL g3116 ( 
.A(n_3010),
.B(n_2539),
.Y(n_3116)
);

OR2x2_ASAP7_75t_L g3117 ( 
.A(n_2827),
.B(n_2666),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2831),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2829),
.A2(n_2580),
.B(n_2566),
.Y(n_3119)
);

BUFx2_ASAP7_75t_L g3120 ( 
.A(n_3002),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3008),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2960),
.A2(n_2563),
.B1(n_2576),
.B2(n_2566),
.Y(n_3122)
);

INVx4_ASAP7_75t_L g3123 ( 
.A(n_2843),
.Y(n_3123)
);

HB1xp67_ASAP7_75t_L g3124 ( 
.A(n_2794),
.Y(n_3124)
);

OAI21xp33_ASAP7_75t_L g3125 ( 
.A1(n_2877),
.A2(n_2764),
.B(n_2666),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2832),
.Y(n_3126)
);

AND2x4_ASAP7_75t_L g3127 ( 
.A(n_2879),
.B(n_2615),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_2894),
.A2(n_2646),
.B1(n_2738),
.B2(n_2643),
.Y(n_3128)
);

HB1xp67_ASAP7_75t_L g3129 ( 
.A(n_2794),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3008),
.Y(n_3130)
);

NAND2xp33_ASAP7_75t_L g3131 ( 
.A(n_2800),
.B(n_2714),
.Y(n_3131)
);

NOR2xp33_ASAP7_75t_R g3132 ( 
.A(n_2972),
.B(n_2683),
.Y(n_3132)
);

OAI211xp5_ASAP7_75t_SL g3133 ( 
.A1(n_2998),
.A2(n_3009),
.B(n_2917),
.C(n_2859),
.Y(n_3133)
);

BUFx12f_ASAP7_75t_L g3134 ( 
.A(n_2940),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_2917),
.A2(n_2738),
.B1(n_2643),
.B2(n_2636),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_2827),
.B(n_2666),
.Y(n_3136)
);

OAI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2960),
.A2(n_2563),
.B1(n_2576),
.B2(n_2580),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2833),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2932),
.Y(n_3139)
);

AO21x2_ASAP7_75t_L g3140 ( 
.A1(n_2819),
.A2(n_2764),
.B(n_2636),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2819),
.B(n_2714),
.Y(n_3141)
);

NAND2xp33_ASAP7_75t_R g3142 ( 
.A(n_2940),
.B(n_2957),
.Y(n_3142)
);

OAI22xp5_ASAP7_75t_SL g3143 ( 
.A1(n_2856),
.A2(n_2580),
.B1(n_2564),
.B2(n_2570),
.Y(n_3143)
);

AOI22xp33_ASAP7_75t_L g3144 ( 
.A1(n_2814),
.A2(n_2780),
.B1(n_2564),
.B2(n_2570),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2856),
.B(n_2547),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_3009),
.A2(n_2580),
.B1(n_2780),
.B2(n_2564),
.Y(n_3146)
);

OAI221xp5_ASAP7_75t_L g3147 ( 
.A1(n_2888),
.A2(n_2573),
.B1(n_2582),
.B2(n_2570),
.C(n_2547),
.Y(n_3147)
);

AOI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2888),
.A2(n_2696),
.B1(n_2692),
.B2(n_2573),
.Y(n_3148)
);

AOI22xp33_ASAP7_75t_L g3149 ( 
.A1(n_2814),
.A2(n_2573),
.B1(n_2582),
.B2(n_2547),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2844),
.Y(n_3150)
);

BUFx6f_ASAP7_75t_L g3151 ( 
.A(n_2843),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2860),
.Y(n_3152)
);

O2A1O1Ixp33_ASAP7_75t_L g3153 ( 
.A1(n_2866),
.A2(n_2696),
.B(n_2692),
.C(n_75),
.Y(n_3153)
);

AOI22xp33_ASAP7_75t_SL g3154 ( 
.A1(n_2976),
.A2(n_2596),
.B1(n_2614),
.B2(n_2582),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2981),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_2976),
.A2(n_2614),
.B1(n_2596),
.B2(n_984),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2893),
.Y(n_3157)
);

NAND3xp33_ASAP7_75t_SL g3158 ( 
.A(n_2802),
.B(n_72),
.C(n_74),
.Y(n_3158)
);

BUFx12f_ASAP7_75t_L g3159 ( 
.A(n_2987),
.Y(n_3159)
);

INVx3_ASAP7_75t_L g3160 ( 
.A(n_2927),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2808),
.A2(n_2614),
.B1(n_2596),
.B2(n_984),
.Y(n_3161)
);

BUFx3_ASAP7_75t_L g3162 ( 
.A(n_2885),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2808),
.A2(n_984),
.B1(n_986),
.B2(n_976),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2906),
.Y(n_3164)
);

AOI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_2859),
.A2(n_984),
.B1(n_986),
.B2(n_976),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2936),
.B(n_72),
.Y(n_3166)
);

AOI22xp33_ASAP7_75t_L g3167 ( 
.A1(n_2967),
.A2(n_984),
.B1(n_986),
.B2(n_976),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2990),
.Y(n_3168)
);

HB1xp67_ASAP7_75t_L g3169 ( 
.A(n_2911),
.Y(n_3169)
);

BUFx2_ASAP7_75t_L g3170 ( 
.A(n_2931),
.Y(n_3170)
);

CKINVDCx11_ASAP7_75t_R g3171 ( 
.A(n_2843),
.Y(n_3171)
);

BUFx3_ASAP7_75t_L g3172 ( 
.A(n_3005),
.Y(n_3172)
);

OAI21x1_ASAP7_75t_L g3173 ( 
.A1(n_2792),
.A2(n_76),
.B(n_77),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_2931),
.B(n_2911),
.Y(n_3174)
);

AND2x4_ASAP7_75t_L g3175 ( 
.A(n_2847),
.B(n_78),
.Y(n_3175)
);

INVx6_ASAP7_75t_L g3176 ( 
.A(n_3005),
.Y(n_3176)
);

AO21x2_ASAP7_75t_L g3177 ( 
.A1(n_2813),
.A2(n_78),
.B(n_79),
.Y(n_3177)
);

INVx4_ASAP7_75t_L g3178 ( 
.A(n_2931),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2868),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2945),
.Y(n_3180)
);

OR2x2_ASAP7_75t_L g3181 ( 
.A(n_2820),
.B(n_80),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_SL g3182 ( 
.A(n_2865),
.B(n_986),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_2943),
.B(n_80),
.Y(n_3183)
);

HB1xp67_ASAP7_75t_L g3184 ( 
.A(n_2820),
.Y(n_3184)
);

CKINVDCx5p33_ASAP7_75t_R g3185 ( 
.A(n_3005),
.Y(n_3185)
);

A2O1A1Ixp33_ASAP7_75t_L g3186 ( 
.A1(n_2809),
.A2(n_2942),
.B(n_2822),
.C(n_2905),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_2967),
.A2(n_987),
.B1(n_986),
.B2(n_83),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_SL g3188 ( 
.A(n_2931),
.B(n_986),
.Y(n_3188)
);

OR2x6_ASAP7_75t_L g3189 ( 
.A(n_2828),
.B(n_987),
.Y(n_3189)
);

A2O1A1Ixp33_ASAP7_75t_L g3190 ( 
.A1(n_2809),
.A2(n_84),
.B(n_81),
.C(n_82),
.Y(n_3190)
);

AND2x4_ASAP7_75t_L g3191 ( 
.A(n_2847),
.B(n_82),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2796),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2796),
.Y(n_3193)
);

BUFx6f_ASAP7_75t_L g3194 ( 
.A(n_2857),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2937),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2929),
.B(n_86),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2989),
.A2(n_987),
.B1(n_88),
.B2(n_86),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2835),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2857),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2835),
.Y(n_3200)
);

BUFx8_ASAP7_75t_L g3201 ( 
.A(n_2857),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_2938),
.Y(n_3202)
);

O2A1O1Ixp33_ASAP7_75t_L g3203 ( 
.A1(n_2942),
.A2(n_90),
.B(n_87),
.C(n_89),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2929),
.Y(n_3204)
);

INVx4_ASAP7_75t_SL g3205 ( 
.A(n_2996),
.Y(n_3205)
);

HB1xp67_ASAP7_75t_L g3206 ( 
.A(n_2984),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2984),
.B(n_87),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_3192),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3121),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3130),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_3204),
.Y(n_3211)
);

AO21x2_ASAP7_75t_L g3212 ( 
.A1(n_3070),
.A2(n_2848),
.B(n_2813),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3024),
.B(n_2854),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3124),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3129),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_3193),
.Y(n_3216)
);

INVx3_ASAP7_75t_L g3217 ( 
.A(n_3178),
.Y(n_3217)
);

AOI21x1_ASAP7_75t_L g3218 ( 
.A1(n_3196),
.A2(n_3207),
.B(n_3070),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3196),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3140),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_3178),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3040),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3040),
.Y(n_3223)
);

INVx4_ASAP7_75t_L g3224 ( 
.A(n_3159),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3140),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_3068),
.B(n_2938),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3059),
.Y(n_3227)
);

BUFx2_ASAP7_75t_SL g3228 ( 
.A(n_3019),
.Y(n_3228)
);

AO21x2_ASAP7_75t_L g3229 ( 
.A1(n_3177),
.A2(n_2876),
.B(n_2909),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3015),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3059),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_3177),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_3189),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3078),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3078),
.Y(n_3235)
);

OAI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_3021),
.A2(n_2812),
.B(n_2970),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3198),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3200),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3037),
.B(n_2854),
.Y(n_3239)
);

HB1xp67_ASAP7_75t_L g3240 ( 
.A(n_3169),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3027),
.B(n_2916),
.Y(n_3241)
);

HB1xp67_ASAP7_75t_L g3242 ( 
.A(n_3072),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3104),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3184),
.B(n_2854),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_3039),
.B(n_2847),
.Y(n_3245)
);

AO21x2_ASAP7_75t_L g3246 ( 
.A1(n_3186),
.A2(n_2909),
.B(n_2963),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3022),
.Y(n_3247)
);

INVx1_ASAP7_75t_SL g3248 ( 
.A(n_3171),
.Y(n_3248)
);

HB1xp67_ASAP7_75t_L g3249 ( 
.A(n_3206),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3023),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3015),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3030),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3034),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_3084),
.A2(n_3133),
.B1(n_3025),
.B2(n_3092),
.Y(n_3254)
);

INVx3_ASAP7_75t_L g3255 ( 
.A(n_3100),
.Y(n_3255)
);

OAI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3190),
.A2(n_2812),
.B(n_3011),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_3168),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3038),
.Y(n_3258)
);

OR2x6_ASAP7_75t_L g3259 ( 
.A(n_3119),
.B(n_3109),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3071),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3029),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3079),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3039),
.B(n_2826),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3029),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3031),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3082),
.Y(n_3266)
);

AND2x4_ASAP7_75t_L g3267 ( 
.A(n_3175),
.B(n_2826),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3087),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_3100),
.Y(n_3269)
);

BUFx3_ASAP7_75t_L g3270 ( 
.A(n_3014),
.Y(n_3270)
);

NAND2x1p5_ASAP7_75t_L g3271 ( 
.A(n_3175),
.B(n_2989),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3031),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_3180),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3174),
.B(n_3067),
.Y(n_3274)
);

OA21x2_ASAP7_75t_L g3275 ( 
.A1(n_3051),
.A2(n_2801),
.B(n_2840),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3016),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_3106),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3091),
.Y(n_3278)
);

OAI21x1_ASAP7_75t_L g3279 ( 
.A1(n_3052),
.A2(n_2793),
.B(n_2797),
.Y(n_3279)
);

INVx2_ASAP7_75t_SL g3280 ( 
.A(n_3176),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3095),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_3067),
.B(n_2826),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3060),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3101),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_3060),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_3120),
.B(n_2971),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3110),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_L g3288 ( 
.A1(n_3025),
.A2(n_2853),
.B1(n_2993),
.B2(n_2841),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3048),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3063),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3017),
.B(n_2971),
.Y(n_3291)
);

OAI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3203),
.A2(n_2944),
.B(n_2899),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3141),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3207),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3065),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3141),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3035),
.Y(n_3297)
);

HB1xp67_ASAP7_75t_L g3298 ( 
.A(n_3181),
.Y(n_3298)
);

AO21x1_ASAP7_75t_SL g3299 ( 
.A1(n_3149),
.A2(n_3003),
.B(n_2985),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3041),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_3042),
.Y(n_3301)
);

BUFx4f_ASAP7_75t_L g3302 ( 
.A(n_3046),
.Y(n_3302)
);

INVxp67_ASAP7_75t_L g3303 ( 
.A(n_3142),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3060),
.B(n_2971),
.Y(n_3304)
);

BUFx2_ASAP7_75t_L g3305 ( 
.A(n_3132),
.Y(n_3305)
);

AO21x2_ASAP7_75t_L g3306 ( 
.A1(n_3049),
.A2(n_3003),
.B(n_2985),
.Y(n_3306)
);

AO21x2_ASAP7_75t_L g3307 ( 
.A1(n_3049),
.A2(n_2878),
.B(n_2951),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3162),
.B(n_2807),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3043),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3096),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3096),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3066),
.B(n_2807),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3117),
.Y(n_3313)
);

BUFx2_ASAP7_75t_L g3314 ( 
.A(n_3170),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3136),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3090),
.B(n_2954),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3105),
.Y(n_3317)
);

BUFx2_ASAP7_75t_L g3318 ( 
.A(n_3066),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3118),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3097),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3126),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3138),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3097),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3069),
.Y(n_3324)
);

NAND2x1p5_ASAP7_75t_L g3325 ( 
.A(n_3191),
.B(n_2935),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3199),
.B(n_2807),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_3099),
.B(n_3172),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3099),
.B(n_2807),
.Y(n_3328)
);

INVxp67_ASAP7_75t_SL g3329 ( 
.A(n_3058),
.Y(n_3329)
);

INVx4_ASAP7_75t_L g3330 ( 
.A(n_3013),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3139),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3032),
.B(n_2958),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3150),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3155),
.Y(n_3334)
);

NOR2xp67_ASAP7_75t_L g3335 ( 
.A(n_3052),
.B(n_2947),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3157),
.Y(n_3336)
);

AND2x2_ASAP7_75t_L g3337 ( 
.A(n_3073),
.B(n_2958),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3164),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_3106),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_3019),
.B(n_2938),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3152),
.Y(n_3341)
);

HB1xp67_ASAP7_75t_L g3342 ( 
.A(n_3076),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3073),
.B(n_2978),
.Y(n_3343)
);

AOI21x1_ASAP7_75t_L g3344 ( 
.A1(n_3191),
.A2(n_2908),
.B(n_2837),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3081),
.B(n_2978),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3012),
.B(n_3018),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3125),
.B(n_2954),
.Y(n_3347)
);

OR2x2_ASAP7_75t_L g3348 ( 
.A(n_3195),
.B(n_2954),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3179),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3064),
.Y(n_3350)
);

O2A1O1Ixp33_ASAP7_75t_SL g3351 ( 
.A1(n_3112),
.A2(n_2905),
.B(n_2898),
.C(n_2944),
.Y(n_3351)
);

HB1xp67_ASAP7_75t_L g3352 ( 
.A(n_3176),
.Y(n_3352)
);

OAI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3203),
.A2(n_3158),
.B(n_3153),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_L g3354 ( 
.A(n_3013),
.B(n_2956),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3205),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3205),
.Y(n_3356)
);

INVx2_ASAP7_75t_SL g3357 ( 
.A(n_3185),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3205),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3109),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3154),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3173),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3189),
.Y(n_3362)
);

OR2x2_ASAP7_75t_L g3363 ( 
.A(n_3028),
.B(n_2954),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3028),
.Y(n_3364)
);

INVx4_ASAP7_75t_L g3365 ( 
.A(n_3046),
.Y(n_3365)
);

NOR2xp67_ASAP7_75t_L g3366 ( 
.A(n_3119),
.B(n_3050),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3351),
.A2(n_3103),
.B(n_3088),
.Y(n_3367)
);

AOI22xp5_ASAP7_75t_SL g3368 ( 
.A1(n_3329),
.A2(n_3166),
.B1(n_3183),
.B2(n_3088),
.Y(n_3368)
);

OAI211xp5_ASAP7_75t_SL g3369 ( 
.A1(n_3254),
.A2(n_3075),
.B(n_3056),
.C(n_3153),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3348),
.Y(n_3370)
);

AOI22xp33_ASAP7_75t_L g3371 ( 
.A1(n_3353),
.A2(n_3056),
.B1(n_3047),
.B2(n_3026),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3247),
.Y(n_3372)
);

BUFx3_ASAP7_75t_L g3373 ( 
.A(n_3257),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3247),
.Y(n_3374)
);

O2A1O1Ixp33_ASAP7_75t_L g3375 ( 
.A1(n_3236),
.A2(n_3026),
.B(n_3146),
.C(n_2898),
.Y(n_3375)
);

OAI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3292),
.A2(n_3271),
.B1(n_3364),
.B2(n_3303),
.Y(n_3376)
);

AOI22xp5_ASAP7_75t_L g3377 ( 
.A1(n_3288),
.A2(n_3086),
.B1(n_3146),
.B2(n_3083),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3364),
.A2(n_3366),
.B1(n_3325),
.B2(n_3256),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3274),
.B(n_3202),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_3209),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_3363),
.A2(n_3083),
.B1(n_3187),
.B2(n_3197),
.Y(n_3381)
);

NAND2x1_ASAP7_75t_L g3382 ( 
.A(n_3318),
.B(n_3012),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_SL g3383 ( 
.A1(n_3308),
.A2(n_3134),
.B1(n_3114),
.B2(n_3086),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3250),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_SL g3385 ( 
.A1(n_3308),
.A2(n_3033),
.B1(n_3147),
.B2(n_3057),
.Y(n_3385)
);

NOR2x1_ASAP7_75t_SL g3386 ( 
.A(n_3259),
.B(n_3109),
.Y(n_3386)
);

AOI221xp5_ASAP7_75t_L g3387 ( 
.A1(n_3219),
.A2(n_2810),
.B1(n_2993),
.B2(n_3147),
.C(n_3036),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_3224),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3250),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_3348),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3220),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_SL g3392 ( 
.A1(n_3271),
.A2(n_3304),
.B1(n_3328),
.B2(n_3360),
.Y(n_3392)
);

BUFx6f_ASAP7_75t_L g3393 ( 
.A(n_3224),
.Y(n_3393)
);

HB1xp67_ASAP7_75t_L g3394 ( 
.A(n_3209),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3360),
.A2(n_3094),
.B1(n_3098),
.B2(n_3062),
.Y(n_3395)
);

BUFx2_ASAP7_75t_L g3396 ( 
.A(n_3305),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3252),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3220),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3294),
.B(n_3144),
.Y(n_3399)
);

AOI221xp5_ASAP7_75t_L g3400 ( 
.A1(n_3219),
.A2(n_2810),
.B1(n_3057),
.B2(n_3033),
.C(n_3122),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3252),
.Y(n_3401)
);

INVx3_ASAP7_75t_L g3402 ( 
.A(n_3330),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3253),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3363),
.A2(n_3347),
.B1(n_3232),
.B2(n_3306),
.Y(n_3404)
);

OAI22xp5_ASAP7_75t_L g3405 ( 
.A1(n_3366),
.A2(n_3050),
.B1(n_3020),
.B2(n_3045),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3306),
.B(n_3298),
.Y(n_3406)
);

OAI221xp5_ASAP7_75t_L g3407 ( 
.A1(n_3271),
.A2(n_3080),
.B1(n_3156),
.B2(n_3148),
.C(n_3053),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3253),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_L g3409 ( 
.A1(n_3306),
.A2(n_3122),
.B1(n_3137),
.B2(n_3074),
.Y(n_3409)
);

BUFx3_ASAP7_75t_L g3410 ( 
.A(n_3257),
.Y(n_3410)
);

AOI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_3328),
.A2(n_3137),
.B1(n_3077),
.B2(n_3128),
.Y(n_3411)
);

INVx4_ASAP7_75t_L g3412 ( 
.A(n_3224),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3325),
.A2(n_3135),
.B1(n_3143),
.B2(n_3102),
.Y(n_3413)
);

AOI221xp5_ASAP7_75t_L g3414 ( 
.A1(n_3283),
.A2(n_3167),
.B1(n_3074),
.B2(n_2853),
.C(n_2920),
.Y(n_3414)
);

AOI22xp33_ASAP7_75t_L g3415 ( 
.A1(n_3232),
.A2(n_3111),
.B1(n_3113),
.B2(n_3093),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3325),
.A2(n_3102),
.B1(n_3123),
.B2(n_3018),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_L g3417 ( 
.A1(n_3232),
.A2(n_3061),
.B1(n_2920),
.B2(n_3108),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3258),
.Y(n_3418)
);

OAI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_3267),
.A2(n_3123),
.B1(n_3151),
.B2(n_3054),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3258),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3241),
.A2(n_3089),
.B1(n_3131),
.B2(n_3116),
.Y(n_3421)
);

OAI22xp33_ASAP7_75t_L g3422 ( 
.A1(n_3335),
.A2(n_3182),
.B1(n_3189),
.B2(n_3151),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3246),
.A2(n_3108),
.B1(n_3127),
.B2(n_2849),
.Y(n_3423)
);

NAND3xp33_ASAP7_75t_L g3424 ( 
.A(n_3243),
.B(n_3182),
.C(n_3161),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3225),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3274),
.B(n_3151),
.Y(n_3426)
);

OAI33xp33_ASAP7_75t_L g3427 ( 
.A1(n_3243),
.A2(n_3115),
.A3(n_3085),
.B1(n_3044),
.B2(n_3188),
.B3(n_91),
.Y(n_3427)
);

AOI22xp33_ASAP7_75t_L g3428 ( 
.A1(n_3246),
.A2(n_3127),
.B1(n_2849),
.B2(n_2841),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3327),
.B(n_3282),
.Y(n_3429)
);

OAI211xp5_ASAP7_75t_L g3430 ( 
.A1(n_3283),
.A2(n_3145),
.B(n_3046),
.C(n_2862),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_L g3431 ( 
.A1(n_3246),
.A2(n_3313),
.B1(n_3315),
.B2(n_3361),
.Y(n_3431)
);

A2O1A1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_3304),
.A2(n_3055),
.B(n_3165),
.C(n_2904),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3267),
.A2(n_3055),
.B1(n_3160),
.B2(n_3194),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3225),
.Y(n_3434)
);

OR2x2_ASAP7_75t_L g3435 ( 
.A(n_3240),
.B(n_2959),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3260),
.Y(n_3436)
);

OR2x2_ASAP7_75t_L g3437 ( 
.A(n_3242),
.B(n_3324),
.Y(n_3437)
);

AOI22xp33_ASAP7_75t_L g3438 ( 
.A1(n_3313),
.A2(n_2878),
.B1(n_2996),
.B2(n_2904),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_3315),
.A2(n_2996),
.B1(n_3007),
.B2(n_2956),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3327),
.B(n_3194),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_3212),
.A2(n_2862),
.B1(n_2855),
.B2(n_2996),
.Y(n_3441)
);

OAI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3267),
.A2(n_3160),
.B1(n_3194),
.B2(n_2845),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3282),
.B(n_3107),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3260),
.Y(n_3444)
);

AOI21xp33_ASAP7_75t_L g3445 ( 
.A1(n_3212),
.A2(n_3007),
.B(n_2956),
.Y(n_3445)
);

AOI22xp33_ASAP7_75t_SL g3446 ( 
.A1(n_3283),
.A2(n_2855),
.B1(n_3201),
.B2(n_2996),
.Y(n_3446)
);

OA21x2_ASAP7_75t_L g3447 ( 
.A1(n_3285),
.A2(n_2907),
.B(n_2874),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3267),
.A2(n_2845),
.B1(n_2828),
.B2(n_3107),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_SL g3449 ( 
.A1(n_3285),
.A2(n_3201),
.B1(n_2959),
.B2(n_3007),
.Y(n_3449)
);

OR2x6_ASAP7_75t_L g3450 ( 
.A(n_3259),
.B(n_2845),
.Y(n_3450)
);

HB1xp67_ASAP7_75t_L g3451 ( 
.A(n_3210),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3263),
.B(n_2871),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3210),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3262),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3257),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3208),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3218),
.B(n_2959),
.Y(n_3457)
);

CKINVDCx5p33_ASAP7_75t_R g3458 ( 
.A(n_3228),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_3212),
.A2(n_3163),
.B1(n_2966),
.B2(n_2926),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3285),
.A2(n_2980),
.B1(n_2986),
.B2(n_2962),
.Y(n_3460)
);

AOI22xp33_ASAP7_75t_L g3461 ( 
.A1(n_3335),
.A2(n_3000),
.B1(n_2999),
.B2(n_3004),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3326),
.A2(n_2842),
.B1(n_2959),
.B2(n_2924),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3263),
.B(n_3213),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3262),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_3305),
.A2(n_2933),
.B1(n_2892),
.B2(n_2902),
.Y(n_3465)
);

NOR2x1_ASAP7_75t_R g3466 ( 
.A(n_3224),
.B(n_3270),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_3249),
.Y(n_3467)
);

BUFx6f_ASAP7_75t_L g3468 ( 
.A(n_3270),
.Y(n_3468)
);

OAI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3218),
.A2(n_2816),
.B1(n_2933),
.B2(n_2892),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3208),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3330),
.B(n_89),
.Y(n_3471)
);

BUFx3_ASAP7_75t_L g3472 ( 
.A(n_3270),
.Y(n_3472)
);

OAI221xp5_ASAP7_75t_L g3473 ( 
.A1(n_3316),
.A2(n_2884),
.B1(n_2902),
.B2(n_2913),
.C(n_2842),
.Y(n_3473)
);

INVx2_ASAP7_75t_SL g3474 ( 
.A(n_3302),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3216),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3222),
.B(n_2913),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3266),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3266),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3268),
.Y(n_3479)
);

AOI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3226),
.A2(n_2884),
.B(n_2915),
.Y(n_3480)
);

HB1xp67_ASAP7_75t_L g3481 ( 
.A(n_3211),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3326),
.A2(n_2850),
.B1(n_2913),
.B2(n_2951),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3268),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3213),
.B(n_2913),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3361),
.A2(n_2850),
.B1(n_2897),
.B2(n_2795),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3278),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3216),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3361),
.A2(n_2870),
.B1(n_2869),
.B2(n_2858),
.Y(n_3488)
);

OAI21x1_ASAP7_75t_L g3489 ( 
.A1(n_3255),
.A2(n_2863),
.B(n_90),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3286),
.B(n_91),
.Y(n_3490)
);

INVx1_ASAP7_75t_SL g3491 ( 
.A(n_3248),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3278),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_3346),
.B(n_92),
.Y(n_3493)
);

AOI221xp5_ASAP7_75t_L g3494 ( 
.A1(n_3312),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.C(n_96),
.Y(n_3494)
);

OAI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3280),
.A2(n_97),
.B1(n_93),
.B2(n_95),
.Y(n_3495)
);

BUFx6f_ASAP7_75t_SL g3496 ( 
.A(n_3365),
.Y(n_3496)
);

AOI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3324),
.A2(n_987),
.B1(n_99),
.B2(n_97),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_L g3498 ( 
.A1(n_3299),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3396),
.B(n_3310),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3429),
.B(n_3310),
.Y(n_3500)
);

HB1xp67_ASAP7_75t_L g3501 ( 
.A(n_3467),
.Y(n_3501)
);

HB1xp67_ASAP7_75t_L g3502 ( 
.A(n_3467),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3371),
.B(n_3222),
.Y(n_3503)
);

BUFx3_ASAP7_75t_L g3504 ( 
.A(n_3472),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3372),
.Y(n_3505)
);

HB1xp67_ASAP7_75t_L g3506 ( 
.A(n_3374),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3384),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3389),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3402),
.B(n_3311),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3397),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3402),
.B(n_3311),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3406),
.B(n_3293),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3391),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_3463),
.B(n_3312),
.Y(n_3514)
);

NOR2x1_ASAP7_75t_L g3515 ( 
.A(n_3373),
.B(n_3330),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3380),
.Y(n_3516)
);

INVx3_ASAP7_75t_L g3517 ( 
.A(n_3393),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3380),
.Y(n_3518)
);

BUFx12f_ASAP7_75t_L g3519 ( 
.A(n_3393),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3394),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3371),
.B(n_3223),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3394),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3443),
.B(n_3320),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3427),
.A2(n_3299),
.B1(n_3345),
.B2(n_3211),
.Y(n_3524)
);

HB1xp67_ASAP7_75t_L g3525 ( 
.A(n_3401),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3398),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3425),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3451),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3434),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3367),
.B(n_3223),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3481),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3481),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3451),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3382),
.B(n_3320),
.Y(n_3534)
);

NOR2xp67_ASAP7_75t_L g3535 ( 
.A(n_3378),
.B(n_3330),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3453),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3426),
.B(n_3323),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3456),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3414),
.B(n_3227),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_R g3540 ( 
.A(n_3455),
.B(n_3302),
.Y(n_3540)
);

INVx3_ASAP7_75t_L g3541 ( 
.A(n_3393),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3453),
.Y(n_3542)
);

INVx1_ASAP7_75t_SL g3543 ( 
.A(n_3491),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_3437),
.B(n_3293),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3440),
.B(n_3323),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3403),
.Y(n_3546)
);

INVx5_ASAP7_75t_L g3547 ( 
.A(n_3393),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3408),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3452),
.B(n_3296),
.Y(n_3549)
);

NOR2xp33_ASAP7_75t_L g3550 ( 
.A(n_3468),
.B(n_3365),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3418),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3470),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3399),
.B(n_3227),
.Y(n_3553)
);

AND2x2_ASAP7_75t_L g3554 ( 
.A(n_3379),
.B(n_3296),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3468),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3475),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3420),
.Y(n_3557)
);

AND2x4_ASAP7_75t_L g3558 ( 
.A(n_3450),
.B(n_3346),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3436),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3468),
.B(n_3350),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3387),
.B(n_3231),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3487),
.Y(n_3562)
);

OAI21xp33_ASAP7_75t_L g3563 ( 
.A1(n_3409),
.A2(n_3234),
.B(n_3231),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3377),
.B(n_3234),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3444),
.Y(n_3565)
);

OR2x2_ASAP7_75t_L g3566 ( 
.A(n_3435),
.B(n_3235),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3468),
.B(n_3350),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3388),
.B(n_3314),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3370),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3412),
.B(n_3314),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3390),
.Y(n_3571)
);

AND2x2_ASAP7_75t_L g3572 ( 
.A(n_3412),
.B(n_3318),
.Y(n_3572)
);

AND2x2_ASAP7_75t_L g3573 ( 
.A(n_3392),
.B(n_3286),
.Y(n_3573)
);

AND2x4_ASAP7_75t_L g3574 ( 
.A(n_3450),
.B(n_3259),
.Y(n_3574)
);

INVxp67_ASAP7_75t_SL g3575 ( 
.A(n_3376),
.Y(n_3575)
);

NOR2xp33_ASAP7_75t_L g3576 ( 
.A(n_3466),
.B(n_3365),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3450),
.B(n_3259),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3454),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3464),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3392),
.B(n_3255),
.Y(n_3580)
);

INVx2_ASAP7_75t_SL g3581 ( 
.A(n_3410),
.Y(n_3581)
);

HB1xp67_ASAP7_75t_L g3582 ( 
.A(n_3477),
.Y(n_3582)
);

AND2x4_ASAP7_75t_L g3583 ( 
.A(n_3478),
.B(n_3479),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3483),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3490),
.B(n_3235),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3486),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_3492),
.Y(n_3587)
);

OR2x2_ASAP7_75t_L g3588 ( 
.A(n_3476),
.B(n_3237),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3457),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3489),
.Y(n_3590)
);

NOR2x1_ASAP7_75t_SL g3591 ( 
.A(n_3413),
.B(n_3259),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3447),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_3386),
.B(n_3244),
.Y(n_3593)
);

INVx1_ASAP7_75t_SL g3594 ( 
.A(n_3493),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3383),
.B(n_3255),
.Y(n_3595)
);

AOI22xp33_ASAP7_75t_SL g3596 ( 
.A1(n_3368),
.A2(n_3345),
.B1(n_3265),
.B2(n_3272),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3424),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3497),
.Y(n_3598)
);

INVx3_ASAP7_75t_L g3599 ( 
.A(n_3496),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3383),
.B(n_3255),
.Y(n_3600)
);

HB1xp67_ASAP7_75t_L g3601 ( 
.A(n_3493),
.Y(n_3601)
);

HB1xp67_ASAP7_75t_L g3602 ( 
.A(n_3447),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3484),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3385),
.B(n_3269),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3411),
.Y(n_3605)
);

INVx2_ASAP7_75t_SL g3606 ( 
.A(n_3458),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3385),
.B(n_3269),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3407),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3419),
.B(n_3269),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3474),
.B(n_3269),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3431),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3496),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3433),
.B(n_3277),
.Y(n_3613)
);

INVx4_ASAP7_75t_L g3614 ( 
.A(n_3471),
.Y(n_3614)
);

AND2x2_ASAP7_75t_L g3615 ( 
.A(n_3416),
.B(n_3277),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3415),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3473),
.Y(n_3617)
);

HB1xp67_ASAP7_75t_L g3618 ( 
.A(n_3405),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3421),
.B(n_3277),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3427),
.A2(n_3211),
.B1(n_3359),
.B2(n_3229),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3376),
.B(n_3237),
.Y(n_3621)
);

OAI22xp33_ASAP7_75t_L g3622 ( 
.A1(n_3400),
.A2(n_3356),
.B1(n_3358),
.B2(n_3355),
.Y(n_3622)
);

AOI222xp33_ASAP7_75t_L g3623 ( 
.A1(n_3369),
.A2(n_3272),
.B1(n_3265),
.B2(n_3244),
.C1(n_3334),
.C2(n_3331),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3375),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3442),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3409),
.B(n_3238),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3506),
.Y(n_3627)
);

INVx1_ASAP7_75t_SL g3628 ( 
.A(n_3543),
.Y(n_3628)
);

NAND2xp33_ASAP7_75t_R g3629 ( 
.A(n_3540),
.B(n_3217),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3611),
.A2(n_3404),
.B1(n_3441),
.B2(n_3381),
.Y(n_3630)
);

NAND2xp33_ASAP7_75t_SL g3631 ( 
.A(n_3604),
.B(n_3365),
.Y(n_3631)
);

OAI221xp5_ASAP7_75t_L g3632 ( 
.A1(n_3575),
.A2(n_3498),
.B1(n_3449),
.B2(n_3441),
.C(n_3381),
.Y(n_3632)
);

NOR2x2_ASAP7_75t_L g3633 ( 
.A(n_3625),
.B(n_3355),
.Y(n_3633)
);

AOI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_3503),
.A2(n_3430),
.B(n_3498),
.Y(n_3634)
);

AND2x4_ASAP7_75t_L g3635 ( 
.A(n_3504),
.B(n_3357),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_R g3636 ( 
.A(n_3606),
.B(n_3504),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3604),
.B(n_3228),
.Y(n_3637)
);

OAI33xp33_ASAP7_75t_L g3638 ( 
.A1(n_3561),
.A2(n_3495),
.A3(n_3215),
.B1(n_3214),
.B2(n_3238),
.B3(n_3469),
.Y(n_3638)
);

NOR3xp33_ASAP7_75t_L g3639 ( 
.A(n_3624),
.B(n_3494),
.C(n_3422),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3607),
.B(n_3302),
.Y(n_3640)
);

AND4x1_ASAP7_75t_L g3641 ( 
.A(n_3576),
.B(n_3395),
.C(n_3423),
.D(n_3340),
.Y(n_3641)
);

AO221x1_ASAP7_75t_L g3642 ( 
.A1(n_3622),
.A2(n_3422),
.B1(n_3448),
.B2(n_3339),
.C(n_3277),
.Y(n_3642)
);

OAI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_3618),
.A2(n_3446),
.B1(n_3428),
.B2(n_3432),
.Y(n_3643)
);

OAI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3521),
.A2(n_3358),
.B1(n_3356),
.B2(n_3469),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3525),
.Y(n_3645)
);

INVxp33_ASAP7_75t_L g3646 ( 
.A(n_3591),
.Y(n_3646)
);

AOI221xp5_ASAP7_75t_L g3647 ( 
.A1(n_3611),
.A2(n_3449),
.B1(n_3265),
.B2(n_3272),
.C(n_3462),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3616),
.A2(n_3446),
.B1(n_3462),
.B2(n_3459),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3607),
.B(n_3302),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3582),
.B(n_3281),
.Y(n_3650)
);

HB1xp67_ASAP7_75t_L g3651 ( 
.A(n_3501),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3584),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3606),
.Y(n_3653)
);

AOI221xp5_ASAP7_75t_L g3654 ( 
.A1(n_3624),
.A2(n_3482),
.B1(n_3459),
.B2(n_3264),
.C(n_3251),
.Y(n_3654)
);

OAI221xp5_ASAP7_75t_L g3655 ( 
.A1(n_3596),
.A2(n_3461),
.B1(n_3438),
.B2(n_3417),
.C(n_3482),
.Y(n_3655)
);

INVx2_ASAP7_75t_SL g3656 ( 
.A(n_3601),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3626),
.B(n_3214),
.Y(n_3657)
);

NAND4xp25_ASAP7_75t_L g3658 ( 
.A(n_3595),
.B(n_3488),
.C(n_3354),
.D(n_3461),
.Y(n_3658)
);

AOI221xp5_ASAP7_75t_L g3659 ( 
.A1(n_3617),
.A2(n_3264),
.B1(n_3251),
.B2(n_3230),
.C(n_3261),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3524),
.A2(n_3460),
.B1(n_3357),
.B2(n_3439),
.Y(n_3660)
);

OAI211xp5_ASAP7_75t_L g3661 ( 
.A1(n_3580),
.A2(n_3488),
.B(n_3342),
.C(n_3445),
.Y(n_3661)
);

AOI22xp33_ASAP7_75t_SL g3662 ( 
.A1(n_3617),
.A2(n_3275),
.B1(n_3233),
.B2(n_3245),
.Y(n_3662)
);

OAI211xp5_ASAP7_75t_L g3663 ( 
.A1(n_3580),
.A2(n_3595),
.B(n_3600),
.C(n_3614),
.Y(n_3663)
);

OR2x6_ASAP7_75t_L g3664 ( 
.A(n_3614),
.B(n_3480),
.Y(n_3664)
);

INVx5_ASAP7_75t_L g3665 ( 
.A(n_3519),
.Y(n_3665)
);

OR2x2_ASAP7_75t_L g3666 ( 
.A(n_3553),
.B(n_3215),
.Y(n_3666)
);

AOI221xp5_ASAP7_75t_L g3667 ( 
.A1(n_3597),
.A2(n_3251),
.B1(n_3264),
.B2(n_3261),
.C(n_3230),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3583),
.Y(n_3668)
);

OAI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_3614),
.A2(n_3598),
.B1(n_3530),
.B2(n_3573),
.Y(n_3669)
);

OAI22xp33_ASAP7_75t_L g3670 ( 
.A1(n_3621),
.A2(n_3233),
.B1(n_3362),
.B2(n_3359),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3502),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3583),
.Y(n_3672)
);

AOI21x1_ASAP7_75t_L g3673 ( 
.A1(n_3612),
.A2(n_3352),
.B(n_3332),
.Y(n_3673)
);

AOI221xp5_ASAP7_75t_L g3674 ( 
.A1(n_3563),
.A2(n_3460),
.B1(n_3276),
.B2(n_3281),
.C(n_3287),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3583),
.Y(n_3675)
);

OAI33xp33_ASAP7_75t_L g3676 ( 
.A1(n_3597),
.A2(n_3276),
.A3(n_3284),
.B1(n_3287),
.B2(n_3331),
.B3(n_3338),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3505),
.B(n_3507),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3546),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3500),
.B(n_3217),
.Y(n_3679)
);

AOI211xp5_ASAP7_75t_L g3680 ( 
.A1(n_3535),
.A2(n_3465),
.B(n_3332),
.C(n_3343),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_3608),
.A2(n_3229),
.B1(n_3275),
.B2(n_3307),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3555),
.Y(n_3682)
);

OAI221xp5_ASAP7_75t_L g3683 ( 
.A1(n_3539),
.A2(n_3275),
.B1(n_3485),
.B2(n_3233),
.C(n_3362),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_3581),
.B(n_3280),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3500),
.B(n_3217),
.Y(n_3685)
);

NAND2x1_ASAP7_75t_L g3686 ( 
.A(n_3600),
.B(n_3593),
.Y(n_3686)
);

BUFx2_ASAP7_75t_L g3687 ( 
.A(n_3519),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_R g3688 ( 
.A(n_3599),
.B(n_3581),
.Y(n_3688)
);

INVx1_ASAP7_75t_SL g3689 ( 
.A(n_3594),
.Y(n_3689)
);

OR2x2_ASAP7_75t_L g3690 ( 
.A(n_3564),
.B(n_3284),
.Y(n_3690)
);

OAI31xp33_ASAP7_75t_SL g3691 ( 
.A1(n_3573),
.A2(n_3279),
.A3(n_3245),
.B(n_3337),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_R g3692 ( 
.A(n_3599),
.B(n_3217),
.Y(n_3692)
);

BUFx3_ASAP7_75t_L g3693 ( 
.A(n_3612),
.Y(n_3693)
);

BUFx3_ASAP7_75t_L g3694 ( 
.A(n_3599),
.Y(n_3694)
);

AOI22xp33_ASAP7_75t_L g3695 ( 
.A1(n_3608),
.A2(n_3229),
.B1(n_3275),
.B2(n_3307),
.Y(n_3695)
);

OAI22xp5_ASAP7_75t_L g3696 ( 
.A1(n_3598),
.A2(n_3605),
.B1(n_3620),
.B2(n_3585),
.Y(n_3696)
);

OR2x6_ASAP7_75t_L g3697 ( 
.A(n_3515),
.B(n_3233),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3508),
.B(n_3334),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3523),
.B(n_3221),
.Y(n_3699)
);

AOI221xp5_ASAP7_75t_L g3700 ( 
.A1(n_3605),
.A2(n_3336),
.B1(n_3338),
.B2(n_3485),
.C(n_3297),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3546),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3523),
.B(n_3554),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3548),
.Y(n_3703)
);

HB1xp67_ASAP7_75t_L g3704 ( 
.A(n_3590),
.Y(n_3704)
);

AOI221xp5_ASAP7_75t_L g3705 ( 
.A1(n_3589),
.A2(n_3336),
.B1(n_3297),
.B2(n_3349),
.C(n_3343),
.Y(n_3705)
);

HB1xp67_ASAP7_75t_L g3706 ( 
.A(n_3590),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3623),
.A2(n_3362),
.B1(n_3233),
.B2(n_3337),
.Y(n_3707)
);

HB1xp67_ASAP7_75t_L g3708 ( 
.A(n_3499),
.Y(n_3708)
);

NAND4xp25_ASAP7_75t_SL g3709 ( 
.A(n_3619),
.B(n_3239),
.C(n_3291),
.D(n_3221),
.Y(n_3709)
);

NAND3xp33_ASAP7_75t_SL g3710 ( 
.A(n_3619),
.B(n_3239),
.C(n_3291),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3548),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3551),
.Y(n_3712)
);

AOI22xp33_ASAP7_75t_L g3713 ( 
.A1(n_3625),
.A2(n_3307),
.B1(n_3233),
.B2(n_3290),
.Y(n_3713)
);

NAND4xp25_ASAP7_75t_L g3714 ( 
.A(n_3550),
.B(n_3221),
.C(n_3339),
.D(n_3279),
.Y(n_3714)
);

NAND4xp25_ASAP7_75t_L g3715 ( 
.A(n_3570),
.B(n_3221),
.C(n_3339),
.D(n_3344),
.Y(n_3715)
);

INVxp67_ASAP7_75t_L g3716 ( 
.A(n_3570),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3499),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3554),
.B(n_3339),
.Y(n_3718)
);

AOI221xp5_ASAP7_75t_L g3719 ( 
.A1(n_3589),
.A2(n_3349),
.B1(n_3290),
.B2(n_3300),
.C(n_3295),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3545),
.B(n_3344),
.Y(n_3720)
);

OAI31xp33_ASAP7_75t_L g3721 ( 
.A1(n_3602),
.A2(n_3289),
.A3(n_3300),
.B(n_3295),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3551),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3557),
.Y(n_3723)
);

INVx2_ASAP7_75t_SL g3724 ( 
.A(n_3547),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3557),
.Y(n_3725)
);

HB1xp67_ASAP7_75t_L g3726 ( 
.A(n_3510),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3555),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3555),
.Y(n_3728)
);

HB1xp67_ASAP7_75t_L g3729 ( 
.A(n_3559),
.Y(n_3729)
);

INVx1_ASAP7_75t_SL g3730 ( 
.A(n_3560),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3565),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3565),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3578),
.B(n_3289),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3545),
.Y(n_3734)
);

BUFx2_ASAP7_75t_L g3735 ( 
.A(n_3560),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3514),
.B(n_3301),
.Y(n_3736)
);

BUFx3_ASAP7_75t_L g3737 ( 
.A(n_3547),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3578),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3514),
.B(n_3301),
.Y(n_3739)
);

BUFx2_ASAP7_75t_L g3740 ( 
.A(n_3567),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3537),
.Y(n_3741)
);

AND2x4_ASAP7_75t_L g3742 ( 
.A(n_3628),
.B(n_3547),
.Y(n_3742)
);

NAND3xp33_ASAP7_75t_L g3743 ( 
.A(n_3669),
.B(n_3518),
.C(n_3516),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_SL g3744 ( 
.A1(n_3642),
.A2(n_3591),
.B1(n_3592),
.B2(n_3603),
.Y(n_3744)
);

OR2x2_ASAP7_75t_L g3745 ( 
.A(n_3628),
.B(n_3544),
.Y(n_3745)
);

NAND3xp33_ASAP7_75t_L g3746 ( 
.A(n_3669),
.B(n_3518),
.C(n_3516),
.Y(n_3746)
);

OA211x2_ASAP7_75t_L g3747 ( 
.A1(n_3686),
.A2(n_3547),
.B(n_3541),
.C(n_3517),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3708),
.B(n_3537),
.Y(n_3748)
);

OAI211xp5_ASAP7_75t_L g3749 ( 
.A1(n_3663),
.A2(n_3547),
.B(n_3522),
.C(n_3528),
.Y(n_3749)
);

INVx2_ASAP7_75t_SL g3750 ( 
.A(n_3636),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3702),
.B(n_3567),
.Y(n_3751)
);

NAND3xp33_ASAP7_75t_L g3752 ( 
.A(n_3696),
.B(n_3522),
.C(n_3520),
.Y(n_3752)
);

NAND3xp33_ASAP7_75t_L g3753 ( 
.A(n_3674),
.B(n_3528),
.C(n_3520),
.Y(n_3753)
);

NOR3xp33_ASAP7_75t_L g3754 ( 
.A(n_3638),
.B(n_3541),
.C(n_3517),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3643),
.A2(n_3592),
.B(n_3536),
.Y(n_3755)
);

NOR3xp33_ASAP7_75t_SL g3756 ( 
.A(n_3631),
.B(n_3536),
.C(n_3533),
.Y(n_3756)
);

AOI221xp5_ASAP7_75t_L g3757 ( 
.A1(n_3696),
.A2(n_3603),
.B1(n_3588),
.B2(n_3532),
.C(n_3531),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3704),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3689),
.B(n_3544),
.Y(n_3759)
);

NAND3xp33_ASAP7_75t_L g3760 ( 
.A(n_3674),
.B(n_3542),
.C(n_3533),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3706),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_3689),
.B(n_3542),
.Y(n_3762)
);

NAND3xp33_ASAP7_75t_L g3763 ( 
.A(n_3632),
.B(n_3532),
.C(n_3531),
.Y(n_3763)
);

NOR3xp33_ASAP7_75t_L g3764 ( 
.A(n_3683),
.B(n_3541),
.C(n_3517),
.Y(n_3764)
);

NAND3xp33_ASAP7_75t_L g3765 ( 
.A(n_3632),
.B(n_3512),
.C(n_3586),
.Y(n_3765)
);

AND2x4_ASAP7_75t_L g3766 ( 
.A(n_3635),
.B(n_3558),
.Y(n_3766)
);

AOI22xp5_ASAP7_75t_L g3767 ( 
.A1(n_3643),
.A2(n_3593),
.B1(n_3577),
.B2(n_3574),
.Y(n_3767)
);

AND2x2_ASAP7_75t_SL g3768 ( 
.A(n_3639),
.B(n_3593),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3633),
.Y(n_3769)
);

NOR2xp33_ASAP7_75t_L g3770 ( 
.A(n_3653),
.B(n_3558),
.Y(n_3770)
);

NOR2xp33_ASAP7_75t_L g3771 ( 
.A(n_3635),
.B(n_3558),
.Y(n_3771)
);

NAND3xp33_ASAP7_75t_L g3772 ( 
.A(n_3630),
.B(n_3651),
.C(n_3634),
.Y(n_3772)
);

NAND4xp75_ASAP7_75t_L g3773 ( 
.A(n_3647),
.B(n_3615),
.C(n_3613),
.D(n_3609),
.Y(n_3773)
);

OR2x2_ASAP7_75t_L g3774 ( 
.A(n_3717),
.B(n_3588),
.Y(n_3774)
);

NOR3xp33_ASAP7_75t_L g3775 ( 
.A(n_3683),
.B(n_3512),
.C(n_3586),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3640),
.B(n_3568),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3656),
.B(n_3579),
.Y(n_3777)
);

BUFx3_ASAP7_75t_L g3778 ( 
.A(n_3687),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3735),
.Y(n_3779)
);

INVx3_ASAP7_75t_L g3780 ( 
.A(n_3737),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3649),
.B(n_3637),
.Y(n_3781)
);

AOI22xp5_ASAP7_75t_L g3782 ( 
.A1(n_3655),
.A2(n_3577),
.B1(n_3574),
.B2(n_3571),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3726),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3729),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3740),
.B(n_3568),
.Y(n_3785)
);

BUFx12f_ASAP7_75t_L g3786 ( 
.A(n_3665),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3716),
.B(n_3579),
.Y(n_3787)
);

OR2x2_ASAP7_75t_L g3788 ( 
.A(n_3690),
.B(n_3587),
.Y(n_3788)
);

OR2x2_ASAP7_75t_L g3789 ( 
.A(n_3657),
.B(n_3734),
.Y(n_3789)
);

NOR4xp75_ASAP7_75t_L g3790 ( 
.A(n_3660),
.B(n_3572),
.C(n_3615),
.D(n_3609),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3730),
.B(n_3587),
.Y(n_3791)
);

OR2x2_ASAP7_75t_L g3792 ( 
.A(n_3741),
.B(n_3730),
.Y(n_3792)
);

OR2x2_ASAP7_75t_L g3793 ( 
.A(n_3666),
.B(n_3566),
.Y(n_3793)
);

NAND3xp33_ASAP7_75t_L g3794 ( 
.A(n_3641),
.B(n_3566),
.C(n_3572),
.Y(n_3794)
);

NOR3xp33_ASAP7_75t_L g3795 ( 
.A(n_3661),
.B(n_3577),
.C(n_3574),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3684),
.B(n_3610),
.Y(n_3796)
);

OA211x2_ASAP7_75t_L g3797 ( 
.A1(n_3709),
.A2(n_3613),
.B(n_3534),
.C(n_3511),
.Y(n_3797)
);

OAI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3660),
.A2(n_3662),
.B(n_3655),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3671),
.B(n_3509),
.Y(n_3799)
);

NOR3xp33_ASAP7_75t_SL g3800 ( 
.A(n_3709),
.B(n_3534),
.C(n_3610),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3678),
.Y(n_3801)
);

NAND3xp33_ASAP7_75t_SL g3802 ( 
.A(n_3648),
.B(n_3511),
.C(n_3509),
.Y(n_3802)
);

NAND3xp33_ASAP7_75t_L g3803 ( 
.A(n_3691),
.B(n_3526),
.C(n_3513),
.Y(n_3803)
);

OR2x2_ASAP7_75t_L g3804 ( 
.A(n_3627),
.B(n_3549),
.Y(n_3804)
);

NOR3xp33_ASAP7_75t_L g3805 ( 
.A(n_3694),
.B(n_3571),
.C(n_3569),
.Y(n_3805)
);

NOR3xp33_ASAP7_75t_L g3806 ( 
.A(n_3693),
.B(n_3569),
.C(n_3549),
.Y(n_3806)
);

HB1xp67_ASAP7_75t_L g3807 ( 
.A(n_3668),
.Y(n_3807)
);

OAI211xp5_ASAP7_75t_L g3808 ( 
.A1(n_3691),
.A2(n_3526),
.B(n_3527),
.C(n_3513),
.Y(n_3808)
);

OR2x2_ASAP7_75t_L g3809 ( 
.A(n_3645),
.B(n_3538),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3684),
.B(n_3538),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3665),
.B(n_3552),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3665),
.B(n_3718),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3665),
.B(n_3699),
.Y(n_3813)
);

NAND3xp33_ASAP7_75t_L g3814 ( 
.A(n_3681),
.B(n_3529),
.C(n_3527),
.Y(n_3814)
);

NAND3xp33_ASAP7_75t_L g3815 ( 
.A(n_3695),
.B(n_3529),
.C(n_3552),
.Y(n_3815)
);

INVxp67_ASAP7_75t_L g3816 ( 
.A(n_3652),
.Y(n_3816)
);

INVx1_ASAP7_75t_SL g3817 ( 
.A(n_3688),
.Y(n_3817)
);

OAI211xp5_ASAP7_75t_SL g3818 ( 
.A1(n_3672),
.A2(n_3562),
.B(n_3556),
.C(n_101),
.Y(n_3818)
);

NOR3xp33_ASAP7_75t_L g3819 ( 
.A(n_3644),
.B(n_3562),
.C(n_3556),
.Y(n_3819)
);

BUFx3_ASAP7_75t_L g3820 ( 
.A(n_3675),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3677),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3679),
.B(n_3309),
.Y(n_3822)
);

NOR2xp33_ASAP7_75t_L g3823 ( 
.A(n_3676),
.B(n_98),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3685),
.B(n_3724),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3646),
.B(n_100),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3682),
.B(n_3309),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3710),
.B(n_101),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3658),
.A2(n_3273),
.B1(n_3319),
.B2(n_3317),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3727),
.B(n_3273),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3728),
.B(n_3317),
.Y(n_3830)
);

NOR2x1_ASAP7_75t_L g3831 ( 
.A(n_3697),
.B(n_102),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3697),
.B(n_3319),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3701),
.B(n_3321),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_3742),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3745),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3759),
.Y(n_3836)
);

AOI31xp33_ASAP7_75t_L g3837 ( 
.A1(n_3817),
.A2(n_3629),
.A3(n_3680),
.B(n_3677),
.Y(n_3837)
);

OR2x2_ASAP7_75t_L g3838 ( 
.A(n_3792),
.B(n_3650),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3798),
.A2(n_3654),
.B1(n_3700),
.B2(n_3664),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3755),
.B(n_3703),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3751),
.B(n_3750),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3823),
.B(n_3711),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3762),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3781),
.B(n_3692),
.Y(n_3844)
);

AOI33xp33_ASAP7_75t_L g3845 ( 
.A1(n_3744),
.A2(n_3722),
.A3(n_3738),
.B1(n_3712),
.B2(n_3732),
.B3(n_3731),
.Y(n_3845)
);

BUFx2_ASAP7_75t_L g3846 ( 
.A(n_3786),
.Y(n_3846)
);

O2A1O1Ixp33_ASAP7_75t_L g3847 ( 
.A1(n_3772),
.A2(n_3664),
.B(n_3725),
.C(n_3723),
.Y(n_3847)
);

OAI221xp5_ASAP7_75t_L g3848 ( 
.A1(n_3772),
.A2(n_3664),
.B1(n_3707),
.B2(n_3713),
.C(n_3721),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3774),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3742),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3778),
.Y(n_3851)
);

AOI221xp5_ASAP7_75t_L g3852 ( 
.A1(n_3765),
.A2(n_3659),
.B1(n_3667),
.B2(n_3705),
.C(n_3670),
.Y(n_3852)
);

AOI22xp5_ASAP7_75t_L g3853 ( 
.A1(n_3775),
.A2(n_3720),
.B1(n_3739),
.B2(n_3736),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3791),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3785),
.B(n_3697),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3801),
.Y(n_3856)
);

AOI221xp5_ASAP7_75t_SL g3857 ( 
.A1(n_3757),
.A2(n_3715),
.B1(n_3714),
.B2(n_3650),
.C(n_3698),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3831),
.Y(n_3858)
);

AOI22xp33_ASAP7_75t_L g3859 ( 
.A1(n_3802),
.A2(n_3733),
.B1(n_3719),
.B2(n_3698),
.Y(n_3859)
);

INVx3_ASAP7_75t_L g3860 ( 
.A(n_3766),
.Y(n_3860)
);

AOI221xp5_ASAP7_75t_SL g3861 ( 
.A1(n_3790),
.A2(n_3733),
.B1(n_3673),
.B2(n_106),
.C(n_103),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3758),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3766),
.B(n_105),
.Y(n_3863)
);

BUFx3_ASAP7_75t_L g3864 ( 
.A(n_3779),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3776),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3810),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3761),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3820),
.Y(n_3868)
);

INVx5_ASAP7_75t_L g3869 ( 
.A(n_3780),
.Y(n_3869)
);

AOI22xp33_ASAP7_75t_L g3870 ( 
.A1(n_3765),
.A2(n_3794),
.B1(n_3818),
.B2(n_3769),
.Y(n_3870)
);

NAND2x1p5_ASAP7_75t_L g3871 ( 
.A(n_3780),
.B(n_105),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3809),
.Y(n_3872)
);

OR2x2_ASAP7_75t_L g3873 ( 
.A(n_3748),
.B(n_106),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3796),
.B(n_107),
.Y(n_3874)
);

INVx2_ASAP7_75t_SL g3875 ( 
.A(n_3813),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3788),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3768),
.Y(n_3877)
);

HB1xp67_ASAP7_75t_L g3878 ( 
.A(n_3752),
.Y(n_3878)
);

AOI22xp33_ASAP7_75t_L g3879 ( 
.A1(n_3794),
.A2(n_3763),
.B1(n_3752),
.B2(n_3803),
.Y(n_3879)
);

AND2x4_ASAP7_75t_L g3880 ( 
.A(n_3770),
.B(n_3321),
.Y(n_3880)
);

OAI211xp5_ASAP7_75t_SL g3881 ( 
.A1(n_3749),
.A2(n_110),
.B(n_107),
.C(n_109),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3787),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3783),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3824),
.B(n_111),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3784),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3812),
.B(n_114),
.Y(n_3886)
);

NAND4xp25_ASAP7_75t_L g3887 ( 
.A(n_3797),
.B(n_117),
.C(n_115),
.D(n_116),
.Y(n_3887)
);

OAI22xp5_ASAP7_75t_L g3888 ( 
.A1(n_3773),
.A2(n_3341),
.B1(n_3333),
.B2(n_3322),
.Y(n_3888)
);

AOI31xp33_ASAP7_75t_L g3889 ( 
.A1(n_3816),
.A2(n_118),
.A3(n_115),
.B(n_117),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3821),
.B(n_119),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3789),
.Y(n_3891)
);

AO31x2_ASAP7_75t_L g3892 ( 
.A1(n_3825),
.A2(n_3333),
.A3(n_3341),
.B(n_3322),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3771),
.B(n_119),
.Y(n_3893)
);

INVx4_ASAP7_75t_L g3894 ( 
.A(n_3811),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3793),
.Y(n_3895)
);

AOI33xp33_ASAP7_75t_L g3896 ( 
.A1(n_3767),
.A2(n_120),
.A3(n_121),
.B1(n_122),
.B2(n_124),
.B3(n_125),
.Y(n_3896)
);

AOI222xp33_ASAP7_75t_L g3897 ( 
.A1(n_3763),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.C1(n_125),
.C2(n_127),
.Y(n_3897)
);

CKINVDCx5p33_ASAP7_75t_R g3898 ( 
.A(n_3827),
.Y(n_3898)
);

NOR3xp33_ASAP7_75t_L g3899 ( 
.A(n_3743),
.B(n_3746),
.C(n_3760),
.Y(n_3899)
);

INVx1_ASAP7_75t_SL g3900 ( 
.A(n_3807),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3804),
.Y(n_3901)
);

OAI31xp33_ASAP7_75t_SL g3902 ( 
.A1(n_3760),
.A2(n_130),
.A3(n_127),
.B(n_128),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3777),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3799),
.Y(n_3904)
);

AOI221xp5_ASAP7_75t_L g3905 ( 
.A1(n_3754),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.C(n_133),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3833),
.Y(n_3906)
);

OAI221xp5_ASAP7_75t_L g3907 ( 
.A1(n_3782),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.C(n_134),
.Y(n_3907)
);

OAI221xp5_ASAP7_75t_L g3908 ( 
.A1(n_3764),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_3908)
);

INVxp67_ASAP7_75t_L g3909 ( 
.A(n_3743),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3746),
.Y(n_3910)
);

INVx1_ASAP7_75t_SL g3911 ( 
.A(n_3832),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3756),
.B(n_135),
.Y(n_3912)
);

AOI22xp5_ASAP7_75t_L g3913 ( 
.A1(n_3803),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.Y(n_3913)
);

INVx1_ASAP7_75t_SL g3914 ( 
.A(n_3826),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3753),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3805),
.Y(n_3916)
);

BUFx3_ASAP7_75t_L g3917 ( 
.A(n_3829),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3800),
.B(n_139),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3806),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3822),
.B(n_142),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3814),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3814),
.Y(n_3922)
);

OR2x6_ASAP7_75t_L g3923 ( 
.A(n_3815),
.B(n_3808),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_SL g3924 ( 
.A(n_3795),
.B(n_987),
.Y(n_3924)
);

OAI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3747),
.A2(n_145),
.B1(n_142),
.B2(n_143),
.Y(n_3925)
);

INVx3_ASAP7_75t_SL g3926 ( 
.A(n_3886),
.Y(n_3926)
);

INVx1_ASAP7_75t_SL g3927 ( 
.A(n_3900),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3860),
.B(n_3830),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3860),
.B(n_3819),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3878),
.Y(n_3930)
);

INVx2_ASAP7_75t_SL g3931 ( 
.A(n_3841),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3878),
.Y(n_3932)
);

OR2x2_ASAP7_75t_L g3933 ( 
.A(n_3909),
.B(n_3815),
.Y(n_3933)
);

AOI32xp33_ASAP7_75t_L g3934 ( 
.A1(n_3899),
.A2(n_3828),
.A3(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3899),
.B(n_143),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3890),
.Y(n_3936)
);

INVx1_ASAP7_75t_SL g3937 ( 
.A(n_3884),
.Y(n_3937)
);

O2A1O1Ixp33_ASAP7_75t_L g3938 ( 
.A1(n_3909),
.A2(n_149),
.B(n_146),
.C(n_147),
.Y(n_3938)
);

OR2x2_ASAP7_75t_L g3939 ( 
.A(n_3901),
.B(n_149),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3871),
.Y(n_3940)
);

NAND4xp75_ASAP7_75t_L g3941 ( 
.A(n_3905),
.B(n_154),
.C(n_152),
.D(n_153),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3890),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3871),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3835),
.Y(n_3944)
);

OAI22xp5_ASAP7_75t_L g3945 ( 
.A1(n_3879),
.A2(n_3923),
.B1(n_3910),
.B2(n_3915),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3836),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3901),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3869),
.Y(n_3948)
);

AOI22xp5_ASAP7_75t_L g3949 ( 
.A1(n_3923),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3849),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3902),
.B(n_155),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3895),
.B(n_156),
.Y(n_3952)
);

INVx2_ASAP7_75t_SL g3953 ( 
.A(n_3869),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3869),
.Y(n_3954)
);

AOI21x1_ASAP7_75t_L g3955 ( 
.A1(n_3921),
.A2(n_157),
.B(n_158),
.Y(n_3955)
);

O2A1O1Ixp33_ASAP7_75t_L g3956 ( 
.A1(n_3922),
.A2(n_161),
.B(n_158),
.C(n_159),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3923),
.A2(n_3879),
.B1(n_3839),
.B2(n_3905),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3843),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3891),
.Y(n_3959)
);

OR2x2_ASAP7_75t_L g3960 ( 
.A(n_3838),
.B(n_162),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3872),
.Y(n_3961)
);

OAI22xp33_ASAP7_75t_L g3962 ( 
.A1(n_3848),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3914),
.B(n_163),
.Y(n_3963)
);

AND2x4_ASAP7_75t_L g3964 ( 
.A(n_3868),
.B(n_165),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3873),
.Y(n_3965)
);

OR2x2_ASAP7_75t_L g3966 ( 
.A(n_3840),
.B(n_165),
.Y(n_3966)
);

AOI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3839),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_3967)
);

NAND2x1_ASAP7_75t_SL g3968 ( 
.A(n_3855),
.B(n_167),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3861),
.B(n_171),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3844),
.B(n_171),
.Y(n_3970)
);

A2O1A1Ixp33_ASAP7_75t_L g3971 ( 
.A1(n_3845),
.A2(n_3913),
.B(n_3847),
.C(n_3870),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3876),
.Y(n_3972)
);

OAI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3870),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3847),
.A2(n_175),
.B(n_176),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3840),
.B(n_175),
.Y(n_3975)
);

AOI32xp33_ASAP7_75t_L g3976 ( 
.A1(n_3881),
.A2(n_177),
.A3(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_3976)
);

AND2x4_ASAP7_75t_L g3977 ( 
.A(n_3864),
.B(n_177),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3920),
.Y(n_3978)
);

NAND2x1_ASAP7_75t_SL g3979 ( 
.A(n_3912),
.B(n_178),
.Y(n_3979)
);

AND2x4_ASAP7_75t_L g3980 ( 
.A(n_3834),
.B(n_182),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3874),
.B(n_182),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3856),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3882),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3862),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3869),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3846),
.B(n_183),
.Y(n_3986)
);

OR2x2_ASAP7_75t_L g3987 ( 
.A(n_3865),
.B(n_183),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3917),
.Y(n_3988)
);

OR2x2_ASAP7_75t_L g3989 ( 
.A(n_3842),
.B(n_184),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3897),
.B(n_185),
.Y(n_3990)
);

AOI22xp5_ASAP7_75t_L g3991 ( 
.A1(n_3848),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3896),
.B(n_186),
.Y(n_3992)
);

OAI22xp33_ASAP7_75t_L g3993 ( 
.A1(n_3837),
.A2(n_187),
.B1(n_189),
.B2(n_191),
.Y(n_3993)
);

AOI211xp5_ASAP7_75t_L g3994 ( 
.A1(n_3881),
.A2(n_3887),
.B(n_3925),
.C(n_3908),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3867),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3858),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3896),
.B(n_189),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3854),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3863),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3889),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3883),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3866),
.B(n_3911),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3851),
.B(n_191),
.Y(n_4003)
);

AOI32xp33_ASAP7_75t_L g4004 ( 
.A1(n_3859),
.A2(n_192),
.A3(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_4004)
);

OR2x2_ASAP7_75t_L g4005 ( 
.A(n_3842),
.B(n_192),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3885),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3903),
.Y(n_4007)
);

INVxp67_ASAP7_75t_L g4008 ( 
.A(n_3924),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3906),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3894),
.B(n_194),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3904),
.Y(n_4011)
);

OAI32xp33_ASAP7_75t_L g4012 ( 
.A1(n_3925),
.A2(n_195),
.A3(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3845),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3893),
.B(n_200),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3916),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3937),
.B(n_3918),
.Y(n_4016)
);

INVx1_ASAP7_75t_SL g4017 ( 
.A(n_3979),
.Y(n_4017)
);

HB1xp67_ASAP7_75t_L g4018 ( 
.A(n_3931),
.Y(n_4018)
);

CKINVDCx16_ASAP7_75t_R g4019 ( 
.A(n_3927),
.Y(n_4019)
);

HB1xp67_ASAP7_75t_L g4020 ( 
.A(n_3930),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3966),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3975),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3926),
.B(n_3875),
.Y(n_4023)
);

AND2x4_ASAP7_75t_L g4024 ( 
.A(n_3928),
.B(n_3894),
.Y(n_4024)
);

INVx3_ASAP7_75t_SL g4025 ( 
.A(n_3977),
.Y(n_4025)
);

OR2x2_ASAP7_75t_L g4026 ( 
.A(n_3945),
.B(n_3850),
.Y(n_4026)
);

HB1xp67_ASAP7_75t_L g4027 ( 
.A(n_3930),
.Y(n_4027)
);

NOR3xp33_ASAP7_75t_SL g4028 ( 
.A(n_3971),
.B(n_3919),
.C(n_3898),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3960),
.Y(n_4029)
);

INVx1_ASAP7_75t_SL g4030 ( 
.A(n_3933),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3968),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3955),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_3964),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3970),
.B(n_3877),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3986),
.B(n_3857),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3980),
.B(n_3859),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_4014),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_3988),
.B(n_3853),
.Y(n_4038)
);

OR2x2_ASAP7_75t_L g4039 ( 
.A(n_3947),
.B(n_3908),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3980),
.B(n_3880),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3939),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3964),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3977),
.Y(n_4043)
);

NAND2xp33_ASAP7_75t_L g4044 ( 
.A(n_4000),
.B(n_3888),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3952),
.Y(n_4045)
);

BUFx2_ASAP7_75t_L g4046 ( 
.A(n_3928),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3981),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_4000),
.B(n_3880),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3965),
.Y(n_4049)
);

NOR2x1_ASAP7_75t_L g4050 ( 
.A(n_3935),
.B(n_3907),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3944),
.B(n_3888),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3963),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_4002),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3976),
.B(n_3907),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3978),
.Y(n_4055)
);

NOR2xp67_ASAP7_75t_SL g4056 ( 
.A(n_3987),
.B(n_3852),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3994),
.B(n_3852),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_3940),
.B(n_201),
.Y(n_4058)
);

AOI222xp33_ASAP7_75t_L g4059 ( 
.A1(n_4013),
.A2(n_3892),
.B1(n_203),
.B2(n_205),
.C1(n_207),
.C2(n_208),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3959),
.Y(n_4060)
);

AND2x4_ASAP7_75t_L g4061 ( 
.A(n_3943),
.B(n_3892),
.Y(n_4061)
);

OAI21xp33_ASAP7_75t_L g4062 ( 
.A1(n_4013),
.A2(n_3892),
.B(n_202),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3932),
.Y(n_4063)
);

OAI32xp33_ASAP7_75t_L g4064 ( 
.A1(n_3973),
.A2(n_3969),
.A3(n_3951),
.B1(n_3990),
.B2(n_4005),
.Y(n_4064)
);

CKINVDCx5p33_ASAP7_75t_R g4065 ( 
.A(n_4003),
.Y(n_4065)
);

NOR4xp25_ASAP7_75t_L g4066 ( 
.A(n_4015),
.B(n_3892),
.C(n_203),
.D(n_205),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3972),
.Y(n_4067)
);

OR2x2_ASAP7_75t_L g4068 ( 
.A(n_3946),
.B(n_202),
.Y(n_4068)
);

NAND4xp25_ASAP7_75t_L g4069 ( 
.A(n_3957),
.B(n_207),
.C(n_208),
.D(n_209),
.Y(n_4069)
);

INVx1_ASAP7_75t_SL g4070 ( 
.A(n_3929),
.Y(n_4070)
);

OR2x6_ASAP7_75t_L g4071 ( 
.A(n_3996),
.B(n_209),
.Y(n_4071)
);

OR2x6_ASAP7_75t_L g4072 ( 
.A(n_3953),
.B(n_210),
.Y(n_4072)
);

INVxp67_ASAP7_75t_SL g4073 ( 
.A(n_3993),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3936),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_4010),
.B(n_210),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3942),
.Y(n_4076)
);

CKINVDCx16_ASAP7_75t_R g4077 ( 
.A(n_3989),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_3999),
.B(n_211),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_4004),
.B(n_211),
.Y(n_4079)
);

INVxp67_ASAP7_75t_L g4080 ( 
.A(n_3941),
.Y(n_4080)
);

OR2x2_ASAP7_75t_L g4081 ( 
.A(n_3958),
.B(n_212),
.Y(n_4081)
);

INVx1_ASAP7_75t_SL g4082 ( 
.A(n_3992),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3950),
.B(n_213),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_4012),
.B(n_213),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3948),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3961),
.B(n_214),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3934),
.B(n_214),
.Y(n_4087)
);

NOR2x1_ASAP7_75t_L g4088 ( 
.A(n_3954),
.B(n_215),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_4011),
.B(n_216),
.Y(n_4089)
);

OR2x2_ASAP7_75t_L g4090 ( 
.A(n_3998),
.B(n_216),
.Y(n_4090)
);

OR2x2_ASAP7_75t_L g4091 ( 
.A(n_3983),
.B(n_217),
.Y(n_4091)
);

AND2x4_ASAP7_75t_L g4092 ( 
.A(n_3985),
.B(n_217),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_4007),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3997),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4015),
.Y(n_4095)
);

NAND4xp25_ASAP7_75t_L g4096 ( 
.A(n_3991),
.B(n_218),
.C(n_220),
.D(n_221),
.Y(n_4096)
);

CKINVDCx6p67_ASAP7_75t_R g4097 ( 
.A(n_3984),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3982),
.Y(n_4098)
);

OAI21xp5_ASAP7_75t_L g4099 ( 
.A1(n_3949),
.A2(n_218),
.B(n_222),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4019),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_4077),
.B(n_3974),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_4046),
.B(n_4009),
.Y(n_4102)
);

NOR2x1_ASAP7_75t_L g4103 ( 
.A(n_4072),
.B(n_3956),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_4030),
.B(n_3995),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_4025),
.B(n_4012),
.Y(n_4105)
);

OAI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_4057),
.A2(n_4030),
.B(n_4088),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4018),
.Y(n_4107)
);

A2O1A1Ixp33_ASAP7_75t_L g4108 ( 
.A1(n_4062),
.A2(n_3967),
.B(n_3938),
.C(n_4001),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4020),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_4023),
.B(n_4006),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4037),
.B(n_3962),
.Y(n_4111)
);

INVxp67_ASAP7_75t_L g4112 ( 
.A(n_4031),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4027),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4070),
.B(n_4008),
.Y(n_4114)
);

OR2x2_ASAP7_75t_L g4115 ( 
.A(n_4070),
.B(n_4097),
.Y(n_4115)
);

NAND3xp33_ASAP7_75t_L g4116 ( 
.A(n_4028),
.B(n_223),
.C(n_225),
.Y(n_4116)
);

INVx2_ASAP7_75t_SL g4117 ( 
.A(n_4024),
.Y(n_4117)
);

XNOR2x2_ASAP7_75t_L g4118 ( 
.A(n_4069),
.B(n_225),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_4024),
.B(n_226),
.Y(n_4119)
);

XNOR2xp5_ASAP7_75t_L g4120 ( 
.A(n_4065),
.B(n_227),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4072),
.Y(n_4121)
);

AOI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_4044),
.A2(n_228),
.B(n_229),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_4035),
.B(n_228),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4092),
.B(n_230),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4072),
.Y(n_4125)
);

INVxp67_ASAP7_75t_L g4126 ( 
.A(n_4056),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4083),
.Y(n_4127)
);

XNOR2xp5_ASAP7_75t_L g4128 ( 
.A(n_4034),
.B(n_230),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_4092),
.B(n_231),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4086),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_4038),
.B(n_233),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_4048),
.B(n_233),
.Y(n_4132)
);

INVxp67_ASAP7_75t_SL g4133 ( 
.A(n_4026),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_4053),
.B(n_235),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_4055),
.B(n_235),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_4049),
.B(n_236),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4089),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_4043),
.B(n_236),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4094),
.B(n_238),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4068),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4081),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_4016),
.B(n_238),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4090),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_4017),
.B(n_239),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_4071),
.Y(n_4145)
);

INVx1_ASAP7_75t_SL g4146 ( 
.A(n_4017),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4091),
.Y(n_4147)
);

INVxp67_ASAP7_75t_L g4148 ( 
.A(n_4036),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_4085),
.B(n_239),
.Y(n_4149)
);

NOR2x1_ASAP7_75t_R g4150 ( 
.A(n_4075),
.B(n_240),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4032),
.Y(n_4151)
);

AND2x4_ASAP7_75t_L g4152 ( 
.A(n_4060),
.B(n_240),
.Y(n_4152)
);

AND2x4_ASAP7_75t_L g4153 ( 
.A(n_4067),
.B(n_242),
.Y(n_4153)
);

AND2x4_ASAP7_75t_L g4154 ( 
.A(n_4098),
.B(n_243),
.Y(n_4154)
);

OAI21xp33_ASAP7_75t_L g4155 ( 
.A1(n_4050),
.A2(n_4082),
.B(n_4051),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4021),
.Y(n_4156)
);

OR2x2_ASAP7_75t_L g4157 ( 
.A(n_4039),
.B(n_243),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_4069),
.B(n_245),
.Y(n_4158)
);

NOR2x1_ASAP7_75t_L g4159 ( 
.A(n_4063),
.B(n_245),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4066),
.B(n_246),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4022),
.B(n_246),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4029),
.Y(n_4162)
);

XNOR2xp5_ASAP7_75t_L g4163 ( 
.A(n_4096),
.B(n_247),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_4082),
.B(n_248),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_4084),
.B(n_4041),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_4058),
.B(n_249),
.Y(n_4166)
);

AOI32xp33_ASAP7_75t_L g4167 ( 
.A1(n_4103),
.A2(n_4062),
.A3(n_4095),
.B1(n_4076),
.B2(n_4074),
.Y(n_4167)
);

OR2x6_ASAP7_75t_L g4168 ( 
.A(n_4100),
.B(n_4144),
.Y(n_4168)
);

OAI221xp5_ASAP7_75t_L g4169 ( 
.A1(n_4155),
.A2(n_4066),
.B1(n_4059),
.B2(n_4054),
.C(n_4073),
.Y(n_4169)
);

AOI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_4146),
.A2(n_4052),
.B1(n_4047),
.B2(n_4059),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4133),
.Y(n_4171)
);

INVx3_ASAP7_75t_L g4172 ( 
.A(n_4119),
.Y(n_4172)
);

OAI21xp33_ASAP7_75t_L g4173 ( 
.A1(n_4105),
.A2(n_4064),
.B(n_4093),
.Y(n_4173)
);

INVx1_ASAP7_75t_SL g4174 ( 
.A(n_4115),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4128),
.Y(n_4175)
);

NAND3xp33_ASAP7_75t_L g4176 ( 
.A(n_4126),
.B(n_4106),
.C(n_4116),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4150),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4150),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4154),
.B(n_4033),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4154),
.B(n_4042),
.Y(n_4180)
);

NAND2x1p5_ASAP7_75t_L g4181 ( 
.A(n_4117),
.B(n_4119),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_SL g4182 ( 
.A1(n_4146),
.A2(n_4045),
.B1(n_4040),
.B2(n_4061),
.Y(n_4182)
);

AOI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_4155),
.A2(n_4080),
.B1(n_4087),
.B2(n_4096),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4120),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4102),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_4132),
.B(n_4071),
.Y(n_4186)
);

AOI321xp33_ASAP7_75t_L g4187 ( 
.A1(n_4151),
.A2(n_4061),
.A3(n_4079),
.B1(n_4078),
.B2(n_4071),
.C(n_4099),
.Y(n_4187)
);

OAI221xp5_ASAP7_75t_L g4188 ( 
.A1(n_4106),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.C(n_252),
.Y(n_4188)
);

NAND2xp33_ASAP7_75t_SL g4189 ( 
.A(n_4104),
.B(n_250),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4157),
.Y(n_4190)
);

AOI22xp33_ASAP7_75t_L g4191 ( 
.A1(n_4148),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_4110),
.B(n_253),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_4132),
.B(n_255),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4123),
.Y(n_4194)
);

INVx1_ASAP7_75t_SL g4195 ( 
.A(n_4101),
.Y(n_4195)
);

INVxp67_ASAP7_75t_L g4196 ( 
.A(n_4131),
.Y(n_4196)
);

NAND3xp33_ASAP7_75t_L g4197 ( 
.A(n_4116),
.B(n_255),
.C(n_256),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4163),
.Y(n_4198)
);

OAI22x1_ASAP7_75t_L g4199 ( 
.A1(n_4112),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_4114),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4107),
.B(n_260),
.Y(n_4201)
);

AOI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_4160),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_4152),
.B(n_261),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4124),
.Y(n_4204)
);

OAI21xp33_ASAP7_75t_L g4205 ( 
.A1(n_4165),
.A2(n_264),
.B(n_265),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4129),
.Y(n_4206)
);

OAI21xp33_ASAP7_75t_L g4207 ( 
.A1(n_4121),
.A2(n_264),
.B(n_265),
.Y(n_4207)
);

AOI31xp33_ASAP7_75t_L g4208 ( 
.A1(n_4162),
.A2(n_266),
.A3(n_267),
.B(n_268),
.Y(n_4208)
);

AOI22xp5_ASAP7_75t_L g4209 ( 
.A1(n_4160),
.A2(n_4137),
.B1(n_4130),
.B2(n_4127),
.Y(n_4209)
);

INVx2_ASAP7_75t_SL g4210 ( 
.A(n_4135),
.Y(n_4210)
);

AOI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_4139),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4134),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4152),
.B(n_270),
.Y(n_4213)
);

OR2x2_ASAP7_75t_L g4214 ( 
.A(n_4109),
.B(n_271),
.Y(n_4214)
);

OAI21xp33_ASAP7_75t_SL g4215 ( 
.A1(n_4113),
.A2(n_4156),
.B(n_4125),
.Y(n_4215)
);

AOI21xp33_ASAP7_75t_L g4216 ( 
.A1(n_4159),
.A2(n_272),
.B(n_273),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4153),
.B(n_272),
.Y(n_4217)
);

AOI22xp33_ASAP7_75t_L g4218 ( 
.A1(n_4140),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_4218)
);

OAI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_4108),
.A2(n_274),
.B(n_275),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4153),
.B(n_276),
.Y(n_4220)
);

AOI221xp5_ASAP7_75t_L g4221 ( 
.A1(n_4122),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.C(n_281),
.Y(n_4221)
);

AOI21xp33_ASAP7_75t_L g4222 ( 
.A1(n_4145),
.A2(n_277),
.B(n_280),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4149),
.B(n_281),
.Y(n_4223)
);

INVx1_ASAP7_75t_SL g4224 ( 
.A(n_4118),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4136),
.Y(n_4225)
);

INVx1_ASAP7_75t_SL g4226 ( 
.A(n_4111),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4141),
.B(n_4143),
.Y(n_4227)
);

XNOR2x2_ASAP7_75t_L g4228 ( 
.A(n_4158),
.B(n_282),
.Y(n_4228)
);

AOI222xp33_ASAP7_75t_L g4229 ( 
.A1(n_4147),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.C1(n_285),
.C2(n_286),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4142),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4164),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4166),
.B(n_283),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4172),
.B(n_4161),
.Y(n_4233)
);

AOI21xp33_ASAP7_75t_SL g4234 ( 
.A1(n_4181),
.A2(n_4138),
.B(n_287),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4172),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4171),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4192),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4179),
.Y(n_4238)
);

HB1xp67_ASAP7_75t_L g4239 ( 
.A(n_4168),
.Y(n_4239)
);

AOI22xp5_ASAP7_75t_L g4240 ( 
.A1(n_4195),
.A2(n_285),
.B1(n_289),
.B2(n_290),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4180),
.Y(n_4241)
);

INVx2_ASAP7_75t_SL g4242 ( 
.A(n_4168),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4194),
.B(n_289),
.Y(n_4243)
);

INVxp33_ASAP7_75t_L g4244 ( 
.A(n_4186),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4210),
.B(n_290),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4208),
.B(n_291),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4185),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4174),
.B(n_292),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_4224),
.B(n_293),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4182),
.B(n_4230),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4228),
.Y(n_4251)
);

NOR2xp33_ASAP7_75t_L g4252 ( 
.A(n_4176),
.B(n_293),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4177),
.B(n_294),
.Y(n_4253)
);

O2A1O1Ixp33_ASAP7_75t_L g4254 ( 
.A1(n_4215),
.A2(n_294),
.B(n_295),
.C(n_296),
.Y(n_4254)
);

OAI211xp5_ASAP7_75t_L g4255 ( 
.A1(n_4167),
.A2(n_295),
.B(n_296),
.C(n_297),
.Y(n_4255)
);

NOR2x1_ASAP7_75t_L g4256 ( 
.A(n_4168),
.B(n_297),
.Y(n_4256)
);

OAI22xp5_ASAP7_75t_L g4257 ( 
.A1(n_4169),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4178),
.B(n_298),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4193),
.Y(n_4259)
);

AOI321xp33_ASAP7_75t_L g4260 ( 
.A1(n_4170),
.A2(n_299),
.A3(n_300),
.B1(n_301),
.B2(n_302),
.C(n_303),
.Y(n_4260)
);

OAI31xp33_ASAP7_75t_L g4261 ( 
.A1(n_4189),
.A2(n_4173),
.A3(n_4231),
.B(n_4197),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4201),
.B(n_301),
.Y(n_4262)
);

A2O1A1Ixp33_ASAP7_75t_L g4263 ( 
.A1(n_4183),
.A2(n_302),
.B(n_303),
.C(n_304),
.Y(n_4263)
);

AOI32xp33_ASAP7_75t_L g4264 ( 
.A1(n_4184),
.A2(n_305),
.A3(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_4264)
);

INVx1_ASAP7_75t_SL g4265 ( 
.A(n_4214),
.Y(n_4265)
);

XNOR2xp5_ASAP7_75t_L g4266 ( 
.A(n_4209),
.B(n_305),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4225),
.B(n_309),
.Y(n_4267)
);

INVx2_ASAP7_75t_SL g4268 ( 
.A(n_4227),
.Y(n_4268)
);

AOI22xp5_ASAP7_75t_L g4269 ( 
.A1(n_4212),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_L g4270 ( 
.A(n_4216),
.B(n_312),
.Y(n_4270)
);

AOI21xp33_ASAP7_75t_L g4271 ( 
.A1(n_4226),
.A2(n_315),
.B(n_317),
.Y(n_4271)
);

INVx3_ASAP7_75t_L g4272 ( 
.A(n_4203),
.Y(n_4272)
);

O2A1O1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_4219),
.A2(n_315),
.B(n_319),
.C(n_320),
.Y(n_4273)
);

HB1xp67_ASAP7_75t_L g4274 ( 
.A(n_4199),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4229),
.B(n_4190),
.Y(n_4275)
);

INVx2_ASAP7_75t_SL g4276 ( 
.A(n_4213),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4217),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4220),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4196),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4223),
.Y(n_4280)
);

XNOR2x2_ASAP7_75t_L g4281 ( 
.A(n_4188),
.B(n_319),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4211),
.B(n_321),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4232),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4175),
.B(n_321),
.Y(n_4284)
);

INVxp67_ASAP7_75t_L g4285 ( 
.A(n_4204),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4202),
.B(n_323),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4206),
.B(n_4205),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_SL g4288 ( 
.A(n_4242),
.B(n_4187),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4239),
.Y(n_4289)
);

NOR3xp33_ASAP7_75t_SL g4290 ( 
.A(n_4255),
.B(n_4198),
.C(n_4200),
.Y(n_4290)
);

INVx2_ASAP7_75t_L g4291 ( 
.A(n_4256),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4235),
.B(n_4268),
.Y(n_4292)
);

CKINVDCx14_ASAP7_75t_R g4293 ( 
.A(n_4248),
.Y(n_4293)
);

INVx1_ASAP7_75t_SL g4294 ( 
.A(n_4262),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4265),
.B(n_4207),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4274),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4246),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4265),
.B(n_4221),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4251),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4237),
.B(n_4191),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4250),
.Y(n_4301)
);

HB1xp67_ASAP7_75t_L g4302 ( 
.A(n_4266),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4233),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4233),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4234),
.B(n_4218),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_4249),
.Y(n_4306)
);

OR2x6_ASAP7_75t_L g4307 ( 
.A(n_4279),
.B(n_4222),
.Y(n_4307)
);

AOI22xp5_ASAP7_75t_L g4308 ( 
.A1(n_4257),
.A2(n_324),
.B1(n_325),
.B2(n_329),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4247),
.B(n_4238),
.Y(n_4309)
);

INVx1_ASAP7_75t_SL g4310 ( 
.A(n_4284),
.Y(n_4310)
);

OR2x2_ASAP7_75t_L g4311 ( 
.A(n_4241),
.B(n_329),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4260),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4272),
.B(n_330),
.Y(n_4313)
);

NAND4xp25_ASAP7_75t_L g4314 ( 
.A(n_4261),
.B(n_332),
.C(n_333),
.D(n_334),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_L g4315 ( 
.A(n_4271),
.B(n_332),
.Y(n_4315)
);

INVx1_ASAP7_75t_SL g4316 ( 
.A(n_4267),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4267),
.Y(n_4317)
);

AOI211xp5_ASAP7_75t_L g4318 ( 
.A1(n_4257),
.A2(n_335),
.B(n_336),
.C(n_337),
.Y(n_4318)
);

CKINVDCx5p33_ASAP7_75t_R g4319 ( 
.A(n_4280),
.Y(n_4319)
);

OAI322xp33_ASAP7_75t_L g4320 ( 
.A1(n_4285),
.A2(n_335),
.A3(n_337),
.B1(n_339),
.B2(n_340),
.C1(n_341),
.C2(n_343),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4272),
.Y(n_4321)
);

INVxp67_ASAP7_75t_L g4322 ( 
.A(n_4252),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4275),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4281),
.Y(n_4324)
);

AOI22xp33_ASAP7_75t_L g4325 ( 
.A1(n_4276),
.A2(n_339),
.B1(n_341),
.B2(n_343),
.Y(n_4325)
);

OA21x2_ASAP7_75t_L g4326 ( 
.A1(n_4271),
.A2(n_344),
.B(n_345),
.Y(n_4326)
);

AND2x2_ASAP7_75t_L g4327 ( 
.A(n_4236),
.B(n_345),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4245),
.Y(n_4328)
);

NOR2xp33_ASAP7_75t_L g4329 ( 
.A(n_4293),
.B(n_4244),
.Y(n_4329)
);

NOR3xp33_ASAP7_75t_L g4330 ( 
.A(n_4288),
.B(n_4253),
.C(n_4258),
.Y(n_4330)
);

NOR3x1_ASAP7_75t_L g4331 ( 
.A(n_4314),
.B(n_4243),
.C(n_4282),
.Y(n_4331)
);

OAI21xp5_ASAP7_75t_L g4332 ( 
.A1(n_4301),
.A2(n_4254),
.B(n_4273),
.Y(n_4332)
);

AOI22xp5_ASAP7_75t_L g4333 ( 
.A1(n_4289),
.A2(n_4323),
.B1(n_4297),
.B2(n_4299),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4292),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4326),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4326),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_4314),
.B(n_4263),
.Y(n_4337)
);

AOI211xp5_ASAP7_75t_L g4338 ( 
.A1(n_4296),
.A2(n_4287),
.B(n_4277),
.C(n_4278),
.Y(n_4338)
);

NOR3xp33_ASAP7_75t_L g4339 ( 
.A(n_4303),
.B(n_4283),
.C(n_4259),
.Y(n_4339)
);

AO22x2_ASAP7_75t_L g4340 ( 
.A1(n_4294),
.A2(n_4286),
.B1(n_4282),
.B2(n_4264),
.Y(n_4340)
);

OA22x2_ASAP7_75t_L g4341 ( 
.A1(n_4308),
.A2(n_4324),
.B1(n_4304),
.B2(n_4321),
.Y(n_4341)
);

AOI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_4310),
.A2(n_4270),
.B1(n_4240),
.B2(n_4269),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4291),
.Y(n_4343)
);

AOI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_4310),
.A2(n_346),
.B1(n_347),
.B2(n_490),
.Y(n_4344)
);

AOI211xp5_ASAP7_75t_L g4345 ( 
.A1(n_4309),
.A2(n_346),
.B(n_347),
.C(n_379),
.Y(n_4345)
);

OA22x2_ASAP7_75t_L g4346 ( 
.A1(n_4312),
.A2(n_4319),
.B1(n_4307),
.B2(n_4295),
.Y(n_4346)
);

AO21x1_ASAP7_75t_L g4347 ( 
.A1(n_4313),
.A2(n_382),
.B(n_385),
.Y(n_4347)
);

NAND3xp33_ASAP7_75t_L g4348 ( 
.A(n_4318),
.B(n_386),
.C(n_387),
.Y(n_4348)
);

AOI211xp5_ASAP7_75t_L g4349 ( 
.A1(n_4316),
.A2(n_389),
.B(n_391),
.C(n_392),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4311),
.Y(n_4350)
);

INVxp67_ASAP7_75t_L g4351 ( 
.A(n_4315),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4327),
.Y(n_4352)
);

AO21x1_ASAP7_75t_L g4353 ( 
.A1(n_4300),
.A2(n_393),
.B(n_394),
.Y(n_4353)
);

OAI22xp33_ASAP7_75t_L g4354 ( 
.A1(n_4333),
.A2(n_4307),
.B1(n_4305),
.B2(n_4316),
.Y(n_4354)
);

AOI22x1_ASAP7_75t_L g4355 ( 
.A1(n_4334),
.A2(n_4317),
.B1(n_4302),
.B2(n_4328),
.Y(n_4355)
);

AOI22xp33_ASAP7_75t_L g4356 ( 
.A1(n_4330),
.A2(n_4306),
.B1(n_4307),
.B2(n_4322),
.Y(n_4356)
);

OAI21xp5_ASAP7_75t_SL g4357 ( 
.A1(n_4329),
.A2(n_4298),
.B(n_4325),
.Y(n_4357)
);

CKINVDCx20_ASAP7_75t_R g4358 ( 
.A(n_4342),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4341),
.B(n_4290),
.Y(n_4359)
);

OAI21xp5_ASAP7_75t_SL g4360 ( 
.A1(n_4343),
.A2(n_4320),
.B(n_396),
.Y(n_4360)
);

NOR2x1_ASAP7_75t_L g4361 ( 
.A(n_4335),
.B(n_395),
.Y(n_4361)
);

HB1xp67_ASAP7_75t_L g4362 ( 
.A(n_4336),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4346),
.B(n_399),
.Y(n_4363)
);

OAI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_4337),
.A2(n_401),
.B1(n_405),
.B2(n_407),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_SL g4365 ( 
.A(n_4338),
.B(n_408),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4340),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4340),
.Y(n_4367)
);

AOI21xp33_ASAP7_75t_L g4368 ( 
.A1(n_4351),
.A2(n_411),
.B(n_412),
.Y(n_4368)
);

OAI32xp33_ASAP7_75t_L g4369 ( 
.A1(n_4339),
.A2(n_489),
.A3(n_418),
.B1(n_421),
.B2(n_425),
.Y(n_4369)
);

NOR4xp25_ASAP7_75t_L g4370 ( 
.A(n_4354),
.B(n_4332),
.C(n_4350),
.D(n_4352),
.Y(n_4370)
);

AOI221xp5_ASAP7_75t_L g4371 ( 
.A1(n_4362),
.A2(n_4353),
.B1(n_4348),
.B2(n_4347),
.C(n_4345),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4359),
.Y(n_4372)
);

HB1xp67_ASAP7_75t_L g4373 ( 
.A(n_4366),
.Y(n_4373)
);

AOI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4367),
.A2(n_4344),
.B1(n_4349),
.B2(n_4331),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4358),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4361),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4355),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4363),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4365),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4360),
.Y(n_4380)
);

NAND2x1p5_ASAP7_75t_L g4381 ( 
.A(n_4377),
.B(n_4356),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4375),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4373),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4376),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_R g4385 ( 
.A(n_4372),
.B(n_4357),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_4370),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4378),
.Y(n_4387)
);

NOR2x1_ASAP7_75t_L g4388 ( 
.A(n_4382),
.B(n_4380),
.Y(n_4388)
);

NAND2x1p5_ASAP7_75t_L g4389 ( 
.A(n_4383),
.B(n_4384),
.Y(n_4389)
);

INVx1_ASAP7_75t_SL g4390 ( 
.A(n_4386),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4381),
.Y(n_4391)
);

NAND2xp33_ASAP7_75t_L g4392 ( 
.A(n_4385),
.B(n_4379),
.Y(n_4392)
);

AOI211xp5_ASAP7_75t_L g4393 ( 
.A1(n_4390),
.A2(n_4387),
.B(n_4371),
.C(n_4374),
.Y(n_4393)
);

OAI211xp5_ASAP7_75t_L g4394 ( 
.A1(n_4388),
.A2(n_4374),
.B(n_4369),
.C(n_4368),
.Y(n_4394)
);

XNOR2xp5_ASAP7_75t_L g4395 ( 
.A(n_4393),
.B(n_4391),
.Y(n_4395)
);

OAI22xp5_ASAP7_75t_SL g4396 ( 
.A1(n_4394),
.A2(n_4389),
.B1(n_4392),
.B2(n_4364),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4395),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4397),
.Y(n_4398)
);

OAI221xp5_ASAP7_75t_SL g4399 ( 
.A1(n_4398),
.A2(n_4396),
.B1(n_4364),
.B2(n_433),
.C(n_436),
.Y(n_4399)
);

AOI21xp5_ASAP7_75t_L g4400 ( 
.A1(n_4399),
.A2(n_415),
.B(n_427),
.Y(n_4400)
);

OAI221xp5_ASAP7_75t_L g4401 ( 
.A1(n_4400),
.A2(n_487),
.B1(n_440),
.B2(n_441),
.C(n_445),
.Y(n_4401)
);

OAI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4401),
.A2(n_439),
.B(n_446),
.Y(n_4402)
);

XNOR2xp5_ASAP7_75t_L g4403 ( 
.A(n_4402),
.B(n_448),
.Y(n_4403)
);

OAI321xp33_ASAP7_75t_L g4404 ( 
.A1(n_4403),
.A2(n_451),
.A3(n_453),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4403),
.B(n_461),
.Y(n_4405)
);

AOI22xp33_ASAP7_75t_L g4406 ( 
.A1(n_4405),
.A2(n_464),
.B1(n_467),
.B2(n_468),
.Y(n_4406)
);

NAND2xp67_ASAP7_75t_L g4407 ( 
.A(n_4404),
.B(n_470),
.Y(n_4407)
);

INVx4_ASAP7_75t_L g4408 ( 
.A(n_4407),
.Y(n_4408)
);

OR2x6_ASAP7_75t_L g4409 ( 
.A(n_4406),
.B(n_471),
.Y(n_4409)
);

AOI221xp5_ASAP7_75t_L g4410 ( 
.A1(n_4408),
.A2(n_472),
.B1(n_475),
.B2(n_477),
.C(n_480),
.Y(n_4410)
);

AOI211xp5_ASAP7_75t_L g4411 ( 
.A1(n_4410),
.A2(n_4409),
.B(n_485),
.C(n_486),
.Y(n_4411)
);


endmodule