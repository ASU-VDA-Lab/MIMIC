module fake_jpeg_10275_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_23),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_10),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_43),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_12),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_14),
.B(n_13),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_42),
.C(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_52),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_35),
.B1(n_37),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_22),
.B1(n_24),
.B2(n_45),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_13),
.B(n_41),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_52),
.C(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_24),
.B1(n_21),
.B2(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_55),
.C(n_39),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_65),
.C(n_50),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_39),
.C(n_34),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_19),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_68),
.B1(n_21),
.B2(n_34),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_17),
.B1(n_21),
.B2(n_4),
.Y(n_75)
);

AOI321xp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_0),
.A3(n_1),
.B1(n_4),
.B2(n_73),
.C(n_7),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_1),
.Y(n_77)
);


endmodule