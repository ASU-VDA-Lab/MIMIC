module fake_jpeg_12169_n_133 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_5),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_28),
.B(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_31),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_38),
.B1(n_29),
.B2(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_13),
.B(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_56),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_20),
.B1(n_23),
.B2(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_40),
.B1(n_25),
.B2(n_2),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_61),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_29),
.A2(n_15),
.B(n_24),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_65),
.B(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_69),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_23),
.C(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_13),
.B1(n_27),
.B2(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_25),
.B1(n_67),
.B2(n_49),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_59),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_78),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_81),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_61),
.B1(n_69),
.B2(n_52),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_51),
.B(n_53),
.C(n_62),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_58),
.B(n_65),
.C(n_67),
.D(n_70),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_97),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_64),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_83),
.B(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_106),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_100),
.C(n_96),
.Y(n_112)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_78),
.C(n_73),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.C(n_95),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_76),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_73),
.B1(n_84),
.B2(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_99),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_111),
.C(n_89),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.C(n_108),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_72),
.C(n_76),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_105),
.C(n_94),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_93),
.B1(n_110),
.B2(n_88),
.Y(n_122)
);

OAI211xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_123),
.B(n_112),
.C(n_92),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_105),
.B1(n_119),
.B2(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_90),
.C(n_82),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_128),
.C(n_74),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_125),
.B(n_63),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.C(n_74),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_52),
.B1(n_60),
.B2(n_63),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_60),
.Y(n_133)
);


endmodule