module fake_ariane_1597_n_1766 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1766);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1766;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_94),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_13),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_11),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_37),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_57),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_76),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_37),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_7),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_25),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_55),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_45),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_44),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_112),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_65),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_47),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_48),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_87),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_14),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_146),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_72),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_41),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_23),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_116),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_105),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_46),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_102),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_148),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_124),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_139),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_92),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_77),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_75),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_6),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_95),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_162),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_70),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_81),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_126),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_80),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_154),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_73),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_3),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_165),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_62),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_18),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_143),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_88),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_52),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_41),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_110),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_26),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_5),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_152),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_28),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_101),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_134),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_93),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_158),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_130),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_122),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_19),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_34),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_61),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_137),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_50),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_40),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_69),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_114),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_153),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_29),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_91),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_40),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_24),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_4),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_131),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_136),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_30),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_78),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_118),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_49),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_150),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_47),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_99),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_98),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_82),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_132),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_27),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_157),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_67),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_85),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_60),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_145),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_20),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_54),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_133),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_35),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_21),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_27),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_83),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_164),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_10),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_144),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_56),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_16),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_0),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_29),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_123),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_135),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_128),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_115),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_4),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_163),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_50),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_38),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_167),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_156),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_39),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_63),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_43),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_2),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_51),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_90),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_35),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_74),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_169),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_265),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_222),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_264),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_239),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_258),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_171),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_312),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_172),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_172),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_203),
.B(n_1),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_322),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_215),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_246),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_240),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_253),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_207),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_209),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_259),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_288),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_240),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_260),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_203),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_298),
.B(n_5),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_171),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_234),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_293),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_263),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_268),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_274),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_276),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_173),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_277),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_181),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_278),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_283),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_6),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_286),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_173),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_188),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_305),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_188),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_181),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_233),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_256),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_245),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_238),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_174),
.B(n_7),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_245),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_170),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_289),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_296),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_316),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_189),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_285),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_177),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_189),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_294),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_180),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_184),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_214),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_176),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_190),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_297),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_316),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_230),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_244),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_331),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_175),
.B(n_182),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_395),
.B(n_254),
.Y(n_420)
);

INVxp33_ASAP7_75t_SL g421 ( 
.A(n_340),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_341),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_341),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_338),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_378),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_385),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_357),
.B(n_301),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_369),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_359),
.B(n_254),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_315),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_357),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g448 ( 
.A1(n_388),
.A2(n_198),
.B(n_186),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_363),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_390),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_363),
.B(n_375),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_315),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_351),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_375),
.B(n_229),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_352),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_397),
.B(n_206),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_352),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_366),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_380),
.B(n_330),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_349),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_403),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_406),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_360),
.B(n_314),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_361),
.B(n_314),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

INVx6_ASAP7_75t_L g484 ( 
.A(n_353),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_368),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_208),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_391),
.A2(n_241),
.B1(n_323),
.B2(n_308),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_R g494 ( 
.A(n_421),
.B(n_345),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_440),
.B(n_389),
.Y(n_495)
);

BUFx8_ASAP7_75t_SL g496 ( 
.A(n_447),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_484),
.A2(n_401),
.B1(n_383),
.B2(n_367),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_484),
.A2(n_404),
.B1(n_411),
.B2(n_281),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_425),
.B(n_348),
.Y(n_501)
);

OAI21xp33_ASAP7_75t_SL g502 ( 
.A1(n_440),
.A2(n_415),
.B(n_414),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_428),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_487),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_469),
.B(n_365),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_426),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_372),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_487),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_473),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_425),
.B(n_409),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_476),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_473),
.B(n_373),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_487),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_447),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_473),
.B(n_374),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_447),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_480),
.B(n_377),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_480),
.B(n_379),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_429),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_473),
.B(n_381),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_421),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_479),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_479),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_492),
.A2(n_337),
.B1(n_371),
.B2(n_343),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_469),
.B(n_382),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_432),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_482),
.B(n_384),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_487),
.B(n_304),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_423),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_482),
.B(n_398),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_492),
.A2(n_439),
.B1(n_484),
.B2(n_477),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_439),
.B(n_415),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_479),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_444),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_477),
.B(n_399),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_475),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_487),
.B(n_304),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_483),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_443),
.B(n_412),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_450),
.B(n_441),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_444),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_444),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_445),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_448),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_433),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_485),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_416),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_484),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_L g575 ( 
.A(n_420),
.B(n_292),
.C(n_201),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_441),
.B(n_402),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_435),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_484),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_489),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_444),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_444),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_489),
.B(n_304),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_484),
.B(n_362),
.Y(n_584)
);

AND2x6_ASAP7_75t_L g585 ( 
.A(n_483),
.B(n_227),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_484),
.A2(n_269),
.B1(n_318),
.B2(n_317),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_444),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_446),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_446),
.Y(n_589)
);

AO21x2_ASAP7_75t_L g590 ( 
.A1(n_420),
.A2(n_211),
.B(n_210),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_435),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_446),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_450),
.B(n_364),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_481),
.B(n_418),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_483),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_445),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_462),
.B(n_178),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_489),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_464),
.A2(n_308),
.B1(n_195),
.B2(n_197),
.Y(n_600)
);

INVx8_ASAP7_75t_L g601 ( 
.A(n_441),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_489),
.B(n_304),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_435),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_488),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_489),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_438),
.B(n_355),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_446),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_446),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_489),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_488),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_455),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_438),
.B(n_405),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_435),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_489),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_446),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_423),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_455),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_442),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_446),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_446),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_464),
.B(n_190),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_445),
.B(n_178),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_448),
.B(n_247),
.Y(n_625)
);

AND3x1_ASAP7_75t_L g626 ( 
.A(n_468),
.B(n_251),
.C(n_250),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_474),
.B(n_227),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_445),
.B(n_179),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_456),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_456),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_456),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_474),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_456),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_474),
.Y(n_635)
);

INVxp67_ASAP7_75t_R g636 ( 
.A(n_478),
.Y(n_636)
);

INVx6_ASAP7_75t_L g637 ( 
.A(n_491),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_454),
.B(n_218),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_442),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_454),
.B(n_339),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_456),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_478),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_456),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_573),
.B(n_491),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_625),
.A2(n_448),
.B1(n_491),
.B2(n_436),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_572),
.B(n_491),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_495),
.B(n_491),
.C(n_490),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_561),
.B(n_491),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_573),
.B(n_491),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_579),
.A2(n_195),
.B1(n_313),
.B2(n_306),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_522),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_601),
.B(n_491),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_490),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_552),
.B(n_486),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_497),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_525),
.B(n_347),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_601),
.B(n_478),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_601),
.B(n_478),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_499),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_499),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_563),
.B(n_486),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_563),
.B(n_486),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_563),
.B(n_486),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_579),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_498),
.A2(n_310),
.B1(n_300),
.B2(n_306),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_507),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_514),
.B(n_468),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_506),
.B(n_350),
.Y(n_669)
);

BUFx6f_ASAP7_75t_SL g670 ( 
.A(n_593),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_468),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_542),
.B(n_354),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_514),
.B(n_468),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_501),
.B(n_356),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_552),
.B(n_358),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_503),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_522),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_606),
.B(n_471),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_558),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_509),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_527),
.A2(n_550),
.B1(n_529),
.B2(n_594),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_594),
.B(n_468),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_504),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_613),
.B(n_434),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_613),
.B(n_434),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_569),
.B(n_456),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_619),
.B(n_508),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_619),
.B(n_434),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_569),
.B(n_456),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_501),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_504),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_558),
.B(n_436),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_553),
.B(n_387),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_513),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_519),
.B(n_437),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_584),
.B(n_460),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_523),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_523),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_569),
.B(n_179),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_496),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_513),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_526),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_524),
.B(n_437),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_521),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_640),
.B(n_458),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_534),
.B(n_437),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_618),
.B(n_541),
.Y(n_707)
);

AND2x6_ASAP7_75t_SL g708 ( 
.A(n_494),
.B(n_262),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_526),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_530),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_574),
.B(n_183),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_630),
.A2(n_448),
.B(n_453),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_638),
.B(n_453),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_574),
.B(n_453),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_496),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_521),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_530),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_531),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_633),
.A2(n_448),
.B(n_458),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_528),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_606),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_574),
.B(n_459),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_597),
.B(n_604),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_606),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_535),
.B(n_459),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_625),
.B(n_183),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_512),
.A2(n_471),
.B(n_448),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_551),
.A2(n_460),
.B1(n_470),
.B2(n_463),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_511),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_618),
.B(n_304),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_565),
.B(n_557),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_546),
.B(n_584),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_528),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_584),
.A2(n_202),
.B1(n_334),
.B2(n_302),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_571),
.B(n_199),
.C(n_197),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_541),
.B(n_185),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_471),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_606),
.B(n_463),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_541),
.B(n_304),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_511),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_532),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_541),
.B(n_304),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_593),
.B(n_517),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_584),
.B(n_199),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_531),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_533),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_465),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_541),
.B(n_185),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_598),
.B(n_300),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_532),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_636),
.B(n_465),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_636),
.B(n_571),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_578),
.B(n_187),
.Y(n_753)
);

NAND2x1_ASAP7_75t_L g754 ( 
.A(n_637),
.B(n_424),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_515),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_590),
.A2(n_470),
.B1(n_472),
.B2(n_467),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_549),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_518),
.B(n_442),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_536),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_590),
.A2(n_472),
.B1(n_467),
.B2(n_466),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_536),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_538),
.B(n_442),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_539),
.B(n_449),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_562),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_535),
.B(n_309),
.C(n_279),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_554),
.B(n_449),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_540),
.B(n_310),
.Y(n_767)
);

OR2x2_ASAP7_75t_SL g768 ( 
.A(n_500),
.B(n_293),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_578),
.B(n_582),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_533),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_549),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_537),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_576),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_560),
.B(n_595),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_590),
.B(n_449),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_637),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_577),
.B(n_449),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_608),
.Y(n_778)
);

INVx4_ASAP7_75t_SL g779 ( 
.A(n_585),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_502),
.B(n_313),
.Y(n_780)
);

NOR2x1p5_ASAP7_75t_L g781 ( 
.A(n_623),
.B(n_323),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_577),
.B(n_451),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_591),
.B(n_451),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_493),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_562),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_537),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_591),
.B(n_451),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_586),
.A2(n_472),
.B1(n_467),
.B2(n_466),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_614),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_SL g790 ( 
.A(n_600),
.B(n_325),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_575),
.B(n_626),
.C(n_570),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_578),
.B(n_187),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_637),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_603),
.B(n_461),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_603),
.B(n_451),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_608),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_615),
.B(n_452),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_615),
.B(n_452),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_568),
.A2(n_452),
.B(n_457),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_543),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_620),
.B(n_452),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_543),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_620),
.B(n_461),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_567),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_567),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_570),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_624),
.A2(n_334),
.B1(n_204),
.B2(n_336),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_639),
.A2(n_457),
.B(n_467),
.C(n_466),
.Y(n_808)
);

INVxp33_ASAP7_75t_L g809 ( 
.A(n_544),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_578),
.B(n_191),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_639),
.B(n_457),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_637),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_635),
.Y(n_813)
);

AOI21x1_ASAP7_75t_L g814 ( 
.A1(n_686),
.A2(n_642),
.B(n_564),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_679),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_646),
.A2(n_648),
.B(n_769),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_651),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_681),
.A2(n_628),
.B1(n_580),
.B2(n_556),
.Y(n_818)
);

BUFx12f_ASAP7_75t_L g819 ( 
.A(n_708),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_667),
.Y(n_820)
);

OAI321xp33_ASAP7_75t_L g821 ( 
.A1(n_767),
.A2(n_461),
.A3(n_466),
.B1(n_472),
.B2(n_457),
.C(n_419),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_696),
.B(n_578),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_654),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_705),
.A2(n_545),
.B(n_544),
.C(n_516),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_657),
.Y(n_825)
);

BUFx8_ASAP7_75t_L g826 ( 
.A(n_670),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_696),
.B(n_582),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_769),
.A2(n_596),
.B(n_568),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_780),
.A2(n_545),
.B(n_510),
.C(n_516),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_686),
.A2(n_596),
.B(n_568),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_682),
.B(n_505),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_689),
.A2(n_596),
.B(n_510),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_682),
.B(n_505),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_680),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_655),
.B(n_505),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_727),
.A2(n_689),
.B(n_808),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_690),
.B(n_510),
.Y(n_837)
);

OAI321xp33_ASAP7_75t_L g838 ( 
.A1(n_666),
.A2(n_461),
.A3(n_419),
.B1(n_212),
.B2(n_282),
.C(n_221),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_694),
.A2(n_329),
.B1(n_326),
.B2(n_325),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_808),
.A2(n_564),
.B(n_555),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_699),
.A2(n_566),
.B(n_555),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_696),
.B(n_582),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_653),
.A2(n_556),
.B(n_516),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_655),
.B(n_556),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_677),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_701),
.A2(n_329),
.B1(n_326),
.B2(n_599),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_704),
.A2(n_605),
.B1(n_580),
.B2(n_599),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_752),
.B(n_582),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_712),
.A2(n_581),
.B(n_566),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_790),
.A2(n_616),
.B(n_599),
.C(n_580),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_751),
.B(n_605),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_716),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_719),
.A2(n_588),
.B(n_581),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_752),
.B(n_674),
.C(n_711),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_751),
.B(n_605),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_693),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_695),
.A2(n_616),
.B(n_607),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_778),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_743),
.B(n_607),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_675),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_700),
.B(n_588),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_720),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_722),
.B(n_687),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_692),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_747),
.B(n_714),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_SL g866 ( 
.A(n_715),
.B(n_242),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_692),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_703),
.B(n_607),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_726),
.A2(n_610),
.B(n_589),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_781),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_721),
.B(n_582),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_733),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_731),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_706),
.A2(n_616),
.B(n_610),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_724),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_713),
.A2(n_617),
.B(n_589),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_732),
.B(n_669),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_672),
.B(n_493),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_741),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_744),
.A2(n_643),
.B1(n_641),
.B2(n_634),
.Y(n_881)
);

OA22x2_ASAP7_75t_L g882 ( 
.A1(n_773),
.A2(n_333),
.B1(n_641),
.B2(n_634),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_768),
.B(n_643),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_726),
.A2(n_632),
.B1(n_631),
.B2(n_629),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_SL g885 ( 
.A(n_755),
.B(n_243),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_784),
.A2(n_632),
.B(n_631),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_670),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_699),
.A2(n_629),
.B(n_621),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_711),
.B(n_493),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_784),
.A2(n_621),
.B(n_617),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_749),
.A2(n_602),
.B1(n_559),
.B2(n_547),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_654),
.Y(n_892)
);

NAND2x1_ASAP7_75t_L g893 ( 
.A(n_678),
.B(n_587),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_665),
.A2(n_547),
.B(n_559),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_652),
.A2(n_583),
.B(n_602),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_662),
.A2(n_583),
.B(n_261),
.C(n_249),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_725),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_750),
.B(n_587),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_730),
.A2(n_592),
.B(n_622),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_654),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_730),
.A2(n_592),
.B(n_622),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_759),
.B(n_587),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_658),
.A2(n_592),
.B(n_622),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_724),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_761),
.B(n_587),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_678),
.B(n_587),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_424),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_659),
.A2(n_622),
.B(n_609),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_764),
.A2(n_592),
.B(n_622),
.C(n_609),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_774),
.A2(n_609),
.B(n_592),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_777),
.A2(n_609),
.B(n_611),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_789),
.B(n_424),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_782),
.A2(n_609),
.B(n_611),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_775),
.A2(n_419),
.B(n_422),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_785),
.B(n_520),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_678),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_721),
.B(n_520),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_783),
.A2(n_611),
.B(n_520),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_654),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_787),
.A2(n_611),
.B(n_520),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_663),
.A2(n_228),
.B(n_232),
.C(n_236),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_804),
.A2(n_272),
.B(n_311),
.C(n_287),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_734),
.B(n_520),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_805),
.A2(n_493),
.B1(n_611),
.B2(n_548),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_796),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_SL g926 ( 
.A1(n_644),
.A2(n_303),
.B(n_290),
.C(n_291),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_799),
.A2(n_548),
.B(n_585),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_791),
.B(n_548),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_735),
.B(n_424),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_724),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_736),
.A2(n_319),
.B(n_295),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_806),
.B(n_548),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_650),
.B(n_548),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_645),
.A2(n_422),
.B(n_424),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_795),
.A2(n_191),
.B(n_192),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_797),
.A2(n_192),
.B(n_193),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_647),
.A2(n_422),
.B(n_321),
.C(n_205),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_668),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_664),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_723),
.A2(n_671),
.B(n_673),
.C(n_738),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_737),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_684),
.B(n_422),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_656),
.Y(n_943)
);

AO21x1_ASAP7_75t_L g944 ( 
.A1(n_736),
.A2(n_753),
.B(n_748),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_798),
.A2(n_193),
.B(n_194),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_794),
.B(n_255),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_794),
.B(n_585),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_801),
.A2(n_194),
.B(n_196),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_813),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_811),
.A2(n_196),
.B(n_200),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_758),
.A2(n_200),
.B(n_204),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_L g952 ( 
.A1(n_807),
.A2(n_328),
.B(n_205),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_728),
.B(n_299),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_809),
.B(n_299),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_803),
.B(n_660),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_685),
.A2(n_688),
.B(n_644),
.C(n_649),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_660),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_678),
.A2(n_302),
.B1(n_307),
.B2(n_336),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_762),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_661),
.B(n_8),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_763),
.A2(n_307),
.B(n_320),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_809),
.A2(n_328),
.B(n_327),
.C(n_324),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_766),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_788),
.B(n_320),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_724),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_661),
.B(n_585),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_729),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_748),
.B(n_327),
.Y(n_968)
);

OAI321xp33_ASAP7_75t_L g969 ( 
.A1(n_756),
.A2(n_227),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C(n_14),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_707),
.A2(n_248),
.B1(n_216),
.B2(n_217),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_683),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_740),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_757),
.B(n_213),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_753),
.Y(n_974)
);

BUFx4f_ASAP7_75t_L g975 ( 
.A(n_729),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_683),
.A2(n_226),
.B(n_225),
.C(n_223),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_691),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_707),
.A2(n_267),
.B(n_220),
.Y(n_978)
);

BUFx4f_ASAP7_75t_L g979 ( 
.A(n_729),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_691),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_676),
.B(n_585),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_697),
.B(n_9),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_757),
.B(n_227),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_697),
.A2(n_270),
.B(n_231),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_698),
.A2(n_271),
.B(n_235),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_698),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_702),
.A2(n_273),
.B(n_237),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_L g988 ( 
.A(n_729),
.B(n_585),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_SL g989 ( 
.A(n_757),
.B(n_266),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_792),
.A2(n_15),
.B(n_17),
.C(n_19),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_709),
.A2(n_275),
.B(n_252),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_709),
.A2(n_219),
.B(n_257),
.C(n_280),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_771),
.B(n_284),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_710),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_740),
.B(n_15),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_710),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_717),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_717),
.B(n_627),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_876),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_845),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_817),
.Y(n_1001)
);

INVxp33_ASAP7_75t_SL g1002 ( 
.A(n_825),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_975),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_941),
.A2(n_771),
.B1(n_760),
.B2(n_810),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_975),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_860),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_854),
.A2(n_810),
.B(n_792),
.C(n_754),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_939),
.B(n_770),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_867),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_820),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_979),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_924),
.A2(n_739),
.B(n_742),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_865),
.A2(n_812),
.B1(n_776),
.B2(n_793),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_878),
.B(n_772),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_943),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_959),
.B(n_963),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_868),
.B(n_718),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_864),
.B(n_718),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_874),
.B(n_812),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_815),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_863),
.B(n_802),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_856),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_879),
.B(n_776),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_955),
.B(n_802),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_924),
.A2(n_739),
.B(n_742),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_858),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_983),
.B(n_793),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_940),
.A2(n_990),
.B(n_839),
.C(n_897),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_839),
.A2(n_800),
.B1(n_786),
.B2(n_772),
.C(n_770),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_938),
.A2(n_800),
.B(n_786),
.C(n_746),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_887),
.B(n_779),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_826),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_925),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_826),
.Y(n_1034)
);

BUFx8_ASAP7_75t_L g1035 ( 
.A(n_819),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_955),
.B(n_746),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_866),
.B(n_745),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_974),
.B(n_885),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_834),
.A2(n_745),
.B1(n_227),
.B2(n_22),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_928),
.A2(n_779),
.B(n_627),
.C(n_304),
.Y(n_1040)
);

AO22x1_ASAP7_75t_L g1041 ( 
.A1(n_953),
.A2(n_627),
.B1(n_779),
.B2(n_22),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_907),
.B(n_20),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_922),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_912),
.B(n_30),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_852),
.B(n_627),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_916),
.B(n_627),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_889),
.A2(n_627),
.B(n_32),
.C(n_33),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_972),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_957),
.Y(n_1049)
);

BUFx8_ASAP7_75t_L g1050 ( 
.A(n_871),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_816),
.A2(n_68),
.B(n_147),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_862),
.B(n_31),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_869),
.A2(n_64),
.B(n_142),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_969),
.B(n_31),
.C(n_33),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_876),
.Y(n_1055)
);

OR2x6_ASAP7_75t_SL g1056 ( 
.A(n_846),
.B(n_34),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_979),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_904),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_946),
.B(n_873),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_850),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_883),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_R g1062 ( 
.A(n_973),
.B(n_89),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_837),
.A2(n_36),
.B(n_44),
.C(n_45),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_946),
.B(n_46),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_846),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_995),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_880),
.B(n_53),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_949),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_954),
.B(n_53),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_964),
.B(n_54),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_899),
.A2(n_79),
.B(n_96),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_962),
.A2(n_97),
.B(n_104),
.C(n_107),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_960),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_958),
.B(n_108),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_901),
.A2(n_109),
.B(n_117),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_982),
.B(n_119),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_823),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_831),
.B(n_138),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_848),
.B(n_168),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_822),
.B(n_827),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_956),
.A2(n_838),
.B(n_921),
.C(n_821),
.Y(n_1081)
);

NAND2x1_ASAP7_75t_L g1082 ( 
.A(n_904),
.B(n_930),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_835),
.A2(n_844),
.B1(n_891),
.B2(n_902),
.Y(n_1083)
);

OAI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_952),
.A2(n_855),
.B(n_851),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_906),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_971),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_994),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_977),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_910),
.A2(n_875),
.B(n_877),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_823),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_842),
.B(n_861),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_898),
.A2(n_902),
.B1(n_905),
.B2(n_847),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_898),
.A2(n_905),
.B1(n_847),
.B2(n_906),
.Y(n_1093)
);

AO32x1_ASAP7_75t_L g1094 ( 
.A1(n_980),
.A2(n_986),
.A3(n_996),
.B1(n_997),
.B2(n_944),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_857),
.A2(n_830),
.B(n_832),
.Y(n_1095)
);

OAI22x1_ASAP7_75t_L g1096 ( 
.A1(n_881),
.A2(n_818),
.B1(n_923),
.B2(n_970),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_882),
.B(n_968),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_823),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_829),
.A2(n_824),
.B(n_937),
.C(n_976),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_831),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_833),
.B(n_859),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_833),
.A2(n_933),
.B1(n_893),
.B2(n_942),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_947),
.B(n_965),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_989),
.B(n_900),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_892),
.Y(n_1105)
);

AO21x1_ASAP7_75t_L g1106 ( 
.A1(n_870),
.A2(n_836),
.B(n_915),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_947),
.A2(n_909),
.B1(n_915),
.B2(n_932),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_836),
.B(n_932),
.C(n_951),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_993),
.B(n_919),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_828),
.A2(n_843),
.B(n_913),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_961),
.A2(n_948),
.B(n_935),
.C(n_945),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_911),
.A2(n_918),
.B(n_920),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_896),
.A2(n_870),
.B(n_936),
.C(n_950),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_882),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_SL g1115 ( 
.A1(n_931),
.A2(n_840),
.B(n_849),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_894),
.A2(n_908),
.B(n_903),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_930),
.B(n_965),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_929),
.A2(n_895),
.B(n_927),
.C(n_840),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_884),
.A2(n_849),
.B1(n_853),
.B2(n_872),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_900),
.B(n_967),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_853),
.A2(n_890),
.B(n_886),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_SL g1122 ( 
.A(n_978),
.B(n_985),
.C(n_991),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_926),
.A2(n_917),
.B(n_987),
.C(n_984),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_900),
.B(n_967),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_927),
.A2(n_981),
.B(n_966),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_919),
.B(n_966),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_919),
.B(n_998),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_934),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_R g1129 ( 
.A(n_988),
.B(n_914),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_814),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_998),
.B(n_841),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_888),
.A2(n_924),
.B(n_646),
.Y(n_1132)
);

BUFx2_ASAP7_75t_SL g1133 ( 
.A(n_815),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_SL g1134 ( 
.A(n_845),
.B(n_535),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_854),
.A2(n_495),
.B(n_690),
.C(n_542),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_R g1136 ( 
.A(n_825),
.B(n_494),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_825),
.A2(n_681),
.B1(n_674),
.B2(n_522),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_940),
.A2(n_824),
.B(n_831),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_878),
.B(n_681),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_878),
.B(n_681),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_878),
.B(n_681),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_876),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_941),
.A2(n_681),
.B1(n_865),
.B2(n_863),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_924),
.A2(n_646),
.B(n_730),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_817),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_868),
.B(n_447),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_SL g1147 ( 
.A1(n_1139),
.A2(n_1140),
.B(n_1141),
.C(n_1082),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1014),
.B(n_1143),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1002),
.B(n_1137),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1150)
);

AND3x4_ASAP7_75t_L g1151 ( 
.A(n_1000),
.B(n_1054),
.C(n_1056),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1069),
.A2(n_1028),
.B(n_1135),
.C(n_1081),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1063),
.B(n_1065),
.C(n_1060),
.Y(n_1153)
);

CKINVDCx9p33_ASAP7_75t_R g1154 ( 
.A(n_1033),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1143),
.A2(n_1144),
.B(n_1118),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1066),
.A2(n_1064),
.B(n_1043),
.C(n_1047),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1039),
.A2(n_1004),
.B(n_1102),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1068),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1010),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1016),
.B(n_1059),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1089),
.A2(n_1095),
.B(n_1092),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1070),
.A2(n_1074),
.B1(n_1039),
.B2(n_1038),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1001),
.B(n_1145),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_1101),
.A2(n_1117),
.B(n_1113),
.C(n_1100),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1007),
.A2(n_1084),
.B(n_1016),
.C(n_1108),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1042),
.A2(n_1109),
.B(n_1076),
.C(n_1080),
.Y(n_1166)
);

AO32x2_ASAP7_75t_L g1167 ( 
.A1(n_1092),
.A2(n_1093),
.A3(n_1119),
.B1(n_1004),
.B2(n_1083),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1093),
.A2(n_1006),
.B1(n_1101),
.B2(n_1102),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1132),
.A2(n_1083),
.B(n_1138),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1022),
.B(n_1061),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1136),
.B(n_1048),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1020),
.B(n_1009),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1057),
.B(n_1085),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1079),
.A2(n_1099),
.B(n_1111),
.C(n_1072),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1073),
.B(n_1017),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1030),
.A2(n_1052),
.B(n_1025),
.C(n_1012),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1106),
.A2(n_1130),
.A3(n_1119),
.B(n_1107),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1107),
.A2(n_1121),
.A3(n_1096),
.B(n_1125),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1018),
.B(n_1133),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_SL g1180 ( 
.A(n_1062),
.B(n_1026),
.C(n_1034),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1077),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1086),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1105),
.B(n_1011),
.Y(n_1183)
);

AO32x2_ASAP7_75t_L g1184 ( 
.A1(n_1013),
.A2(n_1094),
.A3(n_1115),
.B1(n_1114),
.B2(n_1128),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1021),
.B(n_1090),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1078),
.A2(n_1051),
.B(n_1023),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1052),
.A2(n_1044),
.B(n_1067),
.Y(n_1187)
);

NAND2x1p5_ASAP7_75t_L g1188 ( 
.A(n_1003),
.B(n_1005),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1031),
.B(n_1005),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1088),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_1024),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1123),
.A2(n_1097),
.B(n_1091),
.C(n_1078),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1050),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1117),
.A2(n_1013),
.B(n_1103),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1015),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1094),
.A2(n_1024),
.A3(n_1036),
.B(n_1008),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1011),
.B(n_1037),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1011),
.B(n_1104),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1049),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1036),
.B(n_1019),
.Y(n_1200)
);

BUFx4_ASAP7_75t_SL g1201 ( 
.A(n_1035),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1103),
.A2(n_1053),
.B(n_1075),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1050),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1058),
.B(n_1120),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_SL g1205 ( 
.A1(n_1027),
.A2(n_1120),
.B(n_1094),
.C(n_1127),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1071),
.A2(n_1126),
.B(n_1131),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_L g1207 ( 
.A(n_1058),
.B(n_999),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1029),
.A2(n_1045),
.B(n_1142),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1040),
.A2(n_1045),
.B1(n_1087),
.B2(n_1046),
.C(n_1098),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1031),
.B(n_1134),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1055),
.A2(n_1058),
.B1(n_1122),
.B2(n_1124),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1124),
.A2(n_1129),
.B(n_1058),
.Y(n_1212)
);

BUFx4f_ASAP7_75t_L g1213 ( 
.A(n_1032),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1098),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1098),
.B(n_1041),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1046),
.B(n_1035),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1089),
.A2(n_1116),
.B(n_1112),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1069),
.A2(n_1039),
.B(n_681),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1069),
.A2(n_681),
.B(n_1140),
.C(n_1139),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1068),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1139),
.A2(n_681),
.B(n_572),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1146),
.B(n_525),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1139),
.A2(n_681),
.B(n_572),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1070),
.A2(n_674),
.B1(n_675),
.B2(n_657),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1106),
.A2(n_1130),
.A3(n_1132),
.B(n_944),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1068),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1068),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_1143),
.B(n_1016),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_SL g1241 ( 
.A1(n_1139),
.A2(n_1140),
.B(n_1141),
.C(n_940),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1001),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1139),
.A2(n_1141),
.B(n_1140),
.C(n_1069),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1068),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1050),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1139),
.A2(n_681),
.B(n_572),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1143),
.B(n_1016),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_1132),
.A2(n_1115),
.B(n_1112),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1003),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1068),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1139),
.A2(n_681),
.B(n_572),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1081),
.A2(n_1140),
.B(n_1139),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1003),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1001),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1068),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1068),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1001),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1001),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_1026),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1000),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1137),
.A2(n_681),
.B1(n_1140),
.B2(n_1139),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1069),
.A2(n_681),
.B(n_1140),
.C(n_1139),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1139),
.A2(n_681),
.B(n_572),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1132),
.A2(n_1121),
.B(n_1112),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1003),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1106),
.A2(n_1130),
.A3(n_1132),
.B(n_944),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1001),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1065),
.A2(n_1063),
.B1(n_1069),
.B2(n_990),
.C(n_1043),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1069),
.A2(n_681),
.B(n_1140),
.C(n_1139),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1069),
.B(n_983),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1139),
.A2(n_681),
.B(n_572),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1068),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1139),
.A2(n_1140),
.B1(n_1141),
.B2(n_1069),
.Y(n_1286)
);

INVxp67_ASAP7_75t_SL g1287 ( 
.A(n_1001),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1146),
.B(n_675),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1106),
.A2(n_1130),
.A3(n_1132),
.B(n_944),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1144),
.A2(n_924),
.B(n_1112),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1002),
.B(n_825),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1112),
.A2(n_1116),
.B(n_1110),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1220),
.A2(n_1254),
.B1(n_1228),
.B2(n_1232),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1286),
.A2(n_1282),
.B1(n_1225),
.B2(n_1271),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1246),
.A2(n_1284),
.B1(n_1272),
.B2(n_1235),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1158),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1159),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1162),
.A2(n_1283),
.B1(n_1270),
.B2(n_1255),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1255),
.A2(n_1286),
.B1(n_1148),
.B2(n_1157),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1283),
.A2(n_1264),
.B1(n_1280),
.B2(n_1231),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1152),
.A2(n_1149),
.B1(n_1243),
.B2(n_1187),
.Y(n_1301)
);

AOI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1162),
.A2(n_1281),
.B(n_1156),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1153),
.A2(n_1168),
.B1(n_1288),
.B2(n_1160),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1153),
.A2(n_1185),
.B1(n_1155),
.B2(n_1221),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1218),
.A2(n_1247),
.B1(n_1234),
.B2(n_1224),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1151),
.A2(n_1239),
.B1(n_1248),
.B2(n_1222),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1189),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1291),
.Y(n_1309)
);

BUFx2_ASAP7_75t_SL g1310 ( 
.A(n_1267),
.Y(n_1310)
);

CKINVDCx14_ASAP7_75t_R g1311 ( 
.A(n_1213),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1171),
.B(n_1229),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1241),
.B(n_1175),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1191),
.A2(n_1253),
.B1(n_1263),
.B2(n_1237),
.Y(n_1314)
);

INVx8_ASAP7_75t_L g1315 ( 
.A(n_1173),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1238),
.A2(n_1285),
.B1(n_1244),
.B2(n_1260),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1182),
.A2(n_1190),
.B1(n_1265),
.B2(n_1199),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1195),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1180),
.A2(n_1169),
.B(n_1166),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1154),
.Y(n_1320)
);

BUFx4f_ASAP7_75t_SL g1321 ( 
.A(n_1269),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1174),
.A2(n_1165),
.B1(n_1210),
.B2(n_1176),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1200),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1181),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1242),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1287),
.A2(n_1258),
.B1(n_1266),
.B2(n_1163),
.Y(n_1326)
);

INVx2_ASAP7_75t_R g1327 ( 
.A(n_1178),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1216),
.A2(n_1170),
.B1(n_1278),
.B2(n_1172),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1173),
.A2(n_1179),
.B1(n_1215),
.B2(n_1197),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1198),
.A2(n_1281),
.B1(n_1183),
.B2(n_1194),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1203),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1213),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1214),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1196),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1167),
.A2(n_1211),
.B1(n_1252),
.B2(n_1276),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1167),
.A2(n_1257),
.B1(n_1276),
.B2(n_1186),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1257),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1147),
.A2(n_1245),
.B1(n_1193),
.B2(n_1204),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1167),
.A2(n_1202),
.B1(n_1208),
.B2(n_1240),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1201),
.Y(n_1340)
);

CKINVDCx11_ASAP7_75t_R g1341 ( 
.A(n_1188),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1204),
.A2(n_1206),
.B1(n_1251),
.B2(n_1250),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1236),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1207),
.A2(n_1209),
.B1(n_1273),
.B2(n_1227),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1207),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1251),
.A2(n_1249),
.B1(n_1274),
.B2(n_1233),
.Y(n_1346)
);

INVx6_ASAP7_75t_L g1347 ( 
.A(n_1192),
.Y(n_1347)
);

BUFx8_ASAP7_75t_SL g1348 ( 
.A(n_1275),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1217),
.A2(n_1290),
.B1(n_1279),
.B2(n_1261),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1161),
.A2(n_1184),
.B1(n_1219),
.B2(n_1205),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1184),
.A2(n_1219),
.B1(n_1177),
.B2(n_1164),
.Y(n_1351)
);

BUFx8_ASAP7_75t_SL g1352 ( 
.A(n_1184),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1178),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1177),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1277),
.B(n_1289),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1150),
.A2(n_1223),
.B1(n_1230),
.B2(n_1256),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1259),
.A2(n_1262),
.B1(n_1268),
.B2(n_1292),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1220),
.A2(n_878),
.B1(n_1141),
.B2(n_1140),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1151),
.A2(n_1149),
.B1(n_1137),
.B2(n_825),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1267),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1286),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1158),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1220),
.A2(n_878),
.B1(n_1141),
.B2(n_1140),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1154),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1267),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1201),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1154),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1218),
.B(n_1221),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1220),
.A2(n_878),
.B1(n_1141),
.B2(n_1140),
.Y(n_1370)
);

BUFx4_ASAP7_75t_R g1371 ( 
.A(n_1267),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1162),
.A2(n_1283),
.B1(n_347),
.B2(n_350),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1213),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1158),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1267),
.Y(n_1375)
);

BUFx8_ASAP7_75t_L g1376 ( 
.A(n_1203),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1162),
.A2(n_1283),
.B1(n_347),
.B2(n_350),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1201),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1220),
.A2(n_878),
.B1(n_1141),
.B2(n_1140),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1220),
.A2(n_878),
.B1(n_1141),
.B2(n_1140),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1154),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1220),
.A2(n_878),
.B1(n_1141),
.B2(n_1140),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1286),
.A2(n_1137),
.B1(n_681),
.B2(n_1225),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1154),
.Y(n_1384)
);

AOI22x1_ASAP7_75t_SL g1385 ( 
.A1(n_1201),
.A2(n_1034),
.B1(n_825),
.B2(n_246),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1158),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1154),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_R g1388 ( 
.A(n_1148),
.B(n_1062),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1212),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1286),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1158),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1286),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1286),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1162),
.A2(n_1283),
.B1(n_347),
.B2(n_350),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1158),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1212),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1334),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1347),
.A2(n_1352),
.B1(n_1372),
.B2(n_1377),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1348),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1383),
.A2(n_1294),
.B(n_1301),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1347),
.A2(n_1394),
.B1(n_1298),
.B2(n_1354),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1296),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1297),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1396),
.B(n_1389),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1306),
.B(n_1363),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1325),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1389),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1350),
.A2(n_1346),
.B(n_1351),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1305),
.B(n_1369),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1374),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1353),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1395),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1355),
.B(n_1299),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1356),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1358),
.A2(n_1342),
.B(n_1343),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1396),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1323),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1318),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1343),
.A2(n_1350),
.B(n_1351),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1326),
.B(n_1299),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1322),
.A2(n_1330),
.B(n_1293),
.Y(n_1422)
);

AND2x6_ASAP7_75t_L g1423 ( 
.A(n_1347),
.B(n_1338),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1316),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1327),
.B(n_1293),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1319),
.B(n_1315),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1313),
.Y(n_1427)
);

INVx4_ASAP7_75t_SL g1428 ( 
.A(n_1345),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1330),
.A2(n_1307),
.B(n_1314),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1344),
.A2(n_1300),
.B(n_1302),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1314),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_SL g1432 ( 
.A(n_1340),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1324),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1339),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1307),
.A2(n_1370),
.B(n_1382),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1317),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1300),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1360),
.A2(n_1385),
.B1(n_1388),
.B2(n_1312),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1359),
.A2(n_1370),
.B(n_1382),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1384),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1344),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_L g1443 ( 
.A(n_1362),
.B(n_1393),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1336),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1304),
.B(n_1326),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1359),
.B(n_1380),
.C(n_1379),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1295),
.B(n_1392),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1337),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1357),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1349),
.Y(n_1450)
);

AOI21xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1362),
.A2(n_1390),
.B(n_1303),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1390),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1333),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1364),
.B(n_1379),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1335),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1364),
.B(n_1380),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1337),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1295),
.A2(n_1329),
.B(n_1328),
.Y(n_1458)
);

AO21x1_ASAP7_75t_L g1459 ( 
.A1(n_1388),
.A2(n_1373),
.B(n_1332),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1432),
.Y(n_1460)
);

AOI211xp5_ASAP7_75t_L g1461 ( 
.A1(n_1451),
.A2(n_1400),
.B(n_1445),
.C(n_1446),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1440),
.B(n_1368),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1433),
.B(n_1320),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1440),
.B(n_1365),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1451),
.A2(n_1387),
.B(n_1381),
.C(n_1311),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1405),
.B(n_1309),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1406),
.B(n_1310),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1453),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1446),
.A2(n_1311),
.B1(n_1367),
.B2(n_1378),
.C(n_1308),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1371),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1443),
.A2(n_1371),
.B(n_1341),
.C(n_1321),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1441),
.A2(n_1447),
.B1(n_1401),
.B2(n_1454),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1412),
.B(n_1331),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1412),
.B(n_1366),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1406),
.B(n_1375),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1428),
.B(n_1321),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1447),
.A2(n_1361),
.B(n_1376),
.C(n_1437),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1402),
.B(n_1376),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1445),
.A2(n_1456),
.B1(n_1423),
.B2(n_1409),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1399),
.B(n_1414),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1402),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1403),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1430),
.A2(n_1450),
.B(n_1422),
.Y(n_1483)
);

A2O1A1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1439),
.A2(n_1456),
.B(n_1435),
.C(n_1442),
.Y(n_1484)
);

OAI211xp5_ASAP7_75t_L g1485 ( 
.A1(n_1442),
.A2(n_1450),
.B(n_1422),
.C(n_1421),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1427),
.B(n_1459),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1427),
.B(n_1434),
.C(n_1452),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1439),
.A2(n_1435),
.B(n_1421),
.C(n_1429),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1397),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1459),
.B(n_1430),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1410),
.B(n_1413),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1419),
.B(n_1418),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1425),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1425),
.B(n_1438),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1430),
.A2(n_1426),
.B(n_1408),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1426),
.B(n_1411),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1416),
.A2(n_1420),
.B(n_1449),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1407),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1495),
.B(n_1494),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1489),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1481),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1489),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1498),
.B(n_1404),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1495),
.B(n_1408),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1482),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1408),
.Y(n_1508)
);

OAI221xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1461),
.A2(n_1398),
.B1(n_1455),
.B2(n_1444),
.C(n_1431),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_1415),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1490),
.B(n_1458),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1397),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1485),
.A2(n_1458),
.B1(n_1455),
.B2(n_1444),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1493),
.B(n_1408),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1470),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1490),
.B(n_1483),
.Y(n_1516)
);

NOR2xp67_ASAP7_75t_L g1517 ( 
.A(n_1497),
.B(n_1417),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1499),
.B(n_1420),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1471),
.A2(n_1458),
.B1(n_1431),
.B2(n_1424),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1499),
.B(n_1500),
.Y(n_1520)
);

INVxp67_ASAP7_75t_SL g1521 ( 
.A(n_1497),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1484),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1466),
.B(n_1417),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1467),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1484),
.B(n_1458),
.C(n_1436),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1491),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1488),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1488),
.Y(n_1528)
);

AOI222xp33_ASAP7_75t_L g1529 ( 
.A1(n_1519),
.A2(n_1472),
.B1(n_1423),
.B2(n_1485),
.C1(n_1465),
.C2(n_1496),
.Y(n_1529)
);

NAND4xp25_ASAP7_75t_L g1530 ( 
.A(n_1516),
.B(n_1471),
.C(n_1465),
.D(n_1473),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1506),
.B(n_1492),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1514),
.B(n_1520),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1520),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1502),
.Y(n_1534)
);

NOR3xp33_ASAP7_75t_SL g1535 ( 
.A(n_1509),
.B(n_1460),
.C(n_1468),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1512),
.Y(n_1536)
);

OAI211xp5_ASAP7_75t_L g1537 ( 
.A1(n_1516),
.A2(n_1479),
.B(n_1469),
.C(n_1477),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1520),
.Y(n_1538)
);

AOI222xp33_ASAP7_75t_L g1539 ( 
.A1(n_1519),
.A2(n_1423),
.B1(n_1525),
.B2(n_1511),
.C1(n_1522),
.C2(n_1469),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1515),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1504),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1504),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1510),
.B(n_1468),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1506),
.B(n_1487),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1515),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1505),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1526),
.B(n_1511),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1505),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1478),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1505),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1532),
.B(n_1524),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1527),
.B(n_1525),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1550),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1548),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1532),
.B(n_1524),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1534),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1545),
.B(n_1536),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1548),
.B(n_1517),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1548),
.B(n_1517),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1460),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1523),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.B(n_1523),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1545),
.B(n_1512),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1538),
.B(n_1523),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1533),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1538),
.B(n_1550),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1534),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1548),
.B(n_1515),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1544),
.B(n_1475),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1540),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1550),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1503),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1507),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1541),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1542),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1531),
.B(n_1501),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1542),
.Y(n_1585)
);

BUFx2_ASAP7_75t_SL g1586 ( 
.A(n_1548),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1556),
.B(n_1551),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1560),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1582),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1560),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1541),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1572),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1541),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1565),
.B(n_1546),
.Y(n_1596)
);

OAI32xp33_ASAP7_75t_L g1597 ( 
.A1(n_1561),
.A2(n_1530),
.A3(n_1522),
.B1(n_1547),
.B2(n_1549),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1556),
.B(n_1551),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1561),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1556),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1574),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1546),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1556),
.B(n_1530),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1574),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1582),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1577),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1556),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1582),
.B(n_1476),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1578),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1551),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1578),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1564),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1585),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1568),
.B(n_1552),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1555),
.B(n_1527),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1570),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1555),
.B(n_1528),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1568),
.B(n_1552),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1568),
.B(n_1551),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1586),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1587),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1587),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1586),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1605),
.B(n_1611),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1605),
.B(n_1573),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1589),
.B(n_1584),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

OAI322xp33_ASAP7_75t_L g1633 ( 
.A1(n_1600),
.A2(n_1583),
.A3(n_1581),
.B1(n_1549),
.B2(n_1547),
.C1(n_1557),
.C2(n_1569),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1611),
.B(n_1573),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1611),
.B(n_1588),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1588),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1599),
.B(n_1528),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1588),
.B(n_1573),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1591),
.B(n_1620),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1621),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1608),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1592),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1597),
.A2(n_1528),
.B1(n_1521),
.B2(n_1581),
.C(n_1547),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1622),
.B(n_1528),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1598),
.B(n_1559),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1608),
.B(n_1559),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1580),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1621),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1598),
.B(n_1559),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1594),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1597),
.A2(n_1530),
.B(n_1539),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1594),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1615),
.B(n_1553),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1619),
.B(n_1580),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1602),
.B(n_1553),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1601),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1602),
.B(n_1610),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1601),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1603),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1665)
);

OAI32xp33_ASAP7_75t_L g1666 ( 
.A1(n_1638),
.A2(n_1610),
.A3(n_1602),
.B1(n_1628),
.B2(n_1625),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1630),
.Y(n_1667)
);

OR4x1_ASAP7_75t_L g1668 ( 
.A(n_1637),
.B(n_1558),
.C(n_1627),
.D(n_1626),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1664),
.Y(n_1669)
);

XNOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1610),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1654),
.A2(n_1535),
.B1(n_1613),
.B2(n_1628),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1632),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1643),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1643),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1645),
.A2(n_1535),
.B(n_1613),
.C(n_1509),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1632),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1657),
.B(n_1618),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1618),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1636),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1631),
.B(n_1553),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1629),
.A2(n_1539),
.B1(n_1529),
.B2(n_1537),
.C(n_1521),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1629),
.C(n_1641),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1639),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1633),
.A2(n_1613),
.B(n_1539),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1647),
.A2(n_1613),
.B1(n_1551),
.B2(n_1554),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1639),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1644),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1635),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1675),
.A2(n_1637),
.B(n_1634),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1667),
.B(n_1631),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1667),
.B(n_1678),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1669),
.B(n_1649),
.Y(n_1695)
);

O2A1O1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1675),
.A2(n_1663),
.B(n_1644),
.C(n_1661),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1677),
.B(n_1670),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1668),
.Y(n_1698)
);

AOI321xp33_ASAP7_75t_L g1699 ( 
.A1(n_1685),
.A2(n_1662),
.A3(n_1659),
.B1(n_1634),
.B2(n_1640),
.C(n_1651),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1665),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1672),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1682),
.A2(n_1663),
.B(n_1661),
.C(n_1656),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1676),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_SL g1704 ( 
.A1(n_1671),
.A2(n_1656),
.B(n_1653),
.C(n_1558),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1670),
.A2(n_1513),
.B1(n_1529),
.B2(n_1642),
.C(n_1651),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1674),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1679),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1673),
.B(n_1646),
.Y(n_1708)
);

NAND4xp25_ASAP7_75t_SL g1709 ( 
.A(n_1683),
.B(n_1688),
.C(n_1652),
.D(n_1646),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1696),
.A2(n_1666),
.B(n_1684),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1693),
.B(n_1681),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1691),
.B(n_1673),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1692),
.B(n_1648),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1697),
.B(n_1694),
.Y(n_1715)
);

O2A1O1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1698),
.A2(n_1690),
.B(n_1674),
.C(n_1687),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1700),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1705),
.A2(n_1529),
.B1(n_1642),
.B2(n_1660),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1700),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1708),
.B(n_1648),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1706),
.B(n_1652),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1702),
.B(n_1698),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1701),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1715),
.B(n_1706),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1699),
.C(n_1704),
.D(n_1695),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1712),
.B(n_1709),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1717),
.B(n_1690),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1714),
.B(n_1640),
.Y(n_1728)
);

AOI221x1_ASAP7_75t_L g1729 ( 
.A1(n_1722),
.A2(n_1710),
.B1(n_1707),
.B2(n_1703),
.C(n_1689),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1720),
.B(n_1640),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1721),
.B(n_1650),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1711),
.A2(n_1658),
.B1(n_1650),
.B2(n_1655),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_SL g1733 ( 
.A(n_1713),
.B(n_1686),
.C(n_1704),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1717),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1725),
.A2(n_1711),
.B(n_1716),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1732),
.A2(n_1718),
.B1(n_1726),
.B2(n_1668),
.C(n_1733),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_SL g1737 ( 
.A(n_1724),
.B(n_1731),
.Y(n_1737)
);

AOI21xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1727),
.A2(n_1719),
.B(n_1723),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_L g1739 ( 
.A1(n_1729),
.A2(n_1658),
.B(n_1623),
.C(n_1624),
.Y(n_1739)
);

OAI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1735),
.A2(n_1734),
.B1(n_1728),
.B2(n_1730),
.C(n_1660),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1736),
.A2(n_1558),
.B(n_1579),
.C(n_1626),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1738),
.A2(n_1655),
.B1(n_1627),
.B2(n_1609),
.C(n_1617),
.Y(n_1742)
);

AO21x1_ASAP7_75t_L g1743 ( 
.A1(n_1737),
.A2(n_1655),
.B(n_1606),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1549),
.B(n_1617),
.C(n_1616),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1735),
.A2(n_1607),
.B1(n_1616),
.B2(n_1614),
.C(n_1612),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1743),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1740),
.B(n_1603),
.Y(n_1747)
);

OA22x2_ASAP7_75t_L g1748 ( 
.A1(n_1741),
.A2(n_1606),
.B1(n_1614),
.B2(n_1612),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1744),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1745),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1749),
.A2(n_1742),
.B1(n_1563),
.B2(n_1562),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1746),
.B(n_1624),
.Y(n_1752)
);

XOR2xp5_ASAP7_75t_L g1753 ( 
.A(n_1750),
.B(n_1474),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1753),
.Y(n_1754)
);

OAI22x1_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1752),
.B1(n_1747),
.B2(n_1751),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1748),
.B1(n_1609),
.B2(n_1607),
.Y(n_1756)
);

INVxp33_ASAP7_75t_L g1757 ( 
.A(n_1755),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1757),
.A2(n_1576),
.B1(n_1571),
.B2(n_1570),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1756),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1759),
.A2(n_1571),
.B1(n_1570),
.B2(n_1563),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1758),
.A2(n_1571),
.B1(n_1583),
.B2(n_1604),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1595),
.B(n_1593),
.Y(n_1762)
);

AOI21xp33_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1761),
.B(n_1477),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1562),
.B1(n_1563),
.B2(n_1604),
.C(n_1596),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1463),
.B(n_1464),
.C(n_1462),
.Y(n_1766)
);


endmodule