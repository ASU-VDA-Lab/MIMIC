module fake_jpeg_24166_n_307 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_45),
.B1(n_23),
.B2(n_18),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_73),
.B1(n_28),
.B2(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_61),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_18),
.B1(n_25),
.B2(n_23),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_57),
.B(n_63),
.C(n_71),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_38),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_48),
.B(n_41),
.C(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_20),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_21),
.B1(n_32),
.B2(n_20),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_75),
.B(n_36),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_21),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_78),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_21),
.B1(n_32),
.B2(n_35),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_32),
.B1(n_38),
.B2(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_37),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_114),
.B1(n_64),
.B2(n_50),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_19),
.B1(n_28),
.B2(n_30),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_85),
.B(n_108),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_84),
.A2(n_59),
.B1(n_54),
.B2(n_36),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_30),
.B1(n_38),
.B2(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_93),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_26),
.C(n_43),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_116),
.C(n_27),
.Y(n_133)
);

CKINVDCx9p33_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_88),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_91),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

CKINVDCx10_ASAP7_75t_R g144 ( 
.A(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_34),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_99),
.Y(n_134)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_26),
.CON(n_95),
.SN(n_95)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_95),
.A2(n_107),
.B1(n_97),
.B2(n_90),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_103),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_37),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_44),
.B(n_37),
.C(n_33),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_66),
.B1(n_50),
.B2(n_64),
.Y(n_119)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_0),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_57),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_26),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_27),
.B(n_31),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_135),
.B1(n_146),
.B2(n_83),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_16),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_121),
.B(n_133),
.C(n_105),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_51),
.A3(n_44),
.B1(n_54),
.B2(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_108),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_92),
.B1(n_101),
.B2(n_98),
.Y(n_165)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_138),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_81),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_105),
.C(n_88),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_60),
.B1(n_64),
.B2(n_50),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_129),
.A2(n_136),
.B1(n_82),
.B2(n_92),
.Y(n_174)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_132),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_60),
.B1(n_74),
.B2(n_54),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_74),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_74),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_98),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_100),
.B1(n_114),
.B2(n_116),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_181),
.B(n_119),
.Y(n_189)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_157),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_168),
.B1(n_174),
.B2(n_132),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_106),
.B1(n_104),
.B2(n_84),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_165),
.B1(n_172),
.B2(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_81),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_163),
.Y(n_200)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_144),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_160),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_169),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_89),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_87),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_118),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_94),
.B1(n_104),
.B2(n_96),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_104),
.B1(n_99),
.B2(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_145),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_123),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_176),
.B(n_155),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_148),
.C(n_140),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_166),
.B1(n_152),
.B2(n_157),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_134),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_196),
.B(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_137),
.B1(n_147),
.B2(n_134),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_195),
.B1(n_207),
.B2(n_159),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_123),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_122),
.B1(n_136),
.B2(n_131),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_128),
.B(n_124),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_124),
.C(n_138),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_163),
.B(n_178),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_172),
.C(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_205),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_145),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_131),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_121),
.B1(n_117),
.B2(n_113),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_209),
.B1(n_161),
.B2(n_164),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_117),
.B1(n_86),
.B2(n_98),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_97),
.B1(n_90),
.B2(n_58),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_220),
.B1(n_227),
.B2(n_187),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_216),
.A2(n_217),
.B(n_218),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_200),
.B(n_196),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_191),
.B1(n_206),
.B2(n_197),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_175),
.C(n_167),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_184),
.C(n_201),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_224),
.B1(n_186),
.B2(n_204),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_205),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_160),
.B1(n_58),
.B2(n_33),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_160),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_0),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_1),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_201),
.B1(n_202),
.B2(n_33),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_226),
.B1(n_223),
.B2(n_212),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_248),
.B1(n_227),
.B2(n_213),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_193),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_199),
.C(n_188),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_215),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_211),
.C(n_228),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_192),
.C(n_182),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_249),
.B(n_250),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_33),
.C(n_31),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_31),
.C(n_27),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_251),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_216),
.A3(n_218),
.B1(n_226),
.B2(n_222),
.C(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_217),
.B(n_220),
.C(n_214),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_254),
.A2(n_264),
.B1(n_248),
.B2(n_244),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_261),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_R g273 ( 
.A(n_257),
.B(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_231),
.B1(n_230),
.B2(n_229),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_234),
.B(n_239),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_244),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_262),
.B(n_3),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_246),
.C(n_242),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_245),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_261),
.C(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_247),
.C(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.Y(n_287)
);

XNOR2x2_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_250),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_241),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_276),
.B(n_278),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_277),
.A2(n_255),
.B1(n_258),
.B2(n_266),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_266),
.B1(n_264),
.B2(n_257),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_276),
.B(n_279),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_17),
.B(n_14),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_286),
.A2(n_17),
.B(n_14),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_269),
.C(n_275),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_292),
.B(n_293),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_274),
.B(n_279),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_13),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_13),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_13),
.A3(n_12),
.B1(n_5),
.B2(n_6),
.C1(n_2),
.C2(n_8),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_12),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_2),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_299),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_295),
.B(n_12),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_304),
.B(n_6),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_8),
.Y(n_307)
);


endmodule