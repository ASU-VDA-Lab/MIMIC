module fake_jpeg_29579_n_546 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_546);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_61),
.Y(n_125)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_62),
.B(n_64),
.Y(n_133)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_7),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_36),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_72),
.B(n_79),
.Y(n_146)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_83),
.Y(n_149)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_85),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_38),
.B(n_16),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_86),
.Y(n_115)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_90),
.B(n_91),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_37),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_113),
.B(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_64),
.B(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_130),
.Y(n_180)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_82),
.B(n_28),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_99),
.B1(n_102),
.B2(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_140),
.B1(n_160),
.B2(n_60),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_52),
.B1(n_47),
.B2(n_34),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_26),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_86),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_97),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_57),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_159),
.B(n_58),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_95),
.A2(n_51),
.B1(n_52),
.B2(n_34),
.Y(n_160)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_54),
.Y(n_164)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_40),
.B(n_31),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_135),
.B(n_149),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_205),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_176),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_33),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_179),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

INVx6_ASAP7_75t_SL g179 ( 
.A(n_115),
.Y(n_179)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_33),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_186),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_76),
.B1(n_78),
.B2(n_68),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_198),
.B1(n_160),
.B2(n_137),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g242 ( 
.A(n_185),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_45),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_145),
.B1(n_52),
.B2(n_47),
.Y(n_251)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_48),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_209),
.Y(n_231)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

CKINVDCx9p33_ASAP7_75t_R g195 ( 
.A(n_151),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_140),
.A2(n_70),
.B1(n_81),
.B2(n_69),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_118),
.A2(n_101),
.B1(n_96),
.B2(n_51),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_223),
.B1(n_224),
.B2(n_71),
.Y(n_252)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_201),
.B(n_202),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_45),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_133),
.B(n_43),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_215),
.C(n_220),
.Y(n_273)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_127),
.A2(n_51),
.B1(n_40),
.B2(n_20),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_210),
.Y(n_261)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_112),
.A2(n_20),
.B1(n_31),
.B2(n_24),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_219),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_43),
.Y(n_215)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_218),
.B1(n_59),
.B2(n_110),
.Y(n_230)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_217),
.Y(n_265)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_129),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_117),
.B(n_97),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_137),
.A2(n_101),
.B1(n_96),
.B2(n_66),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_167),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_226),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_135),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_227),
.A2(n_258),
.B1(n_187),
.B2(n_216),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_180),
.B(n_154),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_228),
.B(n_264),
.C(n_268),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_236),
.A2(n_23),
.B(n_143),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_171),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_239),
.B(n_12),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_169),
.B(n_223),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_252),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_168),
.A2(n_111),
.B1(n_126),
.B2(n_121),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_251),
.A2(n_253),
.B1(n_59),
.B2(n_79),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_198),
.A2(n_193),
.B1(n_141),
.B2(n_209),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_141),
.B1(n_146),
.B2(n_47),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_146),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_119),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_107),
.C(n_39),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_48),
.C(n_39),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_23),
.C(n_151),
.Y(n_314)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_276),
.A2(n_279),
.B1(n_255),
.B2(n_233),
.Y(n_332)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_237),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_278),
.B(n_288),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_190),
.B1(n_184),
.B2(n_203),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_280),
.A2(n_263),
.B(n_268),
.Y(n_318)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_222),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_294),
.Y(n_337)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

INVx4_ASAP7_75t_SL g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_246),
.A2(n_205),
.B1(n_183),
.B2(n_188),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_287),
.A2(n_242),
.B(n_274),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_231),
.A2(n_79),
.A3(n_199),
.B1(n_44),
.B2(n_26),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_181),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_291),
.B(n_295),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_44),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_292),
.B(n_315),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_224),
.B1(n_23),
.B2(n_37),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_298),
.B(n_240),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_37),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_244),
.B(n_143),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_196),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_303),
.Y(n_338)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_263),
.B(n_231),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

AO22x2_ASAP7_75t_SL g300 ( 
.A1(n_253),
.A2(n_185),
.B1(n_178),
.B2(n_173),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_313),
.B(n_251),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_183),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_302),
.B(n_15),
.Y(n_333)
);

INVx6_ASAP7_75t_SL g303 ( 
.A(n_246),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_229),
.B(n_205),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_273),
.B(n_12),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_23),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_263),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_314),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_231),
.A2(n_236),
.B(n_227),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_228),
.B(n_23),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_257),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_272),
.B1(n_245),
.B2(n_2),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_320),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_324),
.A2(n_353),
.B(n_311),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_296),
.B(n_240),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_342),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_256),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_344),
.C(n_348),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_332),
.A2(n_341),
.B1(n_356),
.B2(n_300),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_333),
.B(n_10),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_313),
.B(n_238),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_339),
.B(n_298),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_276),
.A2(n_243),
.B1(n_255),
.B2(n_267),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_289),
.B(n_259),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_347),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_265),
.C(n_250),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_346),
.A2(n_286),
.B1(n_290),
.B2(n_315),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_242),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_267),
.C(n_254),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_305),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_350),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_292),
.B(n_241),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_351),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_283),
.A2(n_98),
.B(n_87),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_310),
.B1(n_290),
.B2(n_279),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_300),
.A2(n_272),
.B1(n_11),
.B2(n_10),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_0),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_303),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_359),
.B(n_365),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_280),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_361),
.A2(n_368),
.B(n_385),
.Y(n_396)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_281),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_384),
.Y(n_395)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_323),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_374),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_372),
.B(n_382),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_338),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_373),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_319),
.B(n_282),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_277),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_376),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_377),
.A2(n_320),
.B1(n_342),
.B2(n_332),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_300),
.B1(n_310),
.B2(n_317),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_379),
.A2(n_355),
.B1(n_348),
.B2(n_337),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_383),
.Y(n_403)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_322),
.B(n_284),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_285),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_316),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_388),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_331),
.B(n_294),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_344),
.C(n_318),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_328),
.B(n_317),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_322),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_389),
.Y(n_407)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_327),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_327),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_SL g391 ( 
.A(n_324),
.B(n_288),
.C(n_293),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_391),
.A2(n_392),
.B(n_339),
.Y(n_401)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_347),
.A2(n_317),
.B(n_275),
.C(n_297),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_393),
.B(n_424),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_320),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_401),
.B(n_402),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_366),
.B(n_337),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_343),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_417),
.C(n_368),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_377),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_321),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_409),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_382),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_411),
.B(n_421),
.Y(n_443)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_349),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_SL g420 ( 
.A(n_391),
.B(n_357),
.C(n_353),
.Y(n_420)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_380),
.C(n_361),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_358),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_320),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_422),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_371),
.B(n_341),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_407),
.A2(n_346),
.B1(n_363),
.B2(n_373),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_426),
.A2(n_449),
.B(n_419),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_366),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_430),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_429),
.A2(n_399),
.B1(n_400),
.B2(n_414),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_367),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_418),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_358),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_363),
.Y(n_435)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_406),
.B(n_364),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_437),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_388),
.C(n_392),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_452),
.C(n_402),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_390),
.Y(n_440)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_441),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_395),
.A2(n_381),
.B1(n_375),
.B2(n_384),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_445),
.B1(n_448),
.B2(n_334),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_395),
.A2(n_369),
.B1(n_329),
.B2(n_330),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_398),
.A2(n_350),
.B1(n_335),
.B2(n_329),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_398),
.B(n_352),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_450),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_354),
.C(n_336),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_453),
.A2(n_454),
.B1(n_457),
.B2(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_429),
.A2(n_396),
.B1(n_401),
.B2(n_422),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_459),
.C(n_460),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_425),
.A2(n_396),
.B1(n_422),
.B2(n_394),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_425),
.A2(n_394),
.B1(n_393),
.B2(n_420),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_405),
.C(n_414),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_410),
.C(n_419),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_470),
.C(n_474),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_465),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_434),
.A2(n_447),
.B1(n_451),
.B2(n_448),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_435),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_418),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_444),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_427),
.B(n_410),
.C(n_423),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_354),
.C(n_336),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_443),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_477),
.A2(n_471),
.B1(n_473),
.B2(n_456),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_472),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_481),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_434),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_470),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_461),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_466),
.A2(n_447),
.B(n_451),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_490),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_467),
.B(n_446),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_483),
.B(n_487),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_485),
.B(n_460),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_437),
.Y(n_486)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_463),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_491),
.Y(n_494)
);

AND3x1_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_444),
.C(n_440),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_458),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_469),
.Y(n_501)
);

BUFx12_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

INVx11_ASAP7_75t_L g499 ( 
.A(n_493),
.Y(n_499)
);

OA22x2_ASAP7_75t_L g516 ( 
.A1(n_495),
.A2(n_497),
.B1(n_494),
.B2(n_504),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_501),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_476),
.A2(n_487),
.B1(n_489),
.B2(n_477),
.Y(n_500)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

XOR2x2_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_462),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_479),
.B(n_439),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_459),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_335),
.C(n_306),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_488),
.A2(n_475),
.B1(n_455),
.B2(n_456),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_506),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_482),
.A2(n_474),
.B1(n_450),
.B2(n_441),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_495),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_493),
.A2(n_439),
.B1(n_334),
.B2(n_330),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_304),
.B1(n_299),
.B2(n_2),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_508),
.A2(n_493),
.B(n_484),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_510),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_508),
.A2(n_479),
.B(n_484),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_516),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_521),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_503),
.C(n_498),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_512),
.B1(n_522),
.B2(n_6),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_520),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_496),
.B(n_0),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_0),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_L g522 ( 
.A1(n_502),
.A2(n_0),
.B(n_1),
.Y(n_522)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_499),
.C(n_3),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_515),
.B(n_499),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_530),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_527),
.B(n_528),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_501),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_516),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_536),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_525),
.B(n_510),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_523),
.B(n_514),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_539),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_526),
.C(n_516),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_529),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_532),
.C(n_5),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_542),
.A2(n_540),
.B1(n_5),
.B2(n_6),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_1),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_544),
.A2(n_1),
.B(n_5),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_5),
.B(n_6),
.Y(n_546)
);


endmodule