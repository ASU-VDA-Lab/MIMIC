module fake_jpeg_15170_n_24 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_14),
.A2(n_16),
.B1(n_9),
.B2(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_L g16 ( 
.A1(n_9),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_7),
.B(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_17),
.C(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

BUFx24_ASAP7_75t_SL g23 ( 
.A(n_22),
.Y(n_23)
);

BUFx24_ASAP7_75t_SL g24 ( 
.A(n_23),
.Y(n_24)
);


endmodule