module fake_netlist_1_7530_n_1064 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_191, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_1064);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_1064;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_844;
wire n_230;
wire n_209;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_938;
wire n_928;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_1035;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_666;
wire n_621;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_970;
wire n_822;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_899;
wire n_806;
wire n_539;
wire n_1055;
wire n_197;
wire n_201;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_233;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_198;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_12), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_90), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_67), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_96), .Y(n_202) );
BUFx10_ASAP7_75t_L g203 ( .A(n_172), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_85), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_152), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_175), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_86), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_35), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_166), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_169), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_99), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_112), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_58), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_192), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_110), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_22), .B(n_24), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_34), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_50), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_16), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_20), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_142), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_49), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_115), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_62), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_184), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_113), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_87), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_133), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_2), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_165), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_151), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_118), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_5), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_63), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_28), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_194), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_144), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_114), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_157), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_92), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_141), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_138), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_193), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_9), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g251 ( .A(n_187), .B(n_77), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_105), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_33), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_60), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_108), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_93), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_185), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_145), .Y(n_258) );
BUFx8_ASAP7_75t_SL g259 ( .A(n_0), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_28), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_139), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_21), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_98), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_158), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_26), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_181), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_71), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_55), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_67), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_66), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_41), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_140), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_168), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_63), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_109), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_122), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_76), .Y(n_277) );
BUFx10_ASAP7_75t_L g278 ( .A(n_116), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_189), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_146), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_70), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_53), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_120), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_188), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_117), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_72), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_132), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_41), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_190), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_49), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_20), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_126), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_111), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_19), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_186), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_161), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_31), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_7), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_174), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_176), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_167), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_1), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_15), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_82), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_160), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_101), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_51), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_180), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_91), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_24), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_212), .A2(n_75), .B(n_74), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_250), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_250), .B(n_0), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_291), .B(n_1), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_276), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_276), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_276), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_250), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_213), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_276), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_213), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_227), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_227), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
INVx6_ASAP7_75t_L g325 ( .A(n_203), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_212), .A2(n_79), .B(n_78), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_280), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_271), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_280), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_268), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_215), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_215), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_228), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
XNOR2x2_ASAP7_75t_L g337 ( .A(n_208), .B(n_2), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_235), .B(n_3), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_232), .B(n_3), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_237), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_220), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_220), .A2(n_81), .B(n_80), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_271), .B(n_4), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_268), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_282), .B(n_6), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_297), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_225), .A2(n_84), .B(n_83), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_225), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_325), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_313), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_314), .A2(n_286), .B1(n_275), .B2(n_205), .Y(n_355) );
INVx6_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_313), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_316), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_343), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_325), .B(n_266), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_329), .B(n_203), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_341), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_329), .B(n_245), .Y(n_365) );
OA22x2_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_218), .B1(n_219), .B2(n_217), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_341), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
CKINVDCx6p67_ASAP7_75t_R g369 ( .A(n_324), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_325), .B(n_273), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
BUFx8_ASAP7_75t_SL g372 ( .A(n_314), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_325), .B(n_298), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_325), .B(n_298), .Y(n_375) );
INVx8_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_343), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_336), .B(n_206), .Y(n_380) );
INVx5_ASAP7_75t_L g381 ( .A(n_333), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_343), .A2(n_239), .B1(n_254), .B2(n_221), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_326), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_312), .B(n_277), .Y(n_385) );
OAI22xp33_ASAP7_75t_SL g386 ( .A1(n_340), .A2(n_265), .B1(n_267), .B2(n_260), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_333), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_333), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_333), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_311), .B(n_197), .C(n_195), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_338), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_345), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g393 ( .A(n_333), .B(n_202), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_327), .A2(n_200), .B(n_198), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_365), .B(n_338), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_365), .B(n_339), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_370), .B(n_339), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_356), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_391), .B(n_345), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_275), .B1(n_295), .B2(n_205), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_345), .B1(n_318), .B2(n_337), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_361), .B(n_373), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_369), .B(n_196), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_356), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_375), .B(n_318), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_380), .B(n_206), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_362), .B(n_295), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_369), .B(n_199), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_384), .B(n_319), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_356), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_384), .B(n_319), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_376), .B(n_207), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_355), .B(n_337), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_376), .B(n_209), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_392), .B(n_210), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_392), .B(n_382), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_354), .B(n_321), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g418 ( .A(n_386), .B(n_259), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_357), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_354), .B(n_321), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_360), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_364), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_358), .B(n_201), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_385), .B(n_358), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_360), .B(n_279), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_360), .B(n_204), .Y(n_426) );
NOR2x1p5_ASAP7_75t_L g427 ( .A(n_372), .B(n_259), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_379), .B(n_279), .Y(n_428) );
BUFx8_ASAP7_75t_L g429 ( .A(n_351), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_364), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_379), .A2(n_342), .B(n_347), .C(n_327), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_367), .B(n_293), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_390), .B(n_322), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_368), .B(n_293), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_355), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_368), .B(n_296), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_377), .B(n_296), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_366), .A2(n_302), .B1(n_288), .B2(n_274), .C(n_238), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_378), .A2(n_322), .B1(n_332), .B2(n_323), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_394), .A2(n_342), .B(n_327), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_378), .A2(n_253), .B1(n_262), .B2(n_233), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_394), .B(n_300), .Y(n_443) );
BUFx8_ASAP7_75t_L g444 ( .A(n_386), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_389), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_394), .B(n_245), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_389), .B(n_323), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_381), .A2(n_224), .B1(n_270), .B2(n_269), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_393), .B(n_332), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_381), .B(n_344), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_381), .B(n_346), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_349), .A2(n_224), .B1(n_270), .B2(n_269), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_350), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_350), .A2(n_303), .B1(n_310), .B2(n_216), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_352), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_352), .A2(n_290), .B1(n_307), .B2(n_281), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_352), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_353), .B(n_285), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_353), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_371), .B(n_230), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_371), .A2(n_290), .B1(n_307), .B2(n_281), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_459), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_433), .A2(n_342), .B(n_347), .C(n_282), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_399), .B(n_297), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_464), .B(n_7), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_441), .A2(n_347), .B(n_311), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_396), .B(n_203), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_403), .B(n_278), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_431), .A2(n_214), .B(n_211), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_395), .B(n_278), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_431), .A2(n_445), .B(n_447), .C(n_443), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_426), .A2(n_223), .B(n_222), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_402), .B(n_234), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_433), .A2(n_229), .B(n_231), .C(n_226), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_412), .B(n_236), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_409), .A2(n_242), .B(n_246), .C(n_241), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_424), .B(n_243), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_435), .A2(n_248), .B1(n_257), .B2(n_255), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_439), .A2(n_249), .B(n_252), .C(n_247), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_426), .A2(n_423), .B(n_405), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_407), .B(n_272), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_408), .B(n_8), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_423), .A2(n_263), .B(n_256), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_450), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_416), .B(n_258), .Y(n_490) );
INVx11_ASAP7_75t_L g491 ( .A(n_429), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_415), .B(n_261), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_406), .B(n_264), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_409), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_411), .B(n_283), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_411), .B(n_284), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_427), .B(n_251), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_400), .A2(n_289), .B(n_292), .C(n_287), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_419), .A2(n_301), .B(n_299), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_425), .A2(n_306), .B(n_305), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_428), .A2(n_309), .B(n_244), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_414), .B(n_304), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_422), .A2(n_244), .B(n_240), .Y(n_503) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_446), .A2(n_383), .B(n_374), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_398), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_432), .A2(n_436), .B(n_434), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_429), .B(n_228), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_437), .B(n_308), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_404), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_442), .A2(n_418), .B(n_420), .C(n_417), .Y(n_510) );
OR2x6_ASAP7_75t_L g511 ( .A(n_455), .B(n_334), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_452), .A2(n_317), .B(n_320), .C(n_315), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_410), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_453), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_452), .A2(n_317), .B(n_320), .C(n_315), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_440), .A2(n_457), .B1(n_449), .B2(n_448), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_440), .B(n_8), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_461), .A2(n_331), .B(n_330), .C(n_328), .Y(n_518) );
OR2x6_ASAP7_75t_L g519 ( .A(n_444), .B(n_335), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_454), .B(n_9), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_438), .A2(n_331), .B(n_330), .C(n_328), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_463), .A2(n_328), .B1(n_330), .B2(n_331), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_451), .B(n_10), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_456), .B(n_10), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_458), .B(n_11), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_460), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_462), .B(n_13), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_401), .A2(n_14), .B1(n_17), .B2(n_18), .Y(n_528) );
CKINVDCx8_ASAP7_75t_R g529 ( .A(n_407), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_430), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_401), .A2(n_363), .B1(n_359), .B2(n_19), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_396), .B(n_17), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_401), .A2(n_363), .B1(n_21), .B2(n_22), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_399), .A2(n_363), .B1(n_23), .B2(n_25), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_396), .B(n_18), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_396), .B(n_23), .Y(n_536) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_459), .Y(n_537) );
NOR2xp33_ASAP7_75t_R g538 ( .A(n_435), .B(n_25), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_401), .A2(n_26), .B1(n_27), .B2(n_29), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_396), .B(n_27), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_399), .B(n_29), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_399), .A2(n_363), .B1(n_31), .B2(n_32), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_433), .A2(n_363), .B(n_32), .C(n_33), .Y(n_543) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_441), .A2(n_30), .B(n_34), .Y(n_544) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_397), .A2(n_363), .B(n_30), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_413), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_459), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_403), .B(n_36), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_399), .A2(n_39), .B1(n_40), .B2(n_42), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_433), .A2(n_39), .B(n_40), .C(n_42), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_401), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_403), .B(n_43), .Y(n_552) );
INVx4_ASAP7_75t_L g553 ( .A(n_430), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_429), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_429), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_441), .A2(n_89), .B(n_88), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_396), .B(n_44), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_399), .B(n_45), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_396), .B(n_46), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_412), .B(n_46), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_396), .B(n_47), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_430), .Y(n_562) );
NOR2x1_ASAP7_75t_SL g563 ( .A(n_519), .B(n_47), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_535), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_494), .B(n_48), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_491), .Y(n_566) );
BUFx3_ASAP7_75t_L g567 ( .A(n_554), .Y(n_567) );
BUFx10_ASAP7_75t_L g568 ( .A(n_555), .Y(n_568) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_466), .A2(n_48), .A3(n_50), .B(n_51), .Y(n_569) );
OR2x6_ASAP7_75t_L g570 ( .A(n_507), .B(n_52), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_536), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_547), .B(n_54), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_489), .B(n_54), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_541), .B(n_56), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_540), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_541), .B(n_56), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_558), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_511), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_558), .B(n_57), .Y(n_579) );
AOI221x1_ASAP7_75t_L g580 ( .A1(n_545), .A2(n_58), .B1(n_59), .B2(n_60), .C(n_61), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_537), .A2(n_59), .B1(n_61), .B2(n_62), .Y(n_581) );
NAND3x1_ASAP7_75t_L g582 ( .A(n_549), .B(n_64), .C(n_65), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_532), .B(n_64), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_531), .A2(n_65), .B1(n_66), .B2(n_68), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_559), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_471), .B(n_68), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_557), .B(n_69), .Y(n_587) );
AO31x2_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_72), .A3(n_73), .B(n_94), .Y(n_588) );
INVx3_ASAP7_75t_SL g589 ( .A(n_497), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_487), .B(n_548), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_561), .B(n_73), .Y(n_591) );
NOR2x1_ASAP7_75t_SL g592 ( .A(n_519), .B(n_95), .Y(n_592) );
AO32x2_ASAP7_75t_L g593 ( .A1(n_528), .A2(n_97), .A3(n_100), .B1(n_102), .B2(n_103), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_486), .A2(n_104), .B1(n_106), .B2(n_107), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_511), .A2(n_119), .B1(n_121), .B2(n_123), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_467), .B(n_124), .Y(n_596) );
AO32x2_ASAP7_75t_L g597 ( .A1(n_539), .A2(n_125), .A3(n_127), .B1(n_128), .B2(n_129), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_552), .B(n_130), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_553), .Y(n_599) );
AO21x2_ASAP7_75t_L g600 ( .A1(n_556), .A2(n_135), .B(n_136), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_529), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_467), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_538), .B(n_143), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_511), .Y(n_605) );
BUFx3_ASAP7_75t_L g606 ( .A(n_527), .Y(n_606) );
AO31x2_ASAP7_75t_L g607 ( .A1(n_543), .A2(n_148), .A3(n_149), .B(n_150), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_479), .A2(n_153), .B(n_154), .C(n_155), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_470), .B(n_156), .Y(n_609) );
OAI21x1_ASAP7_75t_SL g610 ( .A1(n_553), .A2(n_159), .B(n_163), .Y(n_610) );
INVx3_ASAP7_75t_L g611 ( .A(n_562), .Y(n_611) );
NOR4xp25_ASAP7_75t_L g612 ( .A(n_546), .B(n_177), .C(n_178), .D(n_179), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_516), .A2(n_182), .B(n_183), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_498), .B(n_484), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_520), .Y(n_615) );
AO31x2_ASAP7_75t_L g616 ( .A1(n_518), .A2(n_515), .A3(n_512), .B(n_481), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_508), .A2(n_500), .B(n_478), .Y(n_617) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_550), .A2(n_521), .A3(n_551), .B(n_523), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_495), .A2(n_496), .B(n_493), .Y(n_619) );
BUFx3_ASAP7_75t_L g620 ( .A(n_497), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_482), .A2(n_492), .B(n_501), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_475), .A2(n_468), .B1(n_517), .B2(n_483), .C(n_503), .Y(n_622) );
NOR2xp67_ASAP7_75t_SL g623 ( .A(n_562), .B(n_514), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_490), .A2(n_502), .B(n_480), .Y(n_624) );
OA22x2_ASAP7_75t_L g625 ( .A1(n_533), .A2(n_497), .B1(n_542), .B2(n_534), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_513), .Y(n_626) );
AO31x2_ASAP7_75t_L g627 ( .A1(n_525), .A2(n_526), .A3(n_524), .B(n_522), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_472), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_520), .B(n_560), .Y(n_629) );
AO31x2_ASAP7_75t_L g630 ( .A1(n_488), .A2(n_477), .A3(n_499), .B(n_509), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_505), .Y(n_631) );
AO31x2_ASAP7_75t_L g632 ( .A1(n_466), .A2(n_474), .A3(n_544), .B(n_431), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_494), .B(n_396), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_476), .A2(n_506), .B(n_469), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_473), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_529), .B(n_435), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_535), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_494), .B(n_396), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_535), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_547), .A2(n_391), .B1(n_537), .B2(n_465), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_553), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_535), .Y(n_642) );
AO31x2_ASAP7_75t_L g643 ( .A1(n_466), .A2(n_474), .A3(n_544), .B(n_431), .Y(n_643) );
INVx4_ASAP7_75t_L g644 ( .A(n_491), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_473), .Y(n_645) );
OA21x2_ASAP7_75t_L g646 ( .A1(n_469), .A2(n_466), .B(n_441), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_494), .B(n_396), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_494), .B(n_396), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_529), .B(n_435), .Y(n_649) );
AO31x2_ASAP7_75t_L g650 ( .A1(n_466), .A2(n_474), .A3(n_544), .B(n_431), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_474), .A2(n_445), .B(n_485), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_489), .B(n_391), .Y(n_652) );
BUFx6f_ASAP7_75t_SL g653 ( .A(n_554), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_494), .B(n_396), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_494), .B(n_396), .Y(n_655) );
OA21x2_ASAP7_75t_L g656 ( .A1(n_469), .A2(n_466), .B(n_441), .Y(n_656) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_469), .A2(n_466), .B(n_441), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_535), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_494), .B(n_396), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_474), .A2(n_445), .B(n_485), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_489), .B(n_459), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_476), .A2(n_506), .B(n_469), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_476), .A2(n_506), .B(n_469), .Y(n_663) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_469), .A2(n_504), .B(n_441), .Y(n_664) );
AO31x2_ASAP7_75t_L g665 ( .A1(n_466), .A2(n_474), .A3(n_544), .B(n_431), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_469), .A2(n_504), .B(n_441), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_476), .A2(n_506), .B(n_469), .Y(n_667) );
AO31x2_ASAP7_75t_L g668 ( .A1(n_466), .A2(n_474), .A3(n_544), .B(n_431), .Y(n_668) );
INVx5_ASAP7_75t_L g669 ( .A(n_519), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_633), .B(n_638), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_570), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_634), .A2(n_663), .B(n_662), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_647), .B(n_648), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_574), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_615), .Y(n_675) );
AO21x2_ASAP7_75t_L g676 ( .A1(n_613), .A2(n_666), .B(n_664), .Y(n_676) );
NOR2x1_ASAP7_75t_R g677 ( .A(n_644), .B(n_669), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_574), .A2(n_625), .B1(n_598), .B2(n_622), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_652), .A2(n_636), .B1(n_649), .B2(n_640), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_654), .B(n_655), .Y(n_680) );
OA21x2_ASAP7_75t_L g681 ( .A1(n_651), .A2(n_660), .B(n_580), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_626), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_565), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_659), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_661), .B(n_577), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_602), .Y(n_686) );
CKINVDCx6p67_ASAP7_75t_R g687 ( .A(n_644), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_646), .A2(n_656), .B(n_657), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_669), .B(n_623), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_635), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_614), .B(n_564), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_669), .Y(n_692) );
AO21x2_ASAP7_75t_L g693 ( .A1(n_600), .A2(n_612), .B(n_610), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_571), .A2(n_639), .B(n_658), .C(n_575), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_645), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_590), .B(n_585), .Y(n_696) );
OAI21x1_ASAP7_75t_SL g697 ( .A1(n_592), .A2(n_563), .B(n_595), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_637), .B(n_642), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_581), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_570), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_572), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_629), .B(n_586), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_573), .A2(n_582), .B1(n_579), .B2(n_576), .Y(n_703) );
AO31x2_ASAP7_75t_L g704 ( .A1(n_584), .A2(n_592), .A3(n_563), .B(n_668), .Y(n_704) );
AO21x2_ASAP7_75t_L g705 ( .A1(n_583), .A2(n_591), .B(n_587), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_608), .A2(n_599), .B(n_641), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_624), .A2(n_598), .B(n_609), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_606), .Y(n_708) );
INVx6_ASAP7_75t_L g709 ( .A(n_568), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_628), .A2(n_596), .B(n_631), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_594), .A2(n_605), .B(n_578), .Y(n_711) );
AO31x2_ASAP7_75t_L g712 ( .A1(n_632), .A2(n_668), .A3(n_665), .B(n_650), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_603), .B(n_601), .Y(n_713) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_611), .A2(n_668), .B(n_665), .Y(n_714) );
BUFx3_ASAP7_75t_L g715 ( .A(n_568), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_569), .Y(n_716) );
INVx6_ASAP7_75t_L g717 ( .A(n_567), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_618), .B(n_665), .Y(n_718) );
OAI21x1_ASAP7_75t_L g719 ( .A1(n_632), .A2(n_643), .B(n_650), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_604), .A2(n_632), .B(n_650), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g721 ( .A(n_604), .B(n_620), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_566), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_569), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_630), .B(n_627), .Y(n_724) );
INVx1_ASAP7_75t_SL g725 ( .A(n_589), .Y(n_725) );
AO31x2_ASAP7_75t_L g726 ( .A1(n_643), .A2(n_607), .A3(n_588), .B(n_597), .Y(n_726) );
OAI21x1_ASAP7_75t_L g727 ( .A1(n_607), .A2(n_593), .B(n_597), .Y(n_727) );
BUFx3_ASAP7_75t_L g728 ( .A(n_653), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_618), .B(n_627), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_630), .B(n_627), .Y(n_730) );
OA21x2_ASAP7_75t_L g731 ( .A1(n_607), .A2(n_588), .B(n_593), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_616), .B(n_653), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_616), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_597), .B(n_613), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_626), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_633), .B(n_638), .Y(n_736) );
INVx2_ASAP7_75t_SL g737 ( .A(n_568), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_633), .B(n_638), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_633), .B(n_638), .Y(n_739) );
AND2x4_ASAP7_75t_L g740 ( .A(n_606), .B(n_599), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_652), .B(n_391), .Y(n_741) );
BUFx3_ASAP7_75t_L g742 ( .A(n_644), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_633), .B(n_638), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_633), .B(n_638), .Y(n_744) );
AO31x2_ASAP7_75t_L g745 ( .A1(n_634), .A2(n_662), .A3(n_667), .B(n_663), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g746 ( .A(n_669), .B(n_623), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_634), .A2(n_663), .B(n_662), .Y(n_747) );
BUFx12f_ASAP7_75t_L g748 ( .A(n_644), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_652), .B(n_391), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_626), .Y(n_750) );
OAI21x1_ASAP7_75t_SL g751 ( .A1(n_592), .A2(n_563), .B(n_613), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_606), .B(n_599), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_633), .B(n_638), .Y(n_753) );
AO31x2_ASAP7_75t_L g754 ( .A1(n_634), .A2(n_662), .A3(n_667), .B(n_663), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_626), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_669), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_634), .A2(n_663), .B(n_662), .Y(n_757) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_574), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_626), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_626), .Y(n_760) );
INVxp67_ASAP7_75t_L g761 ( .A(n_574), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g762 ( .A1(n_619), .A2(n_617), .B(n_621), .C(n_510), .Y(n_762) );
BUFx2_ASAP7_75t_L g763 ( .A(n_570), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_626), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_633), .B(n_638), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_626), .Y(n_766) );
OA21x2_ASAP7_75t_L g767 ( .A1(n_634), .A2(n_663), .B(n_662), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_626), .Y(n_768) );
BUFx3_ASAP7_75t_L g769 ( .A(n_709), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_680), .B(n_670), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_682), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_670), .B(n_673), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_735), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_750), .Y(n_774) );
INVx4_ASAP7_75t_L g775 ( .A(n_689), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_767), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_755), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_759), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_760), .Y(n_779) );
OR2x2_ASAP7_75t_L g780 ( .A(n_673), .B(n_736), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_724), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_736), .B(n_738), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_738), .B(n_739), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_764), .Y(n_784) );
OA21x2_ASAP7_75t_L g785 ( .A1(n_727), .A2(n_747), .B(n_672), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_724), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_766), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_730), .Y(n_788) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_684), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_768), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_698), .Y(n_791) );
OA21x2_ASAP7_75t_L g792 ( .A1(n_672), .A2(n_757), .B(n_747), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_695), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_690), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_739), .B(n_743), .Y(n_795) );
OR2x6_ASAP7_75t_L g796 ( .A(n_678), .B(n_689), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_743), .Y(n_797) );
BUFx4f_ASAP7_75t_L g798 ( .A(n_687), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_723), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_744), .B(n_753), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_744), .B(n_753), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_765), .Y(n_802) );
INVx4_ASAP7_75t_L g803 ( .A(n_746), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_765), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_686), .Y(n_805) );
OR2x6_ASAP7_75t_L g806 ( .A(n_678), .B(n_746), .Y(n_806) );
BUFx3_ASAP7_75t_L g807 ( .A(n_709), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g808 ( .A1(n_694), .A2(n_707), .B(n_710), .Y(n_808) );
AO21x2_ASAP7_75t_L g809 ( .A1(n_762), .A2(n_734), .B(n_688), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_758), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_709), .Y(n_811) );
CKINVDCx11_ASAP7_75t_R g812 ( .A(n_748), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_717), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_694), .B(n_756), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_732), .B(n_712), .Y(n_815) );
OR2x6_ASAP7_75t_L g816 ( .A(n_674), .B(n_697), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_685), .Y(n_817) );
INVx4_ASAP7_75t_SL g818 ( .A(n_704), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_745), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_696), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_692), .Y(n_821) );
INVx3_ASAP7_75t_L g822 ( .A(n_740), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_691), .Y(n_823) );
BUFx2_ASAP7_75t_L g824 ( .A(n_692), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_671), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_712), .B(n_691), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_761), .Y(n_827) );
INVx3_ASAP7_75t_L g828 ( .A(n_740), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_754), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_679), .B(n_703), .C(n_707), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_701), .B(n_683), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_761), .Y(n_832) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_700), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_752), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_754), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_675), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_675), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_729), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_716), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_772), .B(n_714), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_772), .B(n_719), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_826), .B(n_718), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_799), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_782), .B(n_712), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_776), .Y(n_845) );
AND2x4_ASAP7_75t_L g846 ( .A(n_781), .B(n_720), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_821), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_782), .B(n_712), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_783), .B(n_733), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_830), .A2(n_702), .B1(n_763), .B2(n_699), .C(n_749), .Y(n_850) );
OR2x2_ASAP7_75t_L g851 ( .A(n_826), .B(n_718), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_783), .B(n_702), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_800), .B(n_741), .Y(n_853) );
OR2x2_ASAP7_75t_L g854 ( .A(n_770), .B(n_726), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_800), .B(n_713), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_801), .B(n_725), .Y(n_856) );
AND2x4_ASAP7_75t_SL g857 ( .A(n_775), .B(n_737), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_801), .B(n_726), .Y(n_858) );
INVxp67_ASAP7_75t_L g859 ( .A(n_789), .Y(n_859) );
INVx8_ASAP7_75t_L g860 ( .A(n_796), .Y(n_860) );
BUFx2_ASAP7_75t_L g861 ( .A(n_810), .Y(n_861) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_810), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_780), .B(n_725), .Y(n_863) );
OAI222xp33_ASAP7_75t_L g864 ( .A1(n_796), .A2(n_721), .B1(n_722), .B2(n_708), .C1(n_728), .C2(n_715), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_795), .B(n_705), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_796), .A2(n_705), .B1(n_711), .B2(n_751), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_793), .B(n_731), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_824), .Y(n_868) );
INVx2_ASAP7_75t_SL g869 ( .A(n_775), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_793), .B(n_731), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_786), .B(n_681), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_795), .B(n_721), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_788), .B(n_704), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_815), .B(n_754), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_824), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_802), .B(n_717), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_804), .B(n_717), .Y(n_877) );
BUFx2_ASAP7_75t_L g878 ( .A(n_816), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_797), .B(n_711), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_838), .B(n_676), .Y(n_880) );
AND2x4_ASAP7_75t_L g881 ( .A(n_818), .B(n_706), .Y(n_881) );
INVx1_ASAP7_75t_SL g882 ( .A(n_812), .Y(n_882) );
BUFx3_ASAP7_75t_L g883 ( .A(n_775), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_820), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_794), .B(n_693), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_791), .B(n_677), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_845), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_843), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_843), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_844), .B(n_792), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_844), .B(n_792), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_848), .B(n_792), .Y(n_892) );
BUFx2_ASAP7_75t_L g893 ( .A(n_847), .Y(n_893) );
OR2x2_ASAP7_75t_L g894 ( .A(n_865), .B(n_815), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_868), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_848), .B(n_785), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_884), .B(n_817), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_841), .B(n_785), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_849), .B(n_831), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_840), .B(n_819), .Y(n_900) );
INVxp67_ASAP7_75t_L g901 ( .A(n_853), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_849), .B(n_831), .Y(n_902) );
AND2x4_ASAP7_75t_L g903 ( .A(n_846), .B(n_818), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_852), .B(n_823), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_842), .B(n_819), .Y(n_905) );
AND2x4_ASAP7_75t_L g906 ( .A(n_846), .B(n_818), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_879), .B(n_771), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_840), .B(n_829), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_858), .B(n_835), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_882), .B(n_722), .Y(n_910) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_875), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_858), .B(n_839), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_859), .B(n_863), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_856), .B(n_812), .Y(n_914) );
BUFx3_ASAP7_75t_L g915 ( .A(n_883), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_867), .B(n_809), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_870), .B(n_809), .Y(n_917) );
AND2x2_ASAP7_75t_SL g918 ( .A(n_878), .B(n_814), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_855), .B(n_773), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_872), .B(n_774), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_888), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_903), .B(n_818), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_887), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_894), .B(n_874), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_888), .Y(n_925) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_895), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_889), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_890), .B(n_885), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_891), .B(n_885), .Y(n_929) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_911), .Y(n_930) );
OR2x2_ASAP7_75t_L g931 ( .A(n_894), .B(n_874), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_891), .B(n_851), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_892), .B(n_873), .Y(n_933) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_893), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_892), .B(n_873), .Y(n_935) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_893), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_915), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_896), .B(n_870), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_896), .B(n_880), .Y(n_939) );
OR2x6_ASAP7_75t_L g940 ( .A(n_915), .B(n_860), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_898), .B(n_880), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_898), .B(n_871), .Y(n_942) );
OR2x2_ASAP7_75t_L g943 ( .A(n_909), .B(n_854), .Y(n_943) );
INVx3_ASAP7_75t_L g944 ( .A(n_903), .Y(n_944) );
OR2x2_ASAP7_75t_L g945 ( .A(n_909), .B(n_854), .Y(n_945) );
AND2x4_ASAP7_75t_L g946 ( .A(n_903), .B(n_881), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_905), .B(n_861), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_915), .Y(n_948) );
NOR2x1p5_ASAP7_75t_L g949 ( .A(n_906), .B(n_883), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_938), .B(n_916), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_926), .B(n_897), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_938), .B(n_916), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_928), .B(n_917), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_949), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_921), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_921), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_923), .Y(n_957) );
OAI21xp33_ASAP7_75t_L g958 ( .A1(n_930), .A2(n_913), .B(n_901), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_932), .B(n_917), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_928), .B(n_899), .Y(n_960) );
INVxp67_ASAP7_75t_L g961 ( .A(n_937), .Y(n_961) );
INVx3_ASAP7_75t_L g962 ( .A(n_940), .Y(n_962) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_934), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_929), .B(n_902), .Y(n_964) );
AOI21xp33_ASAP7_75t_SL g965 ( .A1(n_940), .A2(n_914), .B(n_910), .Y(n_965) );
NOR2x1_ASAP7_75t_L g966 ( .A(n_949), .B(n_883), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_940), .A2(n_850), .B1(n_918), .B2(n_886), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_925), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_941), .B(n_929), .Y(n_969) );
AOI21xp5_ASAP7_75t_SL g970 ( .A1(n_940), .A2(n_869), .B(n_862), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_925), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_941), .B(n_900), .Y(n_972) );
INVx1_ASAP7_75t_SL g973 ( .A(n_948), .Y(n_973) );
INVx3_ASAP7_75t_L g974 ( .A(n_940), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_932), .B(n_905), .Y(n_975) );
NOR2x1_ASAP7_75t_L g976 ( .A(n_944), .B(n_864), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_939), .B(n_907), .Y(n_977) );
NOR2xp33_ASAP7_75t_SL g978 ( .A(n_922), .B(n_798), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_927), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_939), .B(n_912), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_942), .B(n_908), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_975), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_955), .B(n_933), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_975), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_955), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_956), .B(n_933), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_957), .Y(n_987) );
NAND2x1p5_ASAP7_75t_L g988 ( .A(n_966), .B(n_798), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_956), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_959), .B(n_924), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_971), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_971), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_950), .B(n_935), .Y(n_993) );
OAI33xp33_ASAP7_75t_L g994 ( .A1(n_951), .A2(n_919), .A3(n_924), .B1(n_931), .B2(n_920), .B3(n_904), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_967), .A2(n_931), .B1(n_918), .B2(n_944), .Y(n_995) );
OR2x2_ASAP7_75t_L g996 ( .A(n_959), .B(n_943), .Y(n_996) );
NOR2xp67_ASAP7_75t_L g997 ( .A(n_962), .B(n_944), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_979), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_979), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_953), .B(n_943), .Y(n_1000) );
AOI21xp33_ASAP7_75t_SL g1001 ( .A1(n_954), .A2(n_860), .B(n_944), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_950), .B(n_935), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_968), .B(n_942), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_983), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_983), .Y(n_1005) );
O2A1O1Ixp5_ASAP7_75t_L g1006 ( .A1(n_994), .A2(n_962), .B(n_974), .C(n_977), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_988), .A2(n_962), .B1(n_974), .B2(n_954), .Y(n_1007) );
OAI21xp5_ASAP7_75t_L g1008 ( .A1(n_988), .A2(n_976), .B(n_970), .Y(n_1008) );
A2O1A1Ixp33_ASAP7_75t_L g1009 ( .A1(n_997), .A2(n_965), .B(n_958), .C(n_1001), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_995), .A2(n_974), .B1(n_970), .B2(n_978), .C(n_961), .Y(n_1010) );
OAI22xp33_ASAP7_75t_SL g1011 ( .A1(n_995), .A2(n_973), .B1(n_963), .B2(n_869), .Y(n_1011) );
OAI322xp33_ASAP7_75t_L g1012 ( .A1(n_990), .A2(n_960), .A3(n_964), .B1(n_980), .B2(n_945), .C1(n_947), .C2(n_936), .Y(n_1012) );
OAI222xp33_ASAP7_75t_L g1013 ( .A1(n_996), .A2(n_969), .B1(n_806), .B2(n_981), .C1(n_947), .C2(n_972), .Y(n_1013) );
OAI21xp5_ASAP7_75t_L g1014 ( .A1(n_986), .A2(n_798), .B(n_969), .Y(n_1014) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_986), .A2(n_981), .B(n_866), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1003), .Y(n_1016) );
OAI22xp5_ASAP7_75t_SL g1017 ( .A1(n_982), .A2(n_918), .B1(n_806), .B2(n_803), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_1003), .A2(n_857), .B(n_946), .Y(n_1018) );
AOI21xp5_ASAP7_75t_L g1019 ( .A1(n_1009), .A2(n_857), .B(n_984), .Y(n_1019) );
OAI21xp33_ASAP7_75t_L g1020 ( .A1(n_1011), .A2(n_989), .B(n_985), .Y(n_1020) );
OAI21xp33_ASAP7_75t_L g1021 ( .A1(n_1010), .A2(n_992), .B(n_991), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_1018), .A2(n_1000), .B1(n_1002), .B2(n_993), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_1012), .B(n_998), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_1008), .A2(n_860), .B1(n_945), .B2(n_878), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1016), .B(n_952), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1004), .B(n_952), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1005), .B(n_999), .Y(n_1027) );
NOR3xp33_ASAP7_75t_L g1028 ( .A(n_1006), .B(n_833), .C(n_825), .Y(n_1028) );
OAI222xp33_ASAP7_75t_L g1029 ( .A1(n_1022), .A2(n_1023), .B1(n_1019), .B2(n_1024), .C1(n_1007), .C2(n_1025), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1028), .B(n_1015), .Y(n_1030) );
NOR3xp33_ASAP7_75t_SL g1031 ( .A(n_1021), .B(n_1013), .C(n_1017), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_1027), .Y(n_1032) );
NOR3xp33_ASAP7_75t_L g1033 ( .A(n_1020), .B(n_1013), .C(n_1014), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1026), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_1019), .A2(n_857), .B(n_811), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1032), .Y(n_1036) );
OAI211xp5_ASAP7_75t_SL g1037 ( .A1(n_1031), .A2(n_876), .B(n_877), .C(n_813), .Y(n_1037) );
OAI21xp33_ASAP7_75t_L g1038 ( .A1(n_1030), .A2(n_987), .B(n_972), .Y(n_1038) );
OAI221xp5_ASAP7_75t_SL g1039 ( .A1(n_1033), .A2(n_806), .B1(n_816), .B2(n_807), .C(n_769), .Y(n_1039) );
NAND3xp33_ASAP7_75t_SL g1040 ( .A(n_1035), .B(n_803), .C(n_808), .Y(n_1040) );
AND2x4_ASAP7_75t_SL g1041 ( .A(n_1036), .B(n_1034), .Y(n_1041) );
NOR3xp33_ASAP7_75t_L g1042 ( .A(n_1037), .B(n_1029), .C(n_742), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1038), .Y(n_1043) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1039), .Y(n_1044) );
NOR2x1_ASAP7_75t_L g1045 ( .A(n_1044), .B(n_1040), .Y(n_1045) );
AOI31xp33_ASAP7_75t_L g1046 ( .A1(n_1043), .A2(n_811), .A3(n_813), .B(n_834), .Y(n_1046) );
NOR3xp33_ASAP7_75t_L g1047 ( .A(n_1042), .B(n_807), .C(n_769), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_1045), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1046), .Y(n_1049) );
AO22x2_ASAP7_75t_L g1050 ( .A1(n_1047), .A2(n_1042), .B1(n_1041), .B2(n_784), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1049), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1048), .B(n_777), .Y(n_1052) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_1050), .Y(n_1053) );
AND3x1_ASAP7_75t_L g1054 ( .A(n_1051), .B(n_1050), .C(n_828), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_1053), .A2(n_803), .B1(n_806), .B2(n_837), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1052), .Y(n_1056) );
OR2x6_ASAP7_75t_L g1057 ( .A(n_1056), .B(n_822), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_1055), .A2(n_836), .B1(n_946), .B2(n_822), .Y(n_1058) );
NAND3xp33_ASAP7_75t_L g1059 ( .A(n_1054), .B(n_779), .C(n_778), .Y(n_1059) );
AO21x2_ASAP7_75t_L g1060 ( .A1(n_1059), .A2(n_790), .B(n_787), .Y(n_1060) );
OAI21xp5_ASAP7_75t_L g1061 ( .A1(n_1057), .A2(n_832), .B(n_827), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1062 ( .A1(n_1060), .A2(n_1058), .B(n_805), .Y(n_1062) );
OR2x6_ASAP7_75t_L g1063 ( .A(n_1061), .B(n_822), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g1064 ( .A1(n_1063), .A2(n_1062), .B1(n_946), .B2(n_922), .Y(n_1064) );
endmodule