module fake_jpeg_11089_n_649 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_649);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_649;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_61),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_64),
.Y(n_147)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_65),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g173 ( 
.A(n_75),
.Y(n_173)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_82),
.Y(n_193)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_92),
.Y(n_190)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_SL g202 ( 
.A(n_98),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_50),
.B(n_0),
.CON(n_110),
.SN(n_110)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_110),
.B(n_0),
.Y(n_187)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_31),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_116),
.Y(n_137)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_120),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_119),
.Y(n_143)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_42),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_60),
.A2(n_56),
.B1(n_58),
.B2(n_37),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_125),
.A2(n_197),
.B1(n_45),
.B2(n_48),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_128),
.B(n_187),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_32),
.B1(n_23),
.B2(n_34),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_129),
.A2(n_141),
.B1(n_144),
.B2(n_159),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_82),
.A2(n_32),
.B1(n_23),
.B2(n_34),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_66),
.A2(n_32),
.B1(n_34),
.B2(n_52),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_149),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_20),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_162),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_98),
.A2(n_33),
.B1(n_58),
.B2(n_37),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_62),
.B(n_54),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_43),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_91),
.B(n_20),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_85),
.A2(n_37),
.B1(n_58),
.B2(n_42),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_163),
.A2(n_183),
.B1(n_77),
.B2(n_55),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_54),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_175),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_118),
.B(n_44),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_75),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_184),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_110),
.A2(n_56),
.B1(n_58),
.B2(n_37),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_36),
.C(n_21),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_86),
.A2(n_52),
.B1(n_42),
.B2(n_56),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_121),
.B(n_55),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_55),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_188),
.B(n_199),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_113),
.A2(n_52),
.B1(n_42),
.B2(n_59),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_191),
.A2(n_200),
.B1(n_204),
.B2(n_36),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_111),
.A2(n_52),
.B1(n_41),
.B2(n_44),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_55),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_71),
.A2(n_59),
.B1(n_22),
.B2(n_51),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_74),
.A2(n_21),
.B1(n_51),
.B2(n_22),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_205),
.B(n_250),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_122),
.B1(n_120),
.B2(n_103),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_206),
.A2(n_241),
.B1(n_243),
.B2(n_258),
.Y(n_306)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_208),
.Y(n_313)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_210),
.B(n_211),
.Y(n_285)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_202),
.Y(n_212)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_148),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_216),
.B(n_226),
.Y(n_303)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_218),
.Y(n_316)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_129),
.B1(n_191),
.B2(n_144),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_221),
.A2(n_262),
.B1(n_264),
.B2(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_41),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_222),
.B(n_223),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_43),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_143),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_135),
.B(n_49),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_231),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_173),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_239),
.Y(n_307)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_230),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_124),
.B(n_49),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_233),
.A2(n_259),
.B(n_250),
.C(n_267),
.Y(n_311)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_237),
.Y(n_334)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_238),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_173),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_183),
.A2(n_99),
.B1(n_97),
.B2(n_96),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_242),
.Y(n_342)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_157),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_178),
.A2(n_45),
.B1(n_48),
.B2(n_81),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_245),
.A2(n_249),
.B1(n_251),
.B2(n_257),
.Y(n_318)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_246),
.Y(n_293)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_178),
.A2(n_92),
.B1(n_89),
.B2(n_79),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_185),
.A2(n_55),
.B1(n_27),
.B2(n_24),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_252),
.B(n_253),
.Y(n_324)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_254),
.B(n_255),
.Y(n_323)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_256),
.B(n_260),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_185),
.A2(n_27),
.B1(n_24),
.B2(n_18),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_131),
.A2(n_27),
.B1(n_17),
.B2(n_16),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_173),
.A2(n_177),
.B(n_146),
.C(n_204),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_205),
.B(n_227),
.C(n_272),
.Y(n_297)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_266),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_163),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_263),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_179),
.A2(n_27),
.B1(n_17),
.B2(n_14),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_177),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_265),
.B(n_271),
.Y(n_305)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_127),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_267),
.Y(n_329)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_268),
.Y(n_304)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_155),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_177),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_145),
.B(n_0),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_160),
.C(n_147),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_159),
.A2(n_200),
.B1(n_141),
.B2(n_190),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_168),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_274),
.Y(n_335)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_126),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_275),
.Y(n_336)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_189),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_132),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_277),
.A2(n_278),
.B1(n_126),
.B2(n_142),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_164),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_190),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_279),
.Y(n_337)
);

AOI32xp33_ASAP7_75t_L g281 ( 
.A1(n_222),
.A2(n_146),
.A3(n_156),
.B1(n_147),
.B2(n_202),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_281),
.B(n_288),
.C(n_312),
.Y(n_345)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_223),
.B(n_146),
.CI(n_142),
.CON(n_288),
.SN(n_288)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_214),
.B(n_145),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_292),
.B(n_317),
.C(n_321),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_297),
.A2(n_247),
.B1(n_215),
.B2(n_230),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g299 ( 
.A1(n_213),
.A2(n_133),
.B1(n_169),
.B2(n_155),
.Y(n_299)
);

AO21x2_ASAP7_75t_L g355 ( 
.A1(n_299),
.A2(n_311),
.B(n_302),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_214),
.A2(n_153),
.B1(n_133),
.B2(n_201),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_301),
.A2(n_308),
.B1(n_309),
.B2(n_339),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_214),
.A2(n_153),
.B1(n_201),
.B2(n_165),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_231),
.A2(n_150),
.B1(n_132),
.B2(n_165),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_311),
.A2(n_326),
.B1(n_330),
.B2(n_212),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_332),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_160),
.C(n_195),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_211),
.B(n_150),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_340),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_240),
.B(n_138),
.C(n_134),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_208),
.A2(n_171),
.B1(n_138),
.B2(n_134),
.Y(n_326)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_234),
.B(n_171),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_269),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_266),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_248),
.B(n_0),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_250),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_272),
.B(n_1),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_250),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_309),
.B1(n_308),
.B2(n_301),
.Y(n_376)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_SL g396 ( 
.A1(n_345),
.A2(n_366),
.B(n_385),
.Y(n_396)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_346),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_294),
.A2(n_329),
.B1(n_286),
.B2(n_341),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_348),
.A2(n_360),
.B1(n_376),
.B2(n_377),
.Y(n_398)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_220),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_351),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_236),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_286),
.A2(n_243),
.B1(n_244),
.B2(n_242),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_353),
.A2(n_358),
.B1(n_359),
.B2(n_369),
.Y(n_419)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_284),
.Y(n_354)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

OA22x2_ASAP7_75t_L g404 ( 
.A1(n_355),
.A2(n_370),
.B1(n_280),
.B2(n_328),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_307),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_356),
.B(n_361),
.Y(n_401)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_325),
.Y(n_357)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_286),
.A2(n_261),
.B1(n_268),
.B2(n_237),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_306),
.A2(n_238),
.B1(n_255),
.B2(n_256),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_294),
.A2(n_339),
.B1(n_311),
.B2(n_299),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_285),
.B(n_224),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_217),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_364),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_209),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_305),
.A2(n_219),
.B(n_229),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_365),
.A2(n_384),
.B(n_386),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_311),
.A2(n_218),
.B1(n_254),
.B2(n_246),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_311),
.A2(n_299),
.B1(n_292),
.B2(n_297),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_299),
.A2(n_321),
.B1(n_287),
.B2(n_288),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_232),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_392),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_327),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_287),
.A2(n_258),
.B1(n_277),
.B2(n_263),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_303),
.B(n_207),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_379),
.B(n_387),
.Y(n_429)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_279),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_327),
.C(n_314),
.Y(n_397)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_284),
.Y(n_383)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_288),
.A2(n_275),
.B1(n_260),
.B2(n_278),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_313),
.A2(n_235),
.B1(n_3),
.B2(n_4),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_313),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_319),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_282),
.Y(n_388)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_324),
.B(n_1),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_389),
.B(n_333),
.Y(n_437)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g391 ( 
.A(n_283),
.B(n_5),
.C(n_6),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_6),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_6),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_404),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_407),
.C(n_426),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_392),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_8),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_360),
.A2(n_299),
.B1(n_318),
.B2(n_283),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_405),
.B1(n_412),
.B2(n_428),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_348),
.A2(n_335),
.B1(n_336),
.B2(n_314),
.Y(n_405)
);

OAI32xp33_ASAP7_75t_L g406 ( 
.A1(n_371),
.A2(n_351),
.A3(n_350),
.B1(n_347),
.B2(n_369),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_424),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_290),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_355),
.B1(n_367),
.B2(n_370),
.Y(n_412)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_437),
.C(n_393),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_352),
.B(n_290),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_6),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_347),
.B(n_304),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_384),
.A2(n_304),
.B(n_315),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_436),
.B(n_365),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_367),
.B(n_298),
.C(n_338),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_355),
.A2(n_280),
.B1(n_323),
.B2(n_343),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_343),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_345),
.C(n_378),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_382),
.A2(n_323),
.B1(n_293),
.B2(n_282),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_433),
.A2(n_382),
.B1(n_355),
.B2(n_359),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_354),
.B(n_315),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_435),
.B(n_7),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_375),
.A2(n_323),
.B(n_337),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_364),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_446),
.C(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_442),
.A2(n_458),
.B(n_471),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_398),
.A2(n_355),
.B1(n_353),
.B2(n_362),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_461),
.B1(n_423),
.B2(n_427),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_445),
.B(n_468),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_404),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_358),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_396),
.A2(n_346),
.B1(n_344),
.B2(n_349),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_449),
.A2(n_454),
.B1(n_463),
.B2(n_465),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_374),
.C(n_357),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_452),
.C(n_457),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_394),
.A2(n_390),
.B(n_380),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_451),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_298),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_403),
.A2(n_383),
.B1(n_388),
.B2(n_331),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_455),
.Y(n_486)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_411),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_460),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_338),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_403),
.A2(n_373),
.B(n_368),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_459),
.Y(n_503)
);

OA22x2_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_337),
.B1(n_331),
.B2(n_310),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_398),
.A2(n_310),
.B1(n_334),
.B2(n_316),
.Y(n_461)
);

OAI22x1_ASAP7_75t_L g463 ( 
.A1(n_400),
.A2(n_295),
.B1(n_316),
.B2(n_334),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_296),
.C(n_295),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_464),
.B(n_467),
.C(n_466),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_296),
.B1(n_7),
.B2(n_8),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_466),
.B(n_422),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_7),
.C(n_8),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_412),
.A2(n_8),
.B1(n_10),
.B2(n_416),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_469),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_416),
.A2(n_8),
.B1(n_10),
.B2(n_405),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_470),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_425),
.A2(n_394),
.B(n_395),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_473),
.Y(n_493)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_414),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_414),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_475),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_413),
.B(n_10),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_429),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_476),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_413),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_482),
.Y(n_523)
);

XNOR2x2_ASAP7_75t_SL g478 ( 
.A(n_452),
.B(n_424),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_478),
.B(n_415),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_438),
.B(n_397),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_462),
.A2(n_404),
.B1(n_436),
.B2(n_434),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_483),
.B(n_501),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_450),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_492),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_443),
.A2(n_419),
.B1(n_434),
.B2(n_404),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_489),
.A2(n_497),
.B(n_431),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_490),
.A2(n_487),
.B1(n_498),
.B2(n_491),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_421),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_496),
.B(n_505),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_476),
.B(n_401),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_499),
.B(n_500),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_402),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_449),
.A2(n_422),
.B1(n_421),
.B2(n_432),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_502),
.B(n_506),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_439),
.B(n_432),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_451),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_448),
.B(n_427),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_464),
.C(n_467),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_453),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_460),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_442),
.A2(n_471),
.B(n_453),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_510),
.A2(n_453),
.B(n_458),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_512),
.A2(n_520),
.B(n_530),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_513),
.B(n_519),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_484),
.B(n_444),
.C(n_460),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_485),
.C(n_480),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_489),
.A2(n_465),
.B1(n_454),
.B2(n_463),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_515),
.A2(n_525),
.B1(n_529),
.B2(n_536),
.Y(n_546)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_507),
.B(n_475),
.Y(n_517)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_517),
.Y(n_549)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_479),
.Y(n_518)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_518),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_477),
.B(n_461),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_495),
.A2(n_460),
.B(n_474),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_507),
.B(n_440),
.Y(n_521)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_522),
.Y(n_558)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_490),
.A2(n_473),
.B1(n_456),
.B2(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_528),
.A2(n_535),
.B1(n_538),
.B2(n_539),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_495),
.A2(n_441),
.B1(n_459),
.B2(n_410),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_494),
.B(n_402),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_531),
.B(n_534),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_431),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_415),
.Y(n_535)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_504),
.Y(n_539)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_504),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_541),
.A2(n_483),
.B1(n_497),
.B2(n_511),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_542),
.B(n_496),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_544),
.B(n_561),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_482),
.C(n_480),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_545),
.B(n_547),
.C(n_553),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_485),
.C(n_505),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_508),
.C(n_509),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_510),
.C(n_488),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_559),
.C(n_540),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_516),
.A2(n_497),
.B(n_491),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_557),
.B(n_567),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_519),
.C(n_513),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_478),
.Y(n_561)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_562),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_542),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_512),
.A2(n_488),
.B(n_493),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_565),
.A2(n_556),
.B(n_552),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_536),
.A2(n_493),
.B1(n_502),
.B2(n_503),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_566),
.A2(n_524),
.B1(n_528),
.B2(n_518),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_514),
.A2(n_521),
.B(n_537),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_537),
.A2(n_10),
.B1(n_417),
.B2(n_534),
.Y(n_568)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_568),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_550),
.A2(n_520),
.B(n_530),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_569),
.A2(n_579),
.B(n_550),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_533),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_572),
.B(n_582),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_547),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_578),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_549),
.B(n_517),
.Y(n_576)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_576),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_543),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_577),
.B(n_589),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_553),
.B(n_541),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_556),
.A2(n_539),
.B1(n_533),
.B2(n_515),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_580),
.A2(n_583),
.B1(n_568),
.B2(n_557),
.Y(n_599)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_581),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_565),
.B(n_538),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_529),
.C(n_525),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_584),
.B(n_588),
.C(n_544),
.Y(n_591)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_558),
.Y(n_585)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_585),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_560),
.B(n_559),
.C(n_545),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_563),
.Y(n_589)
);

CKINVDCx14_ASAP7_75t_R g590 ( 
.A(n_551),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_590),
.B(n_558),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_591),
.B(n_607),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_576),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_592),
.B(n_595),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_587),
.A2(n_562),
.B(n_555),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_596),
.A2(n_597),
.B(n_605),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_604),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_582),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_600),
.A2(n_603),
.B1(n_571),
.B2(n_583),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_580),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_569),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_589),
.A2(n_546),
.B1(n_566),
.B2(n_567),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_587),
.A2(n_546),
.B(n_522),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_561),
.C(n_564),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_570),
.C(n_584),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_609),
.B(n_610),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_578),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_612),
.B(n_614),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_573),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_599),
.A2(n_571),
.B1(n_587),
.B2(n_574),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_615),
.A2(n_602),
.B1(n_600),
.B2(n_598),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_608),
.B(n_570),
.C(n_575),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_622),
.Y(n_631)
);

BUFx24_ASAP7_75t_SL g617 ( 
.A(n_608),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_617),
.B(n_586),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_620),
.B(n_621),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_597),
.A2(n_577),
.B(n_581),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_586),
.C(n_574),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_618),
.B(n_598),
.Y(n_624)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_624),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_626),
.A2(n_622),
.B(n_607),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_616),
.B(n_596),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_627),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_619),
.A2(n_602),
.B(n_601),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_628),
.A2(n_593),
.B(n_606),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_629),
.B(n_620),
.C(n_605),
.Y(n_637)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_612),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_630),
.A2(n_593),
.B(n_614),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_631),
.A2(n_613),
.B(n_609),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_633),
.B(n_637),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_636),
.B(n_623),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_638),
.A2(n_639),
.B(n_632),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_640),
.B(n_641),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_634),
.B(n_625),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_643),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_644),
.A2(n_642),
.B(n_632),
.Y(n_646)
);

OAI321xp33_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_645),
.A3(n_625),
.B1(n_635),
.B2(n_606),
.C(n_585),
.Y(n_647)
);

OAI32xp33_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_526),
.A3(n_417),
.B1(n_611),
.B2(n_10),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_611),
.Y(n_649)
);


endmodule