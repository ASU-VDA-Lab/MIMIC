module fake_jpeg_18993_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_38),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_69),
.C(n_74),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_67),
.B1(n_78),
.B2(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_79),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_19),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_70),
.B1(n_83),
.B2(n_35),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_37),
.B1(n_19),
.B2(n_32),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_36),
.B1(n_39),
.B2(n_32),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_32),
.B1(n_15),
.B2(n_23),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_37),
.B1(n_22),
.B2(n_26),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_81),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_37),
.B1(n_23),
.B2(n_28),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_35),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_100),
.B1(n_107),
.B2(n_34),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_99),
.B1(n_109),
.B2(n_34),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_22),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_28),
.B1(n_27),
.B2(n_15),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_27),
.B1(n_25),
.B2(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_112),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_67),
.B1(n_78),
.B2(n_58),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_35),
.B1(n_34),
.B2(n_18),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_13),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_57),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_126),
.C(n_87),
.Y(n_171)
);

OAI22x1_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_74),
.B1(n_70),
.B2(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_133),
.B1(n_138),
.B2(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_65),
.B1(n_64),
.B2(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_125),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_66),
.B1(n_64),
.B2(n_76),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_81),
.B1(n_56),
.B2(n_75),
.Y(n_123)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_74),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_130),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_72),
.B1(n_68),
.B2(n_80),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_131),
.B1(n_102),
.B2(n_94),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_31),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_17),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_17),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_109),
.B1(n_112),
.B2(n_90),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_86),
.B(n_111),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_34),
.B1(n_12),
.B2(n_2),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_142),
.A2(n_5),
.B(n_6),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_86),
.B(n_93),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_151),
.B(n_152),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_144),
.B(n_158),
.Y(n_201)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_103),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_96),
.B(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_96),
.B(n_98),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_24),
.B(n_4),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_103),
.B(n_87),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_98),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_133),
.B1(n_141),
.B2(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_126),
.C(n_143),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_16),
.C(n_17),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_20),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_114),
.A2(n_102),
.B1(n_94),
.B2(n_12),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_117),
.B1(n_123),
.B2(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_168),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_178),
.B1(n_144),
.B2(n_149),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_117),
.B(n_130),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_198),
.B(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_204),
.C(n_152),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_179),
.A2(n_193),
.B1(n_194),
.B2(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_30),
.B1(n_18),
.B2(n_16),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_190),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_16),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_191),
.Y(n_206)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_30),
.B1(n_71),
.B2(n_20),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_20),
.B1(n_24),
.B2(n_3),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_202),
.B1(n_203),
.B2(n_163),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_5),
.C(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_227),
.B1(n_193),
.B2(n_190),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_223),
.Y(n_233)
);

OA21x2_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_172),
.B(n_156),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_156),
.C(n_164),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_183),
.C(n_153),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_224),
.B1(n_226),
.B2(n_203),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_166),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_195),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_165),
.B1(n_148),
.B2(n_150),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_178),
.B1(n_200),
.B2(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_155),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_182),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_154),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_160),
.C(n_157),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_198),
.C(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_210),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_181),
.B1(n_186),
.B2(n_196),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_183),
.B1(n_188),
.B2(n_185),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_247),
.C(n_211),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_218),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_199),
.C(n_188),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.C(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_199),
.C(n_185),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_206),
.B(n_179),
.CI(n_194),
.CON(n_244),
.SN(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_213),
.B1(n_207),
.B2(n_208),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_244),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_255),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_206),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_235),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_223),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_145),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_214),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_219),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_221),
.C(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_238),
.C(n_242),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_234),
.C(n_244),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_190),
.B1(n_8),
.B2(n_9),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_207),
.B1(n_230),
.B2(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_232),
.B(n_208),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_8),
.B(n_10),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_237),
.C(n_226),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_259),
.C(n_260),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_231),
.B(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_8),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.C(n_268),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_257),
.B(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_250),
.C(n_254),
.Y(n_281)
);

NAND2x1_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_7),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_7),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_274),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_265),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_286),
.A2(n_278),
.B(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_296),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_268),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_266),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_279),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_277),
.C(n_290),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_283),
.B1(n_285),
.B2(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_292),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_306),
.B(n_307),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_299),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_309),
.A2(n_302),
.B(n_300),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_303),
.B(n_277),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_10),
.C(n_11),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_10),
.Y(n_313)
);


endmodule