module real_jpeg_12413_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_213;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_57),
.B(n_63),
.C(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_3),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_3),
.B(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_58),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_SL g202 ( 
.A1(n_3),
.A2(n_58),
.B(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_25),
.C(n_40),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_103),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_3),
.A2(n_24),
.B1(n_28),
.B2(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_3),
.B(n_81),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_5),
.A2(n_25),
.B1(n_33),
.B2(n_68),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_6),
.A2(n_25),
.B1(n_33),
.B2(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_6),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_25),
.B1(n_33),
.B2(n_73),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_73),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_25),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_11),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_110),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_110),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_13),
.A2(n_25),
.B1(n_33),
.B2(n_110),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_14),
.A2(n_25),
.B1(n_33),
.B2(n_70),
.Y(n_219)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_138),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_20),
.B(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_95),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_21),
.B(n_83),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_52),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_22),
.B(n_53),
.C(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_23),
.B(n_38),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_24),
.A2(n_28),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_24),
.A2(n_28),
.B1(n_217),
.B2(n_225),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_24),
.A2(n_87),
.B(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_28),
.B(n_103),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_29),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_29),
.A2(n_31),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_29),
.A2(n_89),
.B(n_99),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_29),
.A2(n_98),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_33),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_35),
.A2(n_88),
.B(n_98),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_48),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_39),
.B(n_103),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_43),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_45),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_SL g189 ( 
.A(n_44),
.B(n_59),
.C(n_76),
.Y(n_189)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_45),
.A2(n_77),
.B(n_187),
.C(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_45),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_49),
.B(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_93),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_50),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_50),
.A2(n_92),
.B1(n_182),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_50),
.A2(n_92),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_50),
.A2(n_92),
.B1(n_204),
.B2(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_71),
.B2(n_82),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_67),
.B2(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_56),
.B1(n_67),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_69),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_59),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_61),
.B(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_74),
.A2(n_75),
.B1(n_105),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_74),
.A2(n_75),
.B1(n_148),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_74),
.A2(n_75),
.B1(n_164),
.B2(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_92),
.B(n_153),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_95),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.C(n_108),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_96),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_108),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_136),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_121),
.B1(n_134),
.B2(n_135),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_171),
.B(n_250),
.C(n_254),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_140),
.B(n_165),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_155),
.C(n_158),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_149),
.C(n_154),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_154),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_248),
.B(n_249),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_192),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_177),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_184),
.B1(n_185),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_205),
.B(n_247),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_197),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.C(n_203),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_241),
.B(n_246),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_231),
.B(n_240),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_220),
.B(n_230),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_215),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_226),
.B(n_229),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_233),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_236),
.C(n_239),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_245),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_253),
.Y(n_254)
);


endmodule