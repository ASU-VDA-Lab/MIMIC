module fake_jpeg_2088_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_0),
.B(n_1),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_21),
.B(n_36),
.C(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_33),
.B1(n_22),
.B2(n_30),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_77),
.B1(n_96),
.B2(n_99),
.Y(n_116)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_60),
.A2(n_63),
.B(n_98),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_28),
.B1(n_25),
.B2(n_32),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_65),
.A2(n_92),
.B1(n_95),
.B2(n_32),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_20),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_87),
.Y(n_121)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_30),
.B1(n_17),
.B2(n_20),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_56),
.B1(n_46),
.B2(n_21),
.Y(n_106)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_24),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_28),
.B1(n_25),
.B2(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_32),
.B1(n_17),
.B2(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_39),
.A2(n_17),
.B1(n_42),
.B2(n_56),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_12),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_10),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_37),
.B(n_36),
.C(n_34),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_39),
.A2(n_37),
.B1(n_15),
.B2(n_24),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_128),
.B1(n_135),
.B2(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_46),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_31),
.B(n_26),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_78),
.B(n_86),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_82),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_122),
.B(n_125),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_26),
.B1(n_31),
.B2(n_10),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_67),
.B(n_84),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_0),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_0),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_95),
.B1(n_92),
.B2(n_91),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_4),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_61),
.B(n_31),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_64),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_138),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_67),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_64),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_147),
.B1(n_137),
.B2(n_112),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_62),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_143),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_79),
.B1(n_74),
.B2(n_70),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_150),
.B1(n_133),
.B2(n_123),
.Y(n_185)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_74),
.B1(n_70),
.B2(n_62),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_149),
.B(n_108),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_79),
.B(n_81),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_81),
.B1(n_76),
.B2(n_75),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_75),
.B(n_2),
.C(n_3),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_129),
.B(n_9),
.C(n_8),
.D(n_105),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_120),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_121),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_157),
.C(n_160),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_1),
.C(n_2),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_3),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_131),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_4),
.C(n_5),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_106),
.A2(n_122),
.B1(n_113),
.B2(n_128),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_133),
.B1(n_138),
.B2(n_136),
.Y(n_181)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_5),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_6),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_8),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_8),
.C(n_9),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_167),
.C(n_160),
.Y(n_213)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_177),
.Y(n_195)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_179),
.B(n_180),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_119),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_181),
.A2(n_182),
.B1(n_187),
.B2(n_211),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_105),
.B1(n_126),
.B2(n_127),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_201),
.B1(n_155),
.B2(n_174),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_133),
.B(n_112),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_173),
.B(n_151),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_190),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_145),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_119),
.B(n_132),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_203),
.B(n_211),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_132),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_196),
.Y(n_224)
);

AO21x2_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_144),
.B(n_172),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_127),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_205),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_146),
.A2(n_108),
.B1(n_105),
.B2(n_129),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_141),
.A2(n_129),
.B(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_153),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_208),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_169),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_162),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_216),
.B(n_184),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_221),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_153),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_158),
.B(n_152),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_226),
.B(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_187),
.B1(n_191),
.B2(n_193),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_184),
.B(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_235),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_171),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_177),
.B1(n_165),
.B2(n_168),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_233),
.A2(n_236),
.B1(n_207),
.B2(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_176),
.B1(n_182),
.B2(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_240),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_194),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_207),
.B1(n_200),
.B2(n_188),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_217),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_250),
.B1(n_259),
.B2(n_260),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_249),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_205),
.B1(n_202),
.B2(n_211),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_262),
.B1(n_263),
.B2(n_229),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_255),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_223),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_228),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

INVx3_ASAP7_75t_SL g258 ( 
.A(n_216),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_236),
.B1(n_240),
.B2(n_226),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_183),
.B1(n_213),
.B2(n_206),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_214),
.A2(n_183),
.B1(n_196),
.B2(n_210),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_239),
.B1(n_225),
.B2(n_222),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_277),
.B1(n_250),
.B2(n_257),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_221),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_274),
.C(n_275),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_264),
.B(n_261),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_280),
.B1(n_267),
.B2(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_232),
.C(n_220),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_219),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_218),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_279),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_238),
.B1(n_233),
.B2(n_224),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_217),
.C(n_224),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_238),
.B1(n_235),
.B2(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_255),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_296),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_278),
.B1(n_269),
.B2(n_251),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_264),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_276),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_269),
.B(n_251),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_249),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_265),
.B1(n_278),
.B2(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_263),
.CI(n_243),
.CON(n_295),
.SN(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_297),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_247),
.C(n_256),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_297),
.B1(n_284),
.B2(n_295),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_266),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_306),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_295),
.B(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_283),
.B1(n_292),
.B2(n_286),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_242),
.B(n_245),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_262),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_284),
.C(n_289),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_317),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_300),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_178),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_178),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_320),
.Y(n_325)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_328),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_299),
.B(n_309),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_304),
.B(n_306),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_299),
.B(n_304),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_330),
.B(n_331),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_319),
.C(n_302),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_313),
.B(n_245),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_322),
.Y(n_335)
);

AO221x1_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_328),
.B1(n_321),
.B2(n_326),
.C(n_307),
.Y(n_337)
);

AOI31xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_334),
.A3(n_336),
.B(n_210),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_199),
.B(n_178),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_199),
.Y(n_342)
);


endmodule