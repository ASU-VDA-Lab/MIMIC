module real_jpeg_12345_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_289, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_289;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_211;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_0),
.A2(n_38),
.B1(n_68),
.B2(n_69),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_0),
.A2(n_38),
.B1(n_57),
.B2(n_58),
.Y(n_226)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_285),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_4),
.B(n_286),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_47),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_47),
.B1(n_68),
.B2(n_69),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_10),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_24),
.B1(n_57),
.B2(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_24),
.B1(n_68),
.B2(n_69),
.Y(n_206)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_11),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_12),
.A2(n_20),
.B1(n_21),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_28),
.B(n_54),
.C(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_49),
.B1(n_68),
.B2(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_12),
.B(n_26),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_12),
.B(n_66),
.C(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_12),
.B(n_59),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_29),
.C(n_31),
.Y(n_170)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_40),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_39),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_35),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_19),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_34)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_21),
.B(n_170),
.Y(n_169)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_25),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_33),
.B1(n_45),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_27),
.A2(n_37),
.B(n_78),
.Y(n_77)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_27),
.A2(n_46),
.B(n_78),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_28),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_35),
.B(n_42),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_79),
.B(n_284),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_74),
.C(n_77),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_43),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.C(n_61),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_44),
.A2(n_120),
.B1(n_122),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_44),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_44),
.B(n_120),
.C(n_183),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_44),
.A2(n_88),
.B1(n_89),
.B2(n_185),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_44),
.A2(n_185),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_48),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_55),
.B(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_49),
.B(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_49),
.B(n_72),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_50),
.A2(n_61),
.B1(n_259),
.B2(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_50),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_52),
.A2(n_59),
.B1(n_92),
.B2(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_56),
.A2(n_76),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_56),
.A2(n_91),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_58),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_61),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_61),
.B(n_173),
.C(n_260),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_72),
.B(n_73),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_62),
.A2(n_72),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_97),
.Y(n_96)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_67),
.B1(n_95),
.B2(n_97),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_63),
.A2(n_67),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_68),
.B(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_94),
.B(n_96),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_72),
.A2(n_96),
.B(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_73),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_74),
.B(n_77),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_279),
.B(n_283),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_251),
.B(n_276),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_230),
.B(n_250),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_213),
.B(n_229),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_180),
.A3(n_208),
.B1(n_211),
.B2(n_212),
.C(n_289),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_162),
.B(n_179),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_128),
.B(n_161),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_109),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_87),
.B(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_98),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_88),
.A2(n_89),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_89),
.B(n_172),
.C(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_89),
.B(n_185),
.C(n_218),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_93),
.A2(n_132),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_93),
.A2(n_145),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_98),
.A2(n_99),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_104),
.B(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_107),
.A2(n_108),
.B1(n_188),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_108),
.A2(n_118),
.B(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_123),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_125),
.C(n_126),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_120),
.B2(n_122),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_116),
.C(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_120),
.A2(n_245),
.B(n_248),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_120),
.B(n_245),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_127),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_137),
.C(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_125),
.A2(n_127),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_125),
.B(n_205),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_155),
.B(n_160),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_141),
.B(n_154),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_139),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_168),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_146),
.B(n_153),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_187),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B(n_152),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_167),
.C(n_171),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_173),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_195),
.C(n_200),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_172),
.A2(n_173),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_172),
.A2(n_173),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_173),
.B(n_270),
.C(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_190),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_182),
.B(n_186),
.CI(n_190),
.CON(n_210),
.SN(n_210)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_207),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_202),
.B2(n_203),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_203),
.C(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_210),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_228),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_228),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_217),
.C(n_222),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_227),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_236),
.B(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_249),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_243),
.B2(n_244),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_243),
.C(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_255),
.B1(n_256),
.B2(n_263),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_266),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_265),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_265),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_264),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_263),
.C(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_260),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_275),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_275),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_282),
.Y(n_283)
);


endmodule