module fake_netlist_1_10351_n_255 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_255);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_255;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_214;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_88;
wire n_244;
wire n_102;
wire n_141;
wire n_119;
wire n_115;
wire n_97;
wire n_167;
wire n_107;
wire n_158;
wire n_114;
wire n_121;
wire n_171;
wire n_94;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_137;
wire n_87;
wire n_180;
wire n_104;
wire n_160;
wire n_98;
wire n_206;
wire n_154;
wire n_195;
wire n_165;
wire n_146;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_215;
wire n_91;
wire n_155;
wire n_108;
wire n_116;
wire n_209;
wire n_217;
wire n_139;
wire n_229;
wire n_230;
wire n_198;
wire n_169;
wire n_193;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_156;
wire n_124;
wire n_95;
wire n_238;
wire n_128;
wire n_120;
wire n_129;
wire n_90;
wire n_135;
wire n_188;
wire n_247;
wire n_197;
wire n_201;
wire n_242;
wire n_127;
wire n_170;
wire n_157;
wire n_111;
wire n_202;
wire n_210;
wire n_142;
wire n_184;
wire n_245;
wire n_191;
wire n_232;
wire n_200;
wire n_208;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_178;
wire n_118;
wire n_253;
wire n_179;
wire n_131;
wire n_112;
wire n_205;
wire n_86;
wire n_143;
wire n_213;
wire n_235;
wire n_243;
wire n_182;
wire n_166;
wire n_162;
wire n_186;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_248;
wire n_231;
wire n_136;
wire n_176;
wire n_89;
wire n_144;
wire n_183;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_251;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_246;
wire n_153;
wire n_99;
wire n_132;
wire n_109;
wire n_93;
wire n_151;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_225;
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_79), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_20), .Y(n_87) );
INVx3_ASAP7_75t_L g88 ( .A(n_33), .Y(n_88) );
NOR2xp33_ASAP7_75t_L g89 ( .A(n_57), .B(n_71), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_9), .Y(n_90) );
NOR2xp67_ASAP7_75t_L g91 ( .A(n_45), .B(n_69), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_84), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_65), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_49), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_85), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_77), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_61), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_73), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_24), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_76), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_56), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_64), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_80), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_55), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_46), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_38), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_51), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_43), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_52), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_11), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_36), .B(n_28), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_30), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_32), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_72), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_26), .Y(n_121) );
INVx2_ASAP7_75t_SL g122 ( .A(n_44), .Y(n_122) );
BUFx5_ASAP7_75t_L g123 ( .A(n_75), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_13), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_68), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_74), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_70), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_22), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_54), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_8), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_53), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_31), .Y(n_132) );
BUFx10_ASAP7_75t_L g133 ( .A(n_37), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_15), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_63), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_124), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_88), .B(n_0), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_88), .B(n_0), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_104), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_134), .B(n_4), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_90), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_106), .B(n_5), .Y(n_143) );
INVxp67_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_122), .B(n_7), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_137), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_138), .B(n_148), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
NAND2xp33_ASAP7_75t_L g155 ( .A(n_143), .B(n_123), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_159), .B(n_136), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_149), .B(n_133), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_153), .B(n_86), .Y(n_164) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_152), .B(n_141), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_150), .B(n_157), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_155), .B(n_139), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_158), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_156), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_166), .A2(n_96), .B(n_95), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_165), .A2(n_127), .B1(n_131), .B2(n_125), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_167), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_161), .A2(n_130), .B(n_121), .C(n_98), .Y(n_175) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_160), .A2(n_102), .B(n_92), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_163), .A2(n_97), .B(n_103), .C(n_100), .Y(n_177) );
CKINVDCx10_ASAP7_75t_R g178 ( .A(n_168), .Y(n_178) );
OAI21xp33_ASAP7_75t_L g179 ( .A1(n_164), .A2(n_101), .B(n_99), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_173), .B(n_91), .Y(n_180) );
OAI21x1_ASAP7_75t_L g181 ( .A1(n_176), .A2(n_170), .B(n_108), .Y(n_181) );
AO31x2_ASAP7_75t_L g182 ( .A1(n_177), .A2(n_109), .A3(n_110), .B(n_107), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_172), .B(n_105), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_174), .A2(n_169), .B(n_167), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_175), .A2(n_119), .B(n_120), .C(n_118), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_171), .A2(n_114), .B(n_89), .Y(n_186) );
INVx5_ASAP7_75t_L g187 ( .A(n_174), .Y(n_187) );
OAI21xp5_ASAP7_75t_SL g188 ( .A1(n_178), .A2(n_115), .B(n_94), .Y(n_188) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_112), .B(n_111), .Y(n_189) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_181), .A2(n_117), .B(n_116), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_185), .B(n_10), .Y(n_191) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_184), .A2(n_129), .B(n_117), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_187), .Y(n_193) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_186), .A2(n_128), .B(n_126), .Y(n_194) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_180), .A2(n_135), .B(n_132), .Y(n_195) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_180), .A2(n_25), .B(n_23), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_187), .B(n_12), .Y(n_197) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_182), .A2(n_47), .A3(n_83), .B(n_82), .Y(n_198) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_189), .A2(n_29), .B(n_27), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_183), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_200) );
AO22x1_ASAP7_75t_L g201 ( .A1(n_188), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_193), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_197), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_197), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_190), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_192), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_191), .A2(n_19), .B(n_20), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_196), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_198), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_201), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_194), .B(n_21), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_200), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_195), .Y(n_213) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_199), .A2(n_34), .B(n_35), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_193), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_212), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_215), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_202), .B(n_42), .Y(n_218) );
INVxp67_ASAP7_75t_SL g219 ( .A(n_210), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_211), .Y(n_220) );
OR2x2_ASAP7_75t_L g221 ( .A(n_203), .B(n_81), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_204), .B(n_48), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_207), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_208), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_207), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_209), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_219), .B(n_206), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_220), .B(n_205), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_224), .B(n_214), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_217), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_226), .B(n_214), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_223), .B(n_59), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_225), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_235), .Y(n_236) );
AND2x4_ASAP7_75t_SL g237 ( .A(n_231), .B(n_218), .Y(n_237) );
INVx1_ASAP7_75t_SL g238 ( .A(n_237), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_236), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_238), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_239), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_240), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_242), .B(n_241), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_243), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_244), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_245), .B(n_228), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_246), .B(n_233), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_247), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_248), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_249), .A2(n_216), .B1(n_221), .B2(n_222), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_250), .B(n_229), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_251), .Y(n_252) );
NOR2xp33_ASAP7_75t_R g253 ( .A(n_252), .B(n_66), .Y(n_253) );
NOR2x1_ASAP7_75t_L g254 ( .A(n_253), .B(n_232), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_254), .A2(n_229), .B1(n_230), .B2(n_234), .Y(n_255) );
endmodule