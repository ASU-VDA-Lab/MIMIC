module fake_jpeg_4385_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_0),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_2),
.C(n_3),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_8),
.B(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_10),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_11),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_12),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_34),
.B(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

OAI22x1_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_35),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_14),
.B(n_7),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_28),
.C(n_32),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_7),
.B1(n_13),
.B2(n_26),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_25),
.C(n_29),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_38),
.Y(n_48)
);

AOI221xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_37),
.B1(n_41),
.B2(n_39),
.C(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_48),
.C(n_45),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_42),
.Y(n_51)
);


endmodule