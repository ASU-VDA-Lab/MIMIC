module fake_jpeg_9475_n_144 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_19),
.B(n_26),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_29),
.C(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_27),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_35),
.B1(n_37),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_58),
.B1(n_66),
.B2(n_70),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_37),
.B1(n_31),
.B2(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_31),
.B1(n_18),
.B2(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_29),
.B1(n_16),
.B2(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_20),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_46),
.B(n_42),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_82),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_45),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_46),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_42),
.B(n_50),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_63),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_96),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_73),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_55),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_101),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_100),
.B(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_110),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_86),
.A3(n_84),
.B1(n_87),
.B2(n_76),
.C1(n_79),
.C2(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_86),
.C(n_13),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_95),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_101),
.B1(n_94),
.B2(n_100),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_112),
.B1(n_114),
.B2(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_56),
.C(n_15),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_64),
.B1(n_15),
.B2(n_1),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_109),
.B(n_42),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_128),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_109),
.C(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_115),
.B(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_135),
.B(n_137),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_3),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_129),
.B1(n_116),
.B2(n_130),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_125),
.A3(n_120),
.B1(n_121),
.B2(n_11),
.C1(n_3),
.C2(n_8),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_7),
.B1(n_12),
.B2(n_139),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_7),
.B(n_12),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);


endmodule