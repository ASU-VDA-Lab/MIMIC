module fake_jpeg_30351_n_504 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_504);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_504;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_60),
.Y(n_105)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_54),
.B(n_57),
.Y(n_156)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_63),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx6f_ASAP7_75t_SL g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_72),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_86),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_1),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_91),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_34),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx16f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_97),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_27),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_49),
.Y(n_138)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_29),
.B1(n_33),
.B2(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_104),
.A2(n_126),
.B1(n_131),
.B2(n_149),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g195 ( 
.A(n_113),
.Y(n_195)
);

NAND2xp67_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_38),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_26),
.C(n_37),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_51),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_18),
.B1(n_28),
.B2(n_41),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_67),
.B(n_49),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_88),
.B(n_47),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_58),
.A2(n_33),
.B1(n_41),
.B2(n_28),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_47),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_36),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_101),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_69),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_96),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_89),
.Y(n_181)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_163),
.Y(n_255)
);

CKINVDCx9p33_ASAP7_75t_R g164 ( 
.A(n_107),
.Y(n_164)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_39),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_165),
.B(n_169),
.Y(n_241)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_80),
.C(n_53),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_167),
.B(n_177),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_36),
.B1(n_37),
.B2(n_30),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_185),
.B(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_121),
.A2(n_76),
.B1(n_66),
.B2(n_94),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_174),
.A2(n_194),
.B1(n_103),
.B2(n_135),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_70),
.B1(n_77),
.B2(n_61),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_175),
.A2(n_191),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_87),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_184),
.Y(n_221)
);

INVxp67_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_187),
.B(n_143),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_105),
.B(n_85),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_132),
.A2(n_82),
.B1(n_73),
.B2(n_26),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_136),
.B1(n_115),
.B2(n_148),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_30),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_105),
.A2(n_98),
.B1(n_102),
.B2(n_63),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_67),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_41),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_196),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_131),
.A2(n_89),
.B1(n_41),
.B2(n_33),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_33),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_104),
.A2(n_33),
.B(n_28),
.C(n_18),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_115),
.B(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_199),
.B(n_200),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_110),
.B(n_28),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_123),
.B(n_28),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_204),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_18),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_124),
.B(n_18),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_207),
.Y(n_238)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_208),
.Y(n_258)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_113),
.B(n_1),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_217),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_146),
.B(n_3),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_218),
.Y(n_232)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_149),
.B(n_3),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_114),
.B(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_143),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_250),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_153),
.B(n_119),
.C(n_127),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_225),
.B(n_218),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_226),
.B(n_246),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_230),
.B1(n_243),
.B2(n_252),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_229),
.A2(n_212),
.B(n_183),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_177),
.A2(n_136),
.B1(n_155),
.B2(n_134),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_245),
.B1(n_248),
.B2(n_262),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_185),
.A2(n_155),
.B1(n_134),
.B2(n_129),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_129),
.B1(n_125),
.B2(n_118),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_185),
.A2(n_109),
.B1(n_147),
.B2(n_125),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_174),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_179),
.B(n_7),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_167),
.B(n_15),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_15),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_15),
.B1(n_10),
.B2(n_11),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_184),
.B(n_178),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_168),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_191),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_266),
.B(n_294),
.Y(n_330)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_193),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_277),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_194),
.C(n_203),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_274),
.C(n_278),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_272),
.A2(n_276),
.B(n_290),
.Y(n_329)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_203),
.C(n_175),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_164),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_214),
.C(n_212),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_163),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_286),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_239),
.B(n_162),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_281),
.B(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_235),
.B(n_197),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_284),
.B(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_221),
.B(n_163),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_289),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_254),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_240),
.A2(n_216),
.B1(n_215),
.B2(n_173),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_235),
.B(n_210),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_296),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_232),
.B(n_259),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_171),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_232),
.B(n_209),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_298),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_240),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_302),
.Y(n_320)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_236),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_237),
.B1(n_231),
.B2(n_249),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_250),
.B(n_195),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_SL g303 ( 
.A(n_232),
.B(n_220),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_223),
.C(n_232),
.Y(n_305)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_264),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_278),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_245),
.B1(n_233),
.B2(n_229),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_317),
.B1(n_323),
.B2(n_326),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_310),
.B(n_289),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_220),
.B(n_251),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_314),
.A2(n_324),
.B(n_298),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_248),
.B1(n_252),
.B2(n_246),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_318),
.A2(n_340),
.B(n_207),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_295),
.A2(n_262),
.B1(n_232),
.B2(n_260),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_256),
.B(n_241),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_228),
.B1(n_254),
.B2(n_231),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_325),
.A2(n_331),
.B1(n_338),
.B2(n_310),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_274),
.A2(n_270),
.B1(n_265),
.B2(n_282),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_327),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_265),
.A2(n_264),
.B1(n_166),
.B2(n_249),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_257),
.C(n_258),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_180),
.C(n_195),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_276),
.A2(n_261),
.B1(n_205),
.B2(n_201),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_334),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_271),
.A2(n_237),
.B1(n_257),
.B2(n_244),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_271),
.B(n_258),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_283),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_266),
.A2(n_238),
.B1(n_242),
.B2(n_244),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_292),
.A2(n_238),
.B(n_208),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_342),
.B(n_363),
.Y(n_391)
);

INVx13_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

BUFx24_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_353),
.Y(n_375)
);

INVx13_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

AOI322xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_279),
.A3(n_301),
.B1(n_288),
.B2(n_297),
.C1(n_267),
.C2(n_299),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_346),
.B(n_347),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_319),
.B(n_279),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_275),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_330),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_360),
.Y(n_393)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_325),
.A2(n_285),
.B1(n_286),
.B2(n_289),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_356),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_355),
.A2(n_322),
.B1(n_316),
.B2(n_339),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_277),
.B1(n_300),
.B2(n_302),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_357),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_291),
.Y(n_358)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_322),
.Y(n_360)
);

A2O1A1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_298),
.B(n_273),
.C(n_304),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_361),
.A2(n_309),
.B(n_319),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_298),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_364),
.Y(n_384)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_329),
.B(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_335),
.B(n_206),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_368),
.Y(n_400)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_371),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_307),
.A2(n_180),
.B1(n_10),
.B2(n_11),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_333),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_336),
.B(n_321),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_372),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_373),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_363),
.A2(n_318),
.B(n_332),
.Y(n_374)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_379),
.B(n_382),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_359),
.A2(n_308),
.B1(n_329),
.B2(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_392),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_377),
.A2(n_397),
.B1(n_356),
.B2(n_354),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_350),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_315),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_366),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_359),
.A2(n_308),
.B1(n_338),
.B2(n_324),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_336),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_398),
.C(n_305),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_321),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_305),
.C(n_323),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_398),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_409),
.Y(n_434)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_362),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_411),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_370),
.B1(n_347),
.B2(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_406),
.B(n_413),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_393),
.A2(n_349),
.B1(n_353),
.B2(n_341),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_408),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_341),
.B1(n_364),
.B2(n_352),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_365),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_412),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_384),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_375),
.A2(n_358),
.B1(n_344),
.B2(n_361),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_415),
.A2(n_418),
.B1(n_422),
.B2(n_381),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_424),
.B1(n_380),
.B2(n_373),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_375),
.A2(n_368),
.B1(n_309),
.B2(n_316),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_334),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_420),
.C(n_421),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_320),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_320),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_380),
.A2(n_339),
.B1(n_311),
.B2(n_372),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_312),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_423),
.B(n_425),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_377),
.A2(n_357),
.B1(n_312),
.B2(n_367),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_8),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_418),
.Y(n_427)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_430),
.Y(n_449)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_419),
.A2(n_392),
.B1(n_376),
.B2(n_377),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_443),
.B1(n_386),
.B2(n_378),
.Y(n_458)
);

XOR2x1_ASAP7_75t_SL g433 ( 
.A(n_410),
.B(n_382),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_433),
.A2(n_411),
.B(n_401),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_395),
.C(n_391),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_441),
.C(n_409),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_438),
.A2(n_414),
.B1(n_394),
.B2(n_396),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_384),
.C(n_381),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_422),
.A2(n_383),
.B1(n_394),
.B2(n_396),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_378),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_416),
.A2(n_414),
.B(n_383),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_445),
.B(n_416),
.Y(n_453)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_436),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_447),
.B(n_442),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_417),
.Y(n_448)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_448),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_421),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_450),
.B(n_451),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_441),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_454),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_453),
.A2(n_456),
.B1(n_460),
.B2(n_429),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_430),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_440),
.B(n_420),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_459),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_457),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_458),
.A2(n_427),
.B1(n_428),
.B2(n_426),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_432),
.B(n_386),
.Y(n_459)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_463),
.B(n_387),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_434),
.C(n_432),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_470),
.C(n_387),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_446),
.B(n_426),
.Y(n_468)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_468),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_472),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_434),
.C(n_435),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_449),
.A2(n_442),
.B1(n_431),
.B2(n_443),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_473),
.B1(n_463),
.B2(n_462),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_457),
.A2(n_445),
.B1(n_437),
.B2(n_387),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_474),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_476),
.A2(n_481),
.B(n_480),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_484),
.C(n_468),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_482),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_462),
.A2(n_345),
.B(n_343),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_367),
.C(n_345),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_483),
.B(n_470),
.C(n_473),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_471),
.A2(n_343),
.B1(n_12),
.B2(n_13),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_487),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_486),
.A2(n_489),
.B(n_481),
.Y(n_494)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_477),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_461),
.C(n_465),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_491),
.Y(n_495)
);

OA21x2_ASAP7_75t_SL g489 ( 
.A1(n_483),
.A2(n_472),
.B(n_466),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

AO21x1_ASAP7_75t_SL g497 ( 
.A1(n_493),
.A2(n_494),
.B(n_490),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_497),
.B1(n_495),
.B2(n_490),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_498),
.B(n_499),
.C(n_479),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_496),
.A2(n_488),
.B(n_487),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_475),
.C(n_13),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_501),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_502),
.A2(n_10),
.B(n_13),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_14),
.Y(n_504)
);


endmodule