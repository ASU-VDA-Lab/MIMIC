module real_jpeg_14994_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_215;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_53),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_8),
.A2(n_23),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_8),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_8),
.A2(n_23),
.B1(n_36),
.B2(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_47),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_8),
.B(n_56),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_37),
.C(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_8),
.B(n_118),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_8),
.B(n_82),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_8),
.A2(n_24),
.B(n_61),
.C(n_196),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_120)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_122),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_101),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_16),
.B(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_70),
.C(n_85),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_17),
.A2(n_18),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_18),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_45),
.CI(n_54),
.CON(n_18),
.SN(n_18)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_45),
.C(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_20),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_134)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.C(n_26),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_23),
.A2(n_58),
.B(n_62),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_24),
.A2(n_25),
.B1(n_61),
.B2(n_62),
.Y(n_69)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B(n_41),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_34),
.B(n_151),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_34),
.A2(n_44),
.B(n_117),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_44),
.B(n_72),
.Y(n_71)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_36),
.A2(n_37),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_37),
.B(n_171),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_41),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_41),
.B(n_182),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_44),
.B(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_44),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_48),
.B(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_67),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_56),
.A2(n_63),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_57),
.B(n_98),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_59),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_59),
.B(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_63),
.B(n_110),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_85),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_74),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_73),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_73),
.B(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_83),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_75),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_76),
.B(n_82),
.Y(n_203)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_78),
.B(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_78),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_82),
.B(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.C(n_96),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_100),
.B(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_121),
.B(n_166),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_141),
.B(n_218),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_126),
.B(n_129),
.Y(n_219)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_135),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_130),
.A2(n_131),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_135),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_139),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_136),
.B(n_138),
.CI(n_139),
.CON(n_208),
.SN(n_208)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_212),
.B(n_217),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_199),
.B(n_211),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_185),
.B(n_198),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_167),
.B(n_184),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_161),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_161),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_160),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_178),
.B(n_183),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_210),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.C(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);


endmodule