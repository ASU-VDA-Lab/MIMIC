module real_jpeg_104_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_305, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_305;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_286;
wire n_292;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_197;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_293;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_295;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_1),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_108),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_108),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_108),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_3),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_34),
.B1(n_63),
.B2(n_64),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_4),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_138),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_138),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_46),
.B1(n_63),
.B2(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_46),
.Y(n_145)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_168),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_168),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_168),
.Y(n_247)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_49),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_79),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_79),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_14),
.B(n_68),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_14),
.B(n_64),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_14),
.A2(n_57),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_14),
.B(n_26),
.C(n_42),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_159),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_87),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_30),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_14),
.B(n_50),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_14),
.A2(n_64),
.B(n_200),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_110),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_90),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_22),
.A2(n_23),
.B(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_23),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_23),
.A2(n_35),
.B1(n_52),
.B2(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_24),
.A2(n_144),
.B(n_146),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_24),
.A2(n_32),
.B(n_146),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_24),
.A2(n_29),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_25),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_25),
.A2(n_30),
.B1(n_145),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_25),
.A2(n_96),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_25),
.A2(n_30),
.B1(n_159),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_25),
.A2(n_30),
.B1(n_247),
.B2(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_26),
.B(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_29),
.B(n_32),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_29),
.A2(n_98),
.B(n_156),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_30),
.B(n_99),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_35),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_45),
.B(n_47),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_36),
.A2(n_45),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_36),
.A2(n_47),
.B(n_73),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_36),
.A2(n_102),
.B1(n_196),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_48),
.Y(n_75)
);

OAI21x1_ASAP7_75t_R g120 ( 
.A1(n_37),
.A2(n_50),
.B(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_37),
.A2(n_72),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_37),
.A2(n_50),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_37),
.A2(n_50),
.B1(n_233),
.B2(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_40),
.B1(n_83),
.B2(n_85),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_39),
.B(n_63),
.C(n_85),
.Y(n_201)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_40),
.A2(n_83),
.B(n_199),
.C(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_40),
.B(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_65),
.B(n_67),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_55),
.A2(n_62),
.B1(n_107),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_55),
.A2(n_62),
.B1(n_137),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_55),
.A2(n_62),
.B1(n_167),
.B2(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_58),
.B(n_159),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_58),
.B(n_61),
.C(n_64),
.Y(n_160)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_60),
.A2(n_63),
.B(n_158),
.C(n_160),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_62),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_64),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_70),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_76),
.B(n_89),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_75),
.A2(n_101),
.B(n_102),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_87),
.B2(n_88),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_86),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_80),
.A2(n_87),
.B1(n_163),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_81),
.A2(n_118),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_81),
.A2(n_86),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_81),
.A2(n_86),
.B1(n_187),
.B2(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_87),
.B(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_111),
.CI(n_112),
.CON(n_110),
.SN(n_110)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_90),
.A2(n_91),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_103),
.C(n_106),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_92),
.A2(n_93),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_103),
.B(n_106),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_110),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_122),
.B2(n_126),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_296),
.B(n_302),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_181),
.B(n_295),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_169),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_132),
.B(n_169),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_148),
.C(n_150),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_133),
.B(n_148),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_141),
.B2(n_142),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_143),
.B(n_147),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_150),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_161),
.C(n_166),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_151),
.A2(n_152),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_161),
.B(n_166),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_180),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_173),
.B(n_177),
.C(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI321xp33_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_276),
.A3(n_287),
.B1(n_293),
.B2(n_294),
.C(n_305),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_222),
.B(n_275),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_203),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_203),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_194),
.C(n_197),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_185),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_190),
.C(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_194),
.B(n_197),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_202),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_215),
.B2(n_216),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_204),
.B(n_217),
.C(n_220),
.Y(n_288)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_206),
.B(n_210),
.C(n_214),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_270),
.B(n_274),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_260),
.B(n_269),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_241),
.B(n_259),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_234),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_238),
.C(n_240),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_253),
.B(n_258),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_248),
.B(n_252),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_251),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_261),
.B(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_265),
.C(n_267),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_279),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_286),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_281),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_301),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);


endmodule