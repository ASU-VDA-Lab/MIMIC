module fake_jpeg_10717_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_1),
.B1(n_5),
.B2(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_2),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_6),
.B1(n_9),
.B2(n_14),
.Y(n_17)
);

AOI22x1_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_14),
.B1(n_10),
.B2(n_12),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_14),
.C(n_9),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_20),
.B1(n_15),
.B2(n_23),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.C(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_28),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_33),
.B(n_25),
.Y(n_37)
);


endmodule