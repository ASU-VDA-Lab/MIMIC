module fake_netlist_1_5837_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVxp33_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
AND2x2_ASAP7_75t_L g6 ( .A(n_5), .B(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_7), .B(n_4), .Y(n_8) );
AND4x1_ASAP7_75t_L g9 ( .A(n_8), .B(n_3), .C(n_1), .D(n_2), .Y(n_9) );
AO22x2_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_0), .B1(n_2), .B2(n_5), .Y(n_10) );
OAI21xp5_ASAP7_75t_SL g11 ( .A1(n_10), .A2(n_0), .B(n_9), .Y(n_11) );
endmodule