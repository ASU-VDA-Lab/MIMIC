module fake_jpeg_12933_n_286 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_46),
.B(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_68),
.Y(n_104)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_71),
.CON(n_79),
.SN(n_79)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_28),
.B(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_70),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_20),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_76),
.A2(n_78),
.B1(n_86),
.B2(n_87),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_22),
.C(n_25),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_12),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_31),
.B1(n_19),
.B2(n_42),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_79),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_42),
.B1(n_30),
.B2(n_19),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_30),
.B1(n_36),
.B2(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_44),
.B(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_85),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_30),
.B1(n_40),
.B2(n_32),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_91),
.A2(n_108),
.B(n_9),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_34),
.B1(n_40),
.B2(n_36),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_41),
.B1(n_38),
.B2(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_103),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_41),
.B1(n_38),
.B2(n_27),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_110),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_20),
.B1(n_29),
.B2(n_4),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_29),
.B(n_2),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_13),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_14),
.Y(n_122)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_138),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_2),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_123),
.Y(n_163)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_126),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_5),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_128),
.C(n_139),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_96),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_13),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_79),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_139),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_11),
.B(n_12),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_102),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_77),
.B(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_99),
.Y(n_164)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_84),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_123),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_98),
.B1(n_90),
.B2(n_76),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_162),
.B1(n_164),
.B2(n_116),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_165),
.C(n_127),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_90),
.B1(n_97),
.B2(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_99),
.C(n_101),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_117),
.A2(n_84),
.B1(n_109),
.B2(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_109),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_127),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_180),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_125),
.B1(n_116),
.B2(n_135),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_186),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_172),
.B1(n_163),
.B2(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_190),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_182),
.Y(n_218)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_137),
.B(n_134),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_206),
.B(n_123),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_155),
.B(n_121),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_132),
.B1(n_169),
.B2(n_175),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_130),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_205),
.B1(n_170),
.B2(n_125),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_151),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_161),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_131),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_160),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_204),
.B1(n_186),
.B2(n_183),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_214),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_163),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_151),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_165),
.C(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_119),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_220),
.B(n_191),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_128),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_162),
.B1(n_159),
.B2(n_173),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_173),
.B1(n_198),
.B2(n_196),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_141),
.B(n_136),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_241),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_222),
.A2(n_184),
.B1(n_189),
.B2(n_194),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_234),
.B(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_224),
.B1(n_226),
.B2(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_204),
.A3(n_187),
.B1(n_190),
.B2(n_193),
.C1(n_128),
.C2(n_118),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_232),
.B(n_237),
.Y(n_245)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_200),
.B(n_169),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_239),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_226),
.C(n_211),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_208),
.C(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_244),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_248),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_212),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_227),
.C(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_235),
.C(n_214),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_239),
.B1(n_249),
.B2(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_235),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_234),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_238),
.C(n_228),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_249),
.B(n_246),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_240),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_269),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_250),
.B1(n_243),
.B2(n_253),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_266),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_261),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_254),
.B(n_209),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_256),
.B(n_253),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_269),
.Y(n_276)
);

AOI31xp67_ASAP7_75t_SL g274 ( 
.A1(n_265),
.A2(n_259),
.A3(n_254),
.B(n_258),
.Y(n_274)
);

OAI321xp33_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_268),
.A3(n_267),
.B1(n_220),
.B2(n_233),
.C(n_120),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_279),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_270),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_271),
.B(n_273),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_278),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_283),
.B(n_115),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_146),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_124),
.Y(n_286)
);


endmodule