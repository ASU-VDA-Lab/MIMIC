module fake_aes_682_n_1306 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1306);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1306;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g291 ( .A(n_191), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_122), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_42), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_144), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_195), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_121), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_159), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_243), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_231), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_19), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_288), .Y(n_301) );
BUFx5_ASAP7_75t_L g302 ( .A(n_205), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_150), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_154), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_31), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_27), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_168), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_190), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_198), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_2), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_286), .Y(n_312) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_98), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_163), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_29), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_36), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_5), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_141), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_53), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_129), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_124), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_123), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_125), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_21), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_19), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_184), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_200), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_238), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_136), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_197), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_24), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_66), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_0), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_166), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_234), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_162), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_252), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_130), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_143), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_230), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_82), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_158), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_37), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_271), .Y(n_345) );
INVxp33_ASAP7_75t_SL g346 ( .A(n_282), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_100), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_253), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_274), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_217), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_46), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_46), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_213), .Y(n_353) );
BUFx8_ASAP7_75t_SL g354 ( .A(n_176), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_173), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_138), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_40), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_215), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_18), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_132), .Y(n_360) );
BUFx5_ASAP7_75t_L g361 ( .A(n_220), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_54), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_277), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_101), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_161), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_218), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_196), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_4), .Y(n_368) );
BUFx5_ASAP7_75t_L g369 ( .A(n_172), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_15), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_20), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_229), .B(n_64), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_110), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_55), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_211), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_284), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_28), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_108), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_186), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_174), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_179), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_41), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_152), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_105), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_208), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_242), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_104), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_232), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_2), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_24), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_51), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_137), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_31), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_226), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_228), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_212), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_12), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_5), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_262), .Y(n_399) );
CKINVDCx14_ASAP7_75t_R g400 ( .A(n_107), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_40), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_272), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_207), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_287), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_140), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_9), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_155), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_97), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_149), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_169), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_49), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_280), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_32), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_78), .B(n_93), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_214), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_257), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_28), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_146), .Y(n_418) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_15), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_95), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_139), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_273), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_11), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_261), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_42), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_210), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_11), .B(n_34), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_89), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_44), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_34), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_164), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_160), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_114), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_127), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_335), .B(n_0), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_382), .B(n_1), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_348), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_335), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_348), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_300), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_298), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_355), .B(n_1), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_298), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_367), .B(n_3), .Y(n_444) );
BUFx10_ASAP7_75t_L g445 ( .A(n_292), .Y(n_445) );
AND2x2_ASAP7_75t_R g446 ( .A(n_344), .B(n_3), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_298), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_300), .B(n_4), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_311), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_311), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_386), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_358), .B(n_6), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_298), .Y(n_453) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_385), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_319), .B(n_6), .Y(n_455) );
INVx6_ASAP7_75t_L g456 ( .A(n_302), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_304), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_423), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_354), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_319), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_293), .Y(n_461) );
BUFx8_ASAP7_75t_L g462 ( .A(n_302), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_400), .B(n_7), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_352), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_352), .B(n_7), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_291), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_304), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_305), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_460), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_435), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_437), .B(n_428), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_462), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_441), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_437), .B(n_428), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_439), .B(n_368), .C(n_334), .Y(n_477) );
BUFx10_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_456), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_455), .B(n_357), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_441), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_466), .B(n_400), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_456), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_455), .A2(n_419), .B1(n_357), .B2(n_340), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_461), .B(n_436), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_441), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_456), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_451), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_456), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_466), .B(n_371), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_462), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_448), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_451), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g496 ( .A(n_463), .B(n_372), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_462), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_459), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_448), .A2(n_315), .B1(n_316), .B2(n_306), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_448), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_457), .B(n_390), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_443), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_465), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_438), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_443), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_459), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_438), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_463), .B(n_419), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_468), .B(n_313), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_478), .B(n_445), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_506), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_498), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_478), .B(n_445), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_492), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_478), .B(n_457), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_506), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_478), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_511), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_492), .B(n_442), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_506), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_514), .B(n_445), .Y(n_526) );
OR2x6_ASAP7_75t_L g527 ( .A(n_473), .B(n_446), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_470), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_514), .B(n_467), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_469), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_506), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_503), .A2(n_468), .B1(n_449), .B2(n_450), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_511), .Y(n_533) );
BUFx4f_ASAP7_75t_L g534 ( .A(n_473), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_486), .B(n_468), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_486), .B(n_444), .Y(n_536) );
BUFx4f_ASAP7_75t_L g537 ( .A(n_496), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_483), .B(n_452), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_512), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_503), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_492), .B(n_294), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_503), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_497), .B(n_464), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_469), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_503), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_497), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_472), .B(n_432), .Y(n_547) );
NAND3xp33_ASAP7_75t_SL g548 ( .A(n_494), .B(n_458), .C(n_349), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_469), .Y(n_549) );
INVx4_ASAP7_75t_L g550 ( .A(n_497), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_469), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_505), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_505), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_476), .B(n_432), .Y(n_555) );
AO22x1_ASAP7_75t_L g556 ( .A1(n_510), .A2(n_346), .B1(n_331), .B2(n_313), .Y(n_556) );
INVx5_ASAP7_75t_L g557 ( .A(n_512), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_489), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_491), .B(n_440), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_481), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_481), .B(n_398), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_493), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
NAND3xp33_ASAP7_75t_SL g566 ( .A(n_485), .B(n_378), .C(n_329), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_471), .A2(n_347), .B(n_331), .Y(n_567) );
BUFx3_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_496), .A2(n_383), .B1(n_413), .B2(n_401), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_512), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_513), .B(n_440), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_479), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_501), .B(n_449), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_513), .B(n_450), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_493), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_471), .B(n_295), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_474), .B(n_296), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_512), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_500), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_504), .A2(n_324), .B1(n_326), .B2(n_317), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_485), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_504), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_477), .B(n_347), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_474), .B(n_301), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_499), .B(n_332), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_479), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_484), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_484), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_488), .B(n_297), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_488), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_490), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_490), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_482), .B(n_303), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_482), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_495), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_475), .Y(n_597) );
AND2x6_ASAP7_75t_SL g598 ( .A(n_475), .B(n_427), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_495), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_502), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_502), .B(n_351), .Y(n_601) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_546), .B(n_299), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_520), .A2(n_363), .B(n_309), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_554), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_550), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_536), .B(n_359), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_520), .A2(n_363), .B(n_312), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_530), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_530), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_528), .Y(n_611) );
BUFx5_ASAP7_75t_L g612 ( .A(n_522), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_554), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_582), .A2(n_377), .B(n_389), .C(n_370), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_589), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_561), .B(n_391), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_544), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_544), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_538), .A2(n_314), .B(n_308), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_519), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_549), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_536), .B(n_393), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_546), .B(n_327), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_559), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_550), .B(n_330), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_549), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_540), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_567), .A2(n_320), .B(n_318), .Y(n_628) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_568), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_519), .B(n_362), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_517), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_585), .A2(n_323), .B(n_322), .Y(n_632) );
BUFx3_ASAP7_75t_L g633 ( .A(n_568), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_551), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_542), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_535), .B(n_397), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_585), .A2(n_328), .B(n_325), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_519), .Y(n_638) );
INVx4_ASAP7_75t_L g639 ( .A(n_537), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_563), .B(n_406), .Y(n_640) );
BUFx3_ASAP7_75t_L g641 ( .A(n_537), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_580), .A2(n_417), .B1(n_425), .B2(n_411), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_573), .A2(n_430), .B(n_429), .C(n_338), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_569), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_545), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_580), .A2(n_337), .B1(n_342), .B2(n_339), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_526), .A2(n_345), .B(n_343), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_571), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_551), .A2(n_553), .B(n_552), .Y(n_649) );
BUFx3_ASAP7_75t_L g650 ( .A(n_565), .Y(n_650) );
OR2x6_ASAP7_75t_L g651 ( .A(n_527), .B(n_350), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_527), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_573), .A2(n_364), .B(n_366), .C(n_353), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_574), .B(n_333), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_553), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_564), .A2(n_375), .B(n_373), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_570), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_562), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_527), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_562), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_575), .A2(n_379), .B(n_376), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_579), .A2(n_394), .B(n_387), .Y(n_664) );
BUFx4f_ASAP7_75t_L g665 ( .A(n_543), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_570), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_570), .Y(n_667) );
O2A1O1Ixp5_ASAP7_75t_L g668 ( .A1(n_524), .A2(n_414), .B(n_307), .C(n_321), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_583), .A2(n_396), .B(n_395), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_586), .B(n_399), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_543), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_570), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_547), .B(n_360), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_581), .A2(n_404), .B1(n_405), .B2(n_402), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_SL g675 ( .A1(n_584), .A2(n_414), .B(n_508), .C(n_307), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_529), .Y(n_676) );
INVx5_ASAP7_75t_L g677 ( .A(n_598), .Y(n_677) );
BUFx3_ASAP7_75t_L g678 ( .A(n_565), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_578), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_586), .A2(n_408), .B1(n_409), .B2(n_407), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_578), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_548), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_555), .A2(n_412), .B(n_416), .C(n_410), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_515), .A2(n_420), .B1(n_421), .B2(n_418), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_534), .Y(n_685) );
AO221x1_ASAP7_75t_L g686 ( .A1(n_566), .A2(n_385), .B1(n_434), .B2(n_433), .C(n_422), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_560), .A2(n_431), .B(n_321), .C(n_341), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_581), .B(n_374), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_518), .B(n_381), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_524), .A2(n_341), .B(n_310), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_523), .Y(n_691) );
INVx4_ASAP7_75t_L g692 ( .A(n_539), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_541), .A2(n_356), .B(n_310), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_556), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_534), .B(n_403), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_541), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_539), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_576), .A2(n_384), .B(n_356), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_532), .A2(n_415), .B1(n_426), .B2(n_424), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_539), .B(n_365), .Y(n_700) );
INVx4_ASAP7_75t_L g701 ( .A(n_557), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_533), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_578), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_577), .B(n_380), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_557), .B(n_392), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_601), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_558), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_532), .A2(n_384), .B1(n_336), .B2(n_388), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_578), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_584), .A2(n_388), .B(n_336), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_572), .B(n_8), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_557), .B(n_302), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_558), .Y(n_713) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_587), .A2(n_385), .B1(n_9), .B2(n_10), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_572), .A2(n_302), .B1(n_361), .B2(n_369), .Y(n_715) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_557), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_590), .B(n_8), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_558), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_593), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_588), .A2(n_508), .B(n_480), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_592), .A2(n_480), .B(n_475), .Y(n_721) );
INVx2_ASAP7_75t_SL g722 ( .A(n_558), .Y(n_722) );
AO32x2_ASAP7_75t_L g723 ( .A1(n_591), .A2(n_302), .A3(n_361), .B1(n_369), .B2(n_443), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_516), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_591), .Y(n_725) );
NAND2x2_ASAP7_75t_L g726 ( .A(n_594), .B(n_10), .Y(n_726) );
AOI222xp33_ASAP7_75t_L g727 ( .A1(n_648), .A2(n_516), .B1(n_531), .B2(n_525), .C1(n_521), .C2(n_594), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_676), .B(n_521), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_691), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_721), .A2(n_531), .B(n_525), .Y(n_730) );
CKINVDCx11_ASAP7_75t_R g731 ( .A(n_611), .Y(n_731) );
NAND2x1p5_ASAP7_75t_L g732 ( .A(n_639), .B(n_597), .Y(n_732) );
OAI21x1_ASAP7_75t_L g733 ( .A1(n_720), .A2(n_599), .B(n_595), .Y(n_733) );
OAI21x1_ASAP7_75t_L g734 ( .A1(n_649), .A2(n_599), .B(n_595), .Y(n_734) );
AO21x2_ASAP7_75t_L g735 ( .A1(n_675), .A2(n_596), .B(n_600), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_639), .B(n_596), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_702), .Y(n_737) );
OAI21x1_ASAP7_75t_L g738 ( .A1(n_649), .A2(n_600), .B(n_597), .Y(n_738) );
BUFx12f_ASAP7_75t_L g739 ( .A(n_631), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_711), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_641), .B(n_12), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_659), .Y(n_742) );
AO31x2_ASAP7_75t_L g743 ( .A1(n_653), .A2(n_453), .A3(n_443), .B(n_447), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_659), .Y(n_744) );
OA21x2_ASAP7_75t_L g745 ( .A1(n_668), .A2(n_597), .B(n_361), .Y(n_745) );
OAI21x1_ASAP7_75t_L g746 ( .A1(n_712), .A2(n_597), .B(n_361), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_719), .Y(n_747) );
OAI222xp33_ASAP7_75t_L g748 ( .A1(n_651), .A2(n_13), .B1(n_14), .B2(n_16), .C1(n_17), .C2(n_18), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_633), .B(n_13), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_624), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_615), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_706), .Y(n_752) );
OR2x6_ASAP7_75t_L g753 ( .A(n_651), .B(n_385), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g754 ( .A1(n_614), .A2(n_453), .B(n_447), .C(n_454), .Y(n_754) );
BUFx3_ASAP7_75t_L g755 ( .A(n_677), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_692), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_647), .A2(n_480), .B(n_475), .Y(n_757) );
AO21x2_ASAP7_75t_L g758 ( .A1(n_698), .A2(n_361), .B(n_302), .Y(n_758) );
OAI21x1_ASAP7_75t_L g759 ( .A1(n_690), .A2(n_369), .B(n_361), .Y(n_759) );
OA21x2_ASAP7_75t_L g760 ( .A1(n_693), .A2(n_369), .B(n_447), .Y(n_760) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_606), .A2(n_369), .B(n_57), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_606), .A2(n_369), .B(n_58), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_629), .B(n_14), .Y(n_763) );
AO21x2_ASAP7_75t_L g764 ( .A1(n_710), .A2(n_686), .B(n_619), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_671), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_692), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_644), .A2(n_16), .B1(n_17), .B2(n_20), .Y(n_767) );
AOI21x1_ASAP7_75t_L g768 ( .A1(n_700), .A2(n_453), .B(n_447), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_636), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_694), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_670), .B(n_21), .Y(n_771) );
INVx1_ASAP7_75t_SL g772 ( .A(n_659), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_651), .B(n_22), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_670), .A2(n_640), .B1(n_674), .B2(n_654), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_643), .A2(n_447), .B1(n_453), .B2(n_454), .C(n_26), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_665), .B(n_22), .Y(n_776) );
OAI21x1_ASAP7_75t_L g777 ( .A1(n_634), .A2(n_59), .B(n_56), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_628), .A2(n_454), .B(n_453), .Y(n_778) );
OAI21x1_ASAP7_75t_L g779 ( .A1(n_656), .A2(n_61), .B(n_60), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_677), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_628), .A2(n_454), .B(n_475), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_657), .A2(n_63), .B(n_62), .Y(n_782) );
BUFx12f_ASAP7_75t_L g783 ( .A(n_682), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_636), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_627), .A2(n_454), .B(n_475), .Y(n_785) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_726), .Y(n_786) );
OA21x2_ASAP7_75t_L g787 ( .A1(n_715), .A2(n_487), .B(n_480), .Y(n_787) );
OAI21x1_ASAP7_75t_L g788 ( .A1(n_660), .A2(n_67), .B(n_65), .Y(n_788) );
OAI21x1_ASAP7_75t_L g789 ( .A1(n_662), .A2(n_69), .B(n_68), .Y(n_789) );
AOI21x1_ASAP7_75t_L g790 ( .A1(n_705), .A2(n_487), .B(n_480), .Y(n_790) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_661), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_677), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g793 ( .A(n_665), .B(n_23), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_685), .B(n_23), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g795 ( .A1(n_635), .A2(n_487), .B(n_480), .Y(n_795) );
INVxp67_ASAP7_75t_L g796 ( .A(n_616), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_701), .B(n_25), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_680), .A2(n_509), .B1(n_487), .B2(n_27), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_607), .B(n_25), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_666), .A2(n_71), .B(n_70), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_622), .A2(n_674), .B1(n_683), .B2(n_714), .C(n_673), .Y(n_801) );
OAI22x1_ASAP7_75t_L g802 ( .A1(n_652), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_704), .B(n_30), .Y(n_803) );
INVx5_ASAP7_75t_L g804 ( .A(n_716), .Y(n_804) );
OA21x2_ASAP7_75t_L g805 ( .A1(n_604), .A2(n_509), .B(n_487), .Y(n_805) );
INVx4_ASAP7_75t_L g806 ( .A(n_716), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_667), .Y(n_807) );
INVx3_ASAP7_75t_L g808 ( .A(n_701), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_667), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_642), .B(n_688), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_642), .A2(n_509), .B1(n_487), .B2(n_35), .Y(n_811) );
AND2x4_ASAP7_75t_L g812 ( .A(n_716), .B(n_32), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_687), .A2(n_663), .B(n_658), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_667), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_645), .Y(n_815) );
OA21x2_ASAP7_75t_L g816 ( .A1(n_608), .A2(n_509), .B(n_73), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_714), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_696), .B(n_33), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_646), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_724), .Y(n_820) );
OA21x2_ASAP7_75t_L g821 ( .A1(n_632), .A2(n_509), .B(n_74), .Y(n_821) );
NAND2x1p5_ASAP7_75t_L g822 ( .A(n_650), .B(n_33), .Y(n_822) );
OAI21x1_ASAP7_75t_L g823 ( .A1(n_672), .A2(n_75), .B(n_72), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_725), .A2(n_509), .B1(n_36), .B2(n_37), .Y(n_824) );
OAI21x1_ASAP7_75t_L g825 ( .A1(n_679), .A2(n_177), .B(n_285), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_695), .B(n_35), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_664), .B(n_38), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_684), .B(n_38), .Y(n_828) );
OAI21x1_ASAP7_75t_L g829 ( .A1(n_681), .A2(n_178), .B(n_283), .Y(n_829) );
INVxp67_ASAP7_75t_L g830 ( .A(n_699), .Y(n_830) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_717), .B(n_39), .C(n_41), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_703), .A2(n_180), .B(n_281), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g833 ( .A(n_678), .B(n_39), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_625), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_669), .B(n_43), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_689), .B(n_43), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_709), .A2(n_181), .B(n_279), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_605), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_708), .A2(n_44), .B1(n_45), .B2(n_47), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_655), .A2(n_45), .B1(n_47), .B2(n_48), .Y(n_840) );
BUFx12f_ASAP7_75t_L g841 ( .A(n_602), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_655), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_613), .B(n_48), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_697), .B(n_49), .Y(n_844) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_602), .Y(n_845) );
BUFx8_ASAP7_75t_L g846 ( .A(n_723), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_621), .B(n_50), .Y(n_847) );
CKINVDCx16_ASAP7_75t_R g848 ( .A(n_602), .Y(n_848) );
OAI21x1_ASAP7_75t_L g849 ( .A1(n_697), .A2(n_183), .B(n_278), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_723), .B(n_50), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_626), .B(n_51), .Y(n_851) );
INVx4_ASAP7_75t_L g852 ( .A(n_620), .Y(n_852) );
BUFx2_ASAP7_75t_L g853 ( .A(n_707), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_609), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_610), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g856 ( .A1(n_603), .A2(n_185), .B(n_276), .Y(n_856) );
NAND2x1p5_ASAP7_75t_L g857 ( .A(n_620), .B(n_52), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_617), .A2(n_52), .B1(n_53), .B2(n_76), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_718), .A2(n_77), .B1(n_79), .B2(n_80), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_618), .Y(n_860) );
INVxp67_ASAP7_75t_L g861 ( .A(n_623), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_637), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_817), .A2(n_630), .B1(n_713), .B2(n_612), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_801), .A2(n_612), .B1(n_722), .B2(n_638), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_774), .B(n_718), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_729), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_796), .B(n_723), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_750), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_801), .A2(n_612), .B1(n_638), .B2(n_620), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_774), .A2(n_612), .B1(n_638), .B2(n_84), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_751), .B(n_612), .Y(n_871) );
CKINVDCx10_ASAP7_75t_R g872 ( .A(n_731), .Y(n_872) );
INVx3_ASAP7_75t_L g873 ( .A(n_841), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_753), .A2(n_81), .B1(n_83), .B2(n_85), .Y(n_874) );
OAI22xp5_ASAP7_75t_SL g875 ( .A1(n_793), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_739), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_753), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_753), .A2(n_94), .B1(n_96), .B2(n_99), .Y(n_878) );
A2O1A1Ixp33_ASAP7_75t_L g879 ( .A1(n_803), .A2(n_102), .B(n_103), .C(n_106), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_769), .A2(n_109), .B1(n_111), .B2(n_112), .C(n_113), .Y(n_880) );
AOI21xp33_ASAP7_75t_L g881 ( .A1(n_830), .A2(n_290), .B(n_116), .Y(n_881) );
OAI322xp33_ASAP7_75t_L g882 ( .A1(n_773), .A2(n_115), .A3(n_117), .B1(n_118), .B2(n_119), .C1(n_120), .C2(n_126), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_737), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_810), .B(n_275), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_763), .A2(n_128), .B1(n_131), .B2(n_133), .Y(n_885) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_750), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_747), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_757), .A2(n_134), .B(n_135), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_822), .A2(n_142), .B1(n_145), .B2(n_147), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_752), .Y(n_890) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_833), .A2(n_148), .B1(n_151), .B2(n_153), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_815), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_819), .B(n_270), .Y(n_893) );
AO21x2_ASAP7_75t_L g894 ( .A1(n_778), .A2(n_156), .B(n_157), .Y(n_894) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_795), .A2(n_165), .B(n_167), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_741), .B(n_170), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_828), .A2(n_171), .B1(n_175), .B2(n_182), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_820), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_784), .B(n_187), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_794), .A2(n_188), .B1(n_189), .B2(n_192), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_794), .A2(n_193), .B1(n_194), .B2(n_199), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_763), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_902) );
AO21x2_ASAP7_75t_L g903 ( .A1(n_778), .A2(n_204), .B(n_206), .Y(n_903) );
A2O1A1Ixp33_ASAP7_75t_L g904 ( .A1(n_831), .A2(n_209), .B(n_216), .C(n_219), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_765), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_818), .A2(n_221), .B1(n_222), .B2(n_223), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_851), .A2(n_224), .B1(n_225), .B2(n_227), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_771), .A2(n_233), .B1(n_235), .B2(n_236), .C(n_237), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_791), .B(n_239), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_740), .A2(n_240), .B1(n_241), .B2(n_244), .C(n_245), .Y(n_910) );
AO21x2_ASAP7_75t_L g911 ( .A1(n_781), .A2(n_246), .B(n_248), .Y(n_911) );
OAI21xp5_ASAP7_75t_L g912 ( .A1(n_781), .A2(n_249), .B(n_250), .Y(n_912) );
A2O1A1Ixp33_ASAP7_75t_L g913 ( .A1(n_831), .A2(n_251), .B(n_254), .C(n_255), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_728), .Y(n_914) );
OAI21xp33_ASAP7_75t_L g915 ( .A1(n_799), .A2(n_256), .B(n_258), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_741), .A2(n_259), .B1(n_260), .B2(n_263), .Y(n_916) );
AOI33xp33_ASAP7_75t_L g917 ( .A1(n_767), .A2(n_264), .A3(n_265), .B1(n_266), .B2(n_267), .B3(n_268), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_728), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_799), .A2(n_269), .B(n_827), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_804), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_736), .B(n_771), .Y(n_921) );
AO31x2_ASAP7_75t_L g922 ( .A1(n_811), .A2(n_824), .A3(n_798), .B(n_859), .Y(n_922) );
BUFx6f_ASAP7_75t_L g923 ( .A(n_804), .Y(n_923) );
INVx4_ASAP7_75t_L g924 ( .A(n_804), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_749), .B(n_776), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_786), .Y(n_926) );
OA21x2_ASAP7_75t_L g927 ( .A1(n_738), .A2(n_759), .B(n_730), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_749), .A2(n_811), .B1(n_797), .B2(n_839), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_836), .A2(n_826), .B1(n_827), .B2(n_835), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_839), .A2(n_848), .B1(n_862), .B2(n_835), .Y(n_930) );
OAI221xp5_ASAP7_75t_L g931 ( .A1(n_861), .A2(n_775), .B1(n_780), .B2(n_792), .C(n_755), .Y(n_931) );
OA21x2_ASAP7_75t_L g932 ( .A1(n_761), .A2(n_762), .B(n_746), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_842), .B(n_853), .Y(n_933) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_846), .A2(n_812), .B1(n_824), .B2(n_775), .Y(n_934) );
OAI21xp33_ASAP7_75t_L g935 ( .A1(n_798), .A2(n_840), .B(n_858), .Y(n_935) );
AOI21xp33_ASAP7_75t_L g936 ( .A1(n_813), .A2(n_727), .B(n_764), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_736), .B(n_770), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_838), .B(n_860), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_854), .B(n_812), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g940 ( .A(n_806), .B(n_766), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_843), .A2(n_847), .B1(n_727), .B2(n_754), .C(n_857), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g942 ( .A1(n_748), .A2(n_802), .B1(n_847), .B2(n_843), .C(n_834), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_756), .A2(n_808), .B1(n_766), .B2(n_850), .Y(n_943) );
NAND3xp33_ASAP7_75t_L g944 ( .A(n_846), .B(n_859), .C(n_745), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_844), .A2(n_808), .B(n_756), .C(n_856), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_813), .B(n_855), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_783), .Y(n_947) );
AO22x1_ASAP7_75t_L g948 ( .A1(n_806), .A2(n_852), .B1(n_772), .B2(n_845), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_743), .Y(n_949) );
OAI21xp5_ASAP7_75t_L g950 ( .A1(n_734), .A2(n_795), .B(n_785), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_764), .B(n_772), .Y(n_951) );
OAI21x1_ASAP7_75t_L g952 ( .A1(n_790), .A2(n_733), .B(n_768), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g953 ( .A1(n_785), .A2(n_732), .B1(n_745), .B2(n_805), .C(n_814), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_758), .A2(n_735), .B1(n_852), .B2(n_807), .Y(n_954) );
OAI211xp5_ASAP7_75t_SL g955 ( .A1(n_742), .A2(n_809), .B(n_744), .C(n_743), .Y(n_955) );
A2O1A1Ixp33_ASAP7_75t_L g956 ( .A1(n_849), .A2(n_782), .B(n_789), .C(n_788), .Y(n_956) );
NAND2xp5_ASAP7_75t_SL g957 ( .A(n_845), .B(n_779), .Y(n_957) );
OR2x6_ASAP7_75t_L g958 ( .A(n_845), .B(n_777), .Y(n_958) );
OAI21x1_ASAP7_75t_L g959 ( .A1(n_787), .A2(n_837), .B(n_832), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_821), .A2(n_816), .B1(n_787), .B2(n_805), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_758), .B(n_735), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_760), .B(n_816), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_800), .Y(n_963) );
INVx3_ASAP7_75t_L g964 ( .A(n_823), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_760), .A2(n_821), .B1(n_825), .B2(n_829), .Y(n_965) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_774), .A2(n_796), .B1(n_801), .B2(n_528), .C(n_817), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_757), .A2(n_795), .B(n_781), .Y(n_967) );
BUFx12f_ASAP7_75t_L g968 ( .A(n_731), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_729), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_738), .A2(n_730), .B(n_746), .Y(n_970) );
AOI21xp5_ASAP7_75t_L g971 ( .A1(n_757), .A2(n_795), .B(n_781), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_729), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_729), .Y(n_973) );
OR2x6_ASAP7_75t_L g974 ( .A(n_753), .B(n_639), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_729), .Y(n_975) );
AOI21xp5_ASAP7_75t_L g976 ( .A1(n_757), .A2(n_795), .B(n_781), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_817), .A2(n_527), .B1(n_801), .B2(n_566), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_817), .A2(n_527), .B1(n_801), .B2(n_566), .Y(n_978) );
OR2x2_ASAP7_75t_L g979 ( .A(n_750), .B(n_528), .Y(n_979) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_774), .A2(n_796), .B1(n_801), .B2(n_528), .C(n_817), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_796), .A2(n_640), .B1(n_536), .B2(n_582), .C(n_817), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g982 ( .A1(n_757), .A2(n_795), .B(n_781), .Y(n_982) );
CKINVDCx10_ASAP7_75t_R g983 ( .A(n_731), .Y(n_983) );
AO21x2_ASAP7_75t_L g984 ( .A1(n_778), .A2(n_781), .B(n_738), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_914), .B(n_918), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_892), .B(n_969), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_925), .B(n_865), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_946), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_866), .Y(n_989) );
NOR2x1p5_ASAP7_75t_L g990 ( .A(n_944), .B(n_924), .Y(n_990) );
AND2x4_ASAP7_75t_SL g991 ( .A(n_974), .B(n_924), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_979), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_966), .B(n_980), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_883), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_928), .B(n_921), .Y(n_995) );
BUFx3_ASAP7_75t_L g996 ( .A(n_923), .Y(n_996) );
INVx2_ASAP7_75t_L g997 ( .A(n_927), .Y(n_997) );
BUFx6f_ASAP7_75t_L g998 ( .A(n_923), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_887), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_973), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_972), .B(n_975), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_949), .Y(n_1002) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_977), .B(n_978), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_981), .B(n_890), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_905), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_938), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_932), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_932), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_898), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_942), .B(n_929), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_867), .B(n_864), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_934), .B(n_939), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_868), .B(n_886), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_970), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_920), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_893), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_964), .Y(n_1017) );
BUFx3_ASAP7_75t_L g1018 ( .A(n_923), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_930), .B(n_933), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_896), .B(n_919), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_955), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_919), .B(n_869), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_961), .Y(n_1023) );
BUFx6f_ASAP7_75t_L g1024 ( .A(n_952), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_871), .B(n_922), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_963), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_922), .B(n_884), .Y(n_1027) );
BUFx12f_ASAP7_75t_SL g1028 ( .A(n_974), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_964), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_943), .B(n_922), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_974), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_959), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_912), .B(n_940), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_937), .B(n_931), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_912), .B(n_899), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_917), .B(n_916), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_936), .B(n_954), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_951), .B(n_948), .Y(n_1038) );
HB1xp67_ASAP7_75t_L g1039 ( .A(n_873), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_962), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_894), .B(n_903), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_953), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_894), .B(n_903), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_873), .B(n_935), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_902), .B(n_901), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_900), .B(n_911), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_911), .B(n_863), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_944), .B(n_984), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_885), .B(n_870), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_875), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_907), .B(n_945), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_950), .B(n_904), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_909), .B(n_876), .Y(n_1053) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_968), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_958), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_957), .Y(n_1056) );
AOI21xp5_ASAP7_75t_L g1057 ( .A1(n_956), .A2(n_976), .B(n_967), .Y(n_1057) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_947), .Y(n_1058) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_926), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_875), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_889), .B(n_891), .Y(n_1061) );
BUFx3_ASAP7_75t_L g1062 ( .A(n_872), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_913), .B(n_897), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_983), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_960), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_941), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_908), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_879), .B(n_910), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_882), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_880), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_882), .Y(n_1071) );
INVxp67_ASAP7_75t_L g1072 ( .A(n_874), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_971), .Y(n_1073) );
AND2x4_ASAP7_75t_L g1074 ( .A(n_888), .B(n_895), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_906), .B(n_881), .Y(n_1075) );
AND2x4_ASAP7_75t_SL g1076 ( .A(n_965), .B(n_877), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_982), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_878), .B(n_915), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_914), .B(n_918), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_914), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_946), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1025), .B(n_1040), .Y(n_1082) );
INVx4_ASAP7_75t_L g1083 ( .A(n_991), .Y(n_1083) );
INVxp67_ASAP7_75t_SL g1084 ( .A(n_1079), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_990), .B(n_1023), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_1010), .A2(n_1003), .B1(n_993), .B2(n_1004), .C(n_1060), .Y(n_1086) );
INVx5_ASAP7_75t_L g1087 ( .A(n_998), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_1034), .A2(n_1060), .B1(n_1050), .B2(n_1044), .C(n_1072), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1025), .B(n_1040), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1006), .B(n_986), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1009), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1023), .B(n_985), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_1066), .A2(n_1006), .B1(n_992), .B2(n_1005), .C(n_1000), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1080), .B(n_1027), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1080), .B(n_1027), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1096 ( .A1(n_1034), .A2(n_1019), .B1(n_1066), .B2(n_1053), .C(n_1061), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_1015), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_997), .Y(n_1098) );
AO21x2_ASAP7_75t_L g1099 ( .A1(n_1057), .A2(n_1077), .B(n_1073), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_997), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1013), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1011), .B(n_1001), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1001), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1002), .Y(n_1104) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_988), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1026), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_987), .B(n_995), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_987), .B(n_995), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_989), .Y(n_1109) );
OAI21x1_ASAP7_75t_L g1110 ( .A1(n_1032), .A2(n_1008), .B(n_1007), .Y(n_1110) );
OAI21xp5_ASAP7_75t_SL g1111 ( .A1(n_991), .A2(n_1031), .B(n_1064), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_989), .B(n_994), .Y(n_1112) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_1038), .Y(n_1113) );
INVxp33_ASAP7_75t_L g1114 ( .A(n_998), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1011), .B(n_988), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_994), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1019), .B(n_1081), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_999), .Y(n_1118) );
NAND2x1p5_ASAP7_75t_SL g1119 ( .A(n_1036), .B(n_1051), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_999), .Y(n_1120) );
NAND2xp33_ASAP7_75t_L g1121 ( .A(n_990), .B(n_1069), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1000), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1005), .B(n_1030), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1039), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_1069), .A2(n_1071), .B1(n_1020), .B2(n_1031), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_1012), .A2(n_1020), .B1(n_1070), .B2(n_1071), .Y(n_1126) );
NAND3xp33_ASAP7_75t_SL g1127 ( .A(n_1036), .B(n_1068), .C(n_1012), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1016), .B(n_996), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1037), .B(n_1065), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1042), .B(n_1038), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1037), .B(n_1065), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1042), .B(n_1077), .Y(n_1132) );
INVx5_ASAP7_75t_L g1133 ( .A(n_998), .Y(n_1133) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_1018), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1022), .B(n_1073), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1021), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1022), .B(n_1055), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1021), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1055), .B(n_1052), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1052), .B(n_1033), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1028), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_1016), .A2(n_1070), .B1(n_1051), .B2(n_1067), .C(n_1033), .Y(n_1142) );
BUFx3_ASAP7_75t_L g1143 ( .A(n_1058), .Y(n_1143) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_1028), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1047), .B(n_1046), .Y(n_1145) );
NOR2x1_ASAP7_75t_L g1146 ( .A(n_1111), .B(n_1062), .Y(n_1146) );
NAND4xp25_ASAP7_75t_L g1147 ( .A(n_1086), .B(n_1062), .C(n_1054), .D(n_1059), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1091), .Y(n_1148) );
INVx2_ASAP7_75t_SL g1149 ( .A(n_1087), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1085), .B(n_1056), .Y(n_1150) );
OAI21xp5_ASAP7_75t_SL g1151 ( .A1(n_1127), .A2(n_1035), .B(n_1076), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1098), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1109), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1116), .Y(n_1154) );
AND2x4_ASAP7_75t_L g1155 ( .A(n_1085), .B(n_1017), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1082), .B(n_1048), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1082), .B(n_1048), .Y(n_1157) );
NOR3xp33_ASAP7_75t_L g1158 ( .A(n_1136), .B(n_1054), .C(n_1067), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1103), .B(n_1035), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1089), .B(n_1047), .Y(n_1160) );
NAND2xp5_ASAP7_75t_SL g1161 ( .A(n_1093), .B(n_1041), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1102), .B(n_1059), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_1096), .A2(n_1049), .B1(n_1045), .B2(n_1068), .Y(n_1163) );
NAND2x1p5_ASAP7_75t_L g1164 ( .A(n_1083), .B(n_1058), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1118), .Y(n_1165) );
A2O1A1Ixp33_ASAP7_75t_SL g1166 ( .A1(n_1138), .A2(n_1088), .B(n_1124), .C(n_1121), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_1142), .A2(n_1049), .B1(n_1045), .B2(n_1063), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1120), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1107), .B(n_1063), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1122), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1112), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1097), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1101), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_1143), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1100), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1140), .B(n_1029), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1102), .B(n_1107), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1140), .B(n_1029), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1108), .B(n_1076), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1108), .B(n_1014), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1092), .B(n_1046), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1094), .B(n_1043), .Y(n_1182) );
AOI22xp33_ASAP7_75t_SL g1183 ( .A1(n_1144), .A2(n_1078), .B1(n_1041), .B2(n_1043), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1104), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1092), .B(n_1078), .Y(n_1185) );
NAND2xp5_ASAP7_75t_SL g1186 ( .A(n_1083), .B(n_1024), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1143), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1084), .B(n_1024), .Y(n_1188) );
NOR2xp33_ASAP7_75t_SL g1189 ( .A(n_1083), .B(n_1144), .Y(n_1189) );
OA21x2_ASAP7_75t_L g1190 ( .A1(n_1110), .A2(n_1074), .B(n_1075), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1106), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1095), .B(n_1074), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1115), .B(n_1074), .Y(n_1193) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1105), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1145), .B(n_1075), .Y(n_1195) );
INVxp67_ASAP7_75t_L g1196 ( .A(n_1172), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1160), .B(n_1182), .Y(n_1197) );
INVxp67_ASAP7_75t_L g1198 ( .A(n_1194), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1152), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1177), .B(n_1113), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1184), .Y(n_1201) );
INVx1_ASAP7_75t_SL g1202 ( .A(n_1174), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1160), .B(n_1145), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1182), .B(n_1137), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1156), .B(n_1137), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1156), .B(n_1113), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1157), .B(n_1135), .Y(n_1207) );
NOR2x1_ASAP7_75t_R g1208 ( .A(n_1174), .B(n_1134), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1157), .B(n_1135), .Y(n_1209) );
NOR3xp33_ASAP7_75t_SL g1210 ( .A(n_1147), .B(n_1125), .C(n_1128), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1173), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1191), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1169), .B(n_1185), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1169), .B(n_1129), .Y(n_1214) );
NAND2xp5_ASAP7_75t_SL g1215 ( .A(n_1189), .B(n_1141), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1148), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1193), .B(n_1139), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1153), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1154), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1195), .B(n_1129), .Y(n_1220) );
AND5x1_ASAP7_75t_L g1221 ( .A(n_1166), .B(n_1119), .C(n_1121), .D(n_1126), .E(n_1130), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1165), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1168), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1170), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1180), .Y(n_1225) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_1188), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1227 ( .A1(n_1163), .A2(n_1131), .B1(n_1117), .B2(n_1123), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1195), .B(n_1131), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1192), .B(n_1123), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1181), .B(n_1115), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1175), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1207), .B(n_1171), .Y(n_1232) );
INVx1_ASAP7_75t_SL g1233 ( .A(n_1202), .Y(n_1233) );
AOI32xp33_ASAP7_75t_L g1234 ( .A1(n_1197), .A2(n_1146), .A3(n_1187), .B1(n_1158), .B2(n_1163), .Y(n_1234) );
INVx1_ASAP7_75t_SL g1235 ( .A(n_1200), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1197), .B(n_1192), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1223), .Y(n_1237) );
AND2x4_ASAP7_75t_L g1238 ( .A(n_1226), .B(n_1150), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1207), .B(n_1176), .Y(n_1239) );
AOI22xp5_ASAP7_75t_L g1240 ( .A1(n_1227), .A2(n_1151), .B1(n_1167), .B2(n_1183), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1223), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1224), .Y(n_1242) );
INVx4_ASAP7_75t_L g1243 ( .A(n_1208), .Y(n_1243) );
AOI21xp5_ASAP7_75t_L g1244 ( .A1(n_1215), .A2(n_1166), .B(n_1186), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1224), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1210), .A2(n_1167), .B1(n_1164), .B2(n_1162), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1198), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1209), .B(n_1178), .Y(n_1248) );
AOI211x1_ASAP7_75t_L g1249 ( .A1(n_1213), .A2(n_1161), .B(n_1159), .C(n_1090), .Y(n_1249) );
CKINVDCx14_ASAP7_75t_R g1250 ( .A(n_1200), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1209), .B(n_1178), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1205), .B(n_1176), .Y(n_1252) );
NAND3xp33_ASAP7_75t_SL g1253 ( .A(n_1196), .B(n_1164), .C(n_1186), .Y(n_1253) );
AND2x4_ASAP7_75t_L g1254 ( .A(n_1225), .B(n_1150), .Y(n_1254) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1199), .Y(n_1255) );
NAND3xp33_ASAP7_75t_L g1256 ( .A(n_1211), .B(n_1161), .C(n_1190), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1216), .Y(n_1257) );
INVx2_ASAP7_75t_L g1258 ( .A(n_1199), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1247), .Y(n_1259) );
OAI21x1_ASAP7_75t_SL g1260 ( .A1(n_1243), .A2(n_1230), .B(n_1228), .Y(n_1260) );
AOI21xp33_ASAP7_75t_L g1261 ( .A1(n_1234), .A2(n_1132), .B(n_1149), .Y(n_1261) );
NAND2xp5_ASAP7_75t_SL g1262 ( .A(n_1243), .B(n_1206), .Y(n_1262) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1255), .Y(n_1263) );
INVxp67_ASAP7_75t_SL g1264 ( .A(n_1247), .Y(n_1264) );
A2O1A1Ixp33_ASAP7_75t_L g1265 ( .A1(n_1250), .A2(n_1206), .B(n_1204), .C(n_1217), .Y(n_1265) );
INVxp67_ASAP7_75t_L g1266 ( .A(n_1233), .Y(n_1266) );
XNOR2x1_ASAP7_75t_L g1267 ( .A(n_1240), .B(n_1179), .Y(n_1267) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_1249), .B(n_1218), .C(n_1219), .Y(n_1268) );
OAI22xp33_ASAP7_75t_L g1269 ( .A1(n_1253), .A2(n_1214), .B1(n_1117), .B2(n_1220), .Y(n_1269) );
NAND2xp5_ASAP7_75t_SL g1270 ( .A(n_1256), .B(n_1222), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1235), .B(n_1204), .Y(n_1271) );
AOI32xp33_ASAP7_75t_L g1272 ( .A1(n_1246), .A2(n_1203), .A3(n_1229), .B1(n_1205), .B2(n_1150), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1251), .B(n_1229), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1237), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1241), .Y(n_1275) );
INVx1_ASAP7_75t_SL g1276 ( .A(n_1238), .Y(n_1276) );
OAI21xp33_ASAP7_75t_L g1277 ( .A1(n_1272), .A2(n_1254), .B(n_1238), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1264), .Y(n_1278) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_1265), .A2(n_1238), .B1(n_1244), .B2(n_1239), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1262), .B(n_1232), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1259), .Y(n_1281) );
NAND2x1_ASAP7_75t_L g1282 ( .A(n_1260), .B(n_1254), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1274), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1275), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1268), .B(n_1252), .Y(n_1285) );
A2O1A1Ixp33_ASAP7_75t_SL g1286 ( .A1(n_1261), .A2(n_1257), .B(n_1258), .C(n_1255), .Y(n_1286) );
AOI21xp5_ASAP7_75t_L g1287 ( .A1(n_1269), .A2(n_1231), .B(n_1258), .Y(n_1287) );
NAND4xp25_ASAP7_75t_L g1288 ( .A(n_1279), .B(n_1277), .C(n_1286), .D(n_1287), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1278), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1290 ( .A(n_1280), .B(n_1266), .Y(n_1290) );
O2A1O1Ixp33_ASAP7_75t_L g1291 ( .A1(n_1285), .A2(n_1270), .B(n_1276), .C(n_1271), .Y(n_1291) );
AOI211xp5_ASAP7_75t_L g1292 ( .A1(n_1287), .A2(n_1254), .B(n_1242), .C(n_1245), .Y(n_1292) );
INVxp67_ASAP7_75t_L g1293 ( .A(n_1281), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_1282), .A2(n_1267), .B1(n_1273), .B2(n_1248), .Y(n_1294) );
AOI221xp5_ASAP7_75t_L g1295 ( .A1(n_1288), .A2(n_1284), .B1(n_1283), .B2(n_1119), .C(n_1263), .Y(n_1295) );
NOR2x1_ASAP7_75t_R g1296 ( .A(n_1289), .B(n_1087), .Y(n_1296) );
NAND2x1p5_ASAP7_75t_L g1297 ( .A(n_1290), .B(n_1087), .Y(n_1297) );
AND2x4_ASAP7_75t_L g1298 ( .A(n_1293), .B(n_1236), .Y(n_1298) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_1295), .A2(n_1294), .B1(n_1292), .B2(n_1291), .Y(n_1299) );
NAND3xp33_ASAP7_75t_SL g1300 ( .A(n_1297), .B(n_1221), .C(n_1132), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g1301 ( .A1(n_1299), .A2(n_1298), .B1(n_1296), .B2(n_1212), .Y(n_1301) );
OAI22xp5_ASAP7_75t_SL g1302 ( .A1(n_1301), .A2(n_1300), .B1(n_1087), .B2(n_1133), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1302), .Y(n_1303) );
AOI21xp33_ASAP7_75t_SL g1304 ( .A1(n_1303), .A2(n_1190), .B(n_1201), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_1304), .A2(n_1201), .B1(n_1155), .B2(n_1099), .Y(n_1305) );
AOI21xp5_ASAP7_75t_L g1306 ( .A1(n_1305), .A2(n_1106), .B(n_1114), .Y(n_1306) );
endmodule