module fake_jpeg_19174_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_39),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_40),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_68),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_71),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_39),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_85),
.Y(n_94)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_80),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_41),
.B1(n_42),
.B2(n_29),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_38),
.B1(n_53),
.B2(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_41),
.B1(n_17),
.B2(n_20),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_81),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_24),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_16),
.B1(n_21),
.B2(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_16),
.B1(n_26),
.B2(n_18),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_49),
.Y(n_114)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_55),
.B1(n_43),
.B2(n_31),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_115),
.B1(n_61),
.B2(n_113),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_49),
.C(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_114),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_49),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_80),
.B(n_78),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_82),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_62),
.A2(n_55),
.B1(n_43),
.B2(n_34),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_115),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_64),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_123),
.B1(n_128),
.B2(n_130),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_85),
.B1(n_77),
.B2(n_64),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_131),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_86),
.B1(n_72),
.B2(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_118),
.B1(n_108),
.B2(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_109),
.B(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_114),
.B1(n_117),
.B2(n_102),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_69),
.B1(n_88),
.B2(n_89),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_55),
.B1(n_71),
.B2(n_69),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_97),
.B(n_95),
.C(n_30),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_90),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_109),
.B1(n_105),
.B2(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_146),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_111),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_95),
.B1(n_97),
.B2(n_88),
.Y(n_147)
);

OAI22x1_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_145),
.B1(n_139),
.B2(n_136),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_100),
.C(n_120),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_172),
.C(n_143),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_108),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_144),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_163),
.B(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_98),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_116),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_107),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_170),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_34),
.B(n_18),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_87),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_173),
.B(n_122),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_33),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_191),
.B(n_195),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_121),
.B1(n_122),
.B2(n_142),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_188),
.B1(n_193),
.B2(n_194),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_133),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_196),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_177),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_132),
.B1(n_138),
.B2(n_141),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_135),
.B(n_134),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_166),
.B(n_183),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_145),
.B1(n_139),
.B2(n_136),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_136),
.B1(n_95),
.B2(n_25),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_30),
.C(n_25),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_25),
.B1(n_22),
.B2(n_33),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_198),
.B1(n_173),
.B2(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_195),
.B1(n_179),
.B2(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_187),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_207),
.C(n_211),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_161),
.C(n_154),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_157),
.B1(n_173),
.B2(n_168),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_185),
.B(n_164),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_175),
.A2(n_174),
.B(n_153),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_216),
.B1(n_203),
.B2(n_199),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_174),
.B(n_172),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_189),
.Y(n_224)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_215),
.A2(n_182),
.B1(n_184),
.B2(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_231),
.B1(n_200),
.B2(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_189),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_226),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_232),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_212),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_196),
.C(n_192),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_229),
.C(n_22),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_176),
.B1(n_188),
.B2(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_176),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_8),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_194),
.C(n_198),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_22),
.B1(n_9),
.B2(n_15),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_235),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_204),
.B(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_28),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_243),
.B1(n_236),
.B2(n_238),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_218),
.B1(n_225),
.B2(n_230),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_8),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_8),
.C(n_14),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_245),
.C(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_224),
.C(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_235),
.C(n_244),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_222),
.B(n_9),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_245),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_7),
.C(n_12),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_9),
.B(n_15),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_262),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_260),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_247),
.A3(n_246),
.B1(n_6),
.B2(n_11),
.C1(n_12),
.C2(n_5),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_259),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_234),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_240),
.B(n_7),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_247),
.B(n_12),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_1),
.B(n_3),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_246),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_260),
.C(n_255),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_272),
.B(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_267),
.C(n_266),
.Y(n_275)
);

AOI221xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_276),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_1),
.B(n_3),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_4),
.B(n_5),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_4),
.Y(n_279)
);


endmodule