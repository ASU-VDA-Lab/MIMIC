module fake_jpeg_17267_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_15),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_13),
.B(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_15),
.C(n_12),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_17),
.B(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_15),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_23),
.Y(n_44)
);

AOI32xp33_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_17),
.A3(n_14),
.B1(n_9),
.B2(n_13),
.Y(n_36)
);

FAx1_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_37),
.CI(n_39),
.CON(n_51),
.SN(n_51)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_43),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_50),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_37),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_35),
.C(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_48),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_53),
.B(n_55),
.C(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_11),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_64),
.B1(n_46),
.B2(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_0),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_73),
.C(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_7),
.Y(n_77)
);


endmodule