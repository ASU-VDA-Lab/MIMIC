module fake_netlist_1_802_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_2), .B(n_1), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
INVx3_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
AND2x4_ASAP7_75t_SL g7 ( .A(n_5), .B(n_4), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
OAI22xp33_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_6), .B1(n_4), .B2(n_2), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_1), .Y(n_10) );
O2A1O1Ixp33_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_8), .B(n_7), .C(n_2), .Y(n_11) );
AND4x1_ASAP7_75t_SL g12 ( .A(n_10), .B(n_0), .C(n_2), .D(n_3), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
NOR2x1_ASAP7_75t_L g14 ( .A(n_11), .B(n_0), .Y(n_14) );
OAI31xp33_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_0), .A3(n_12), .B(n_14), .Y(n_15) );
NAND2x1p5_ASAP7_75t_L g16 ( .A(n_15), .B(n_0), .Y(n_16) );
endmodule