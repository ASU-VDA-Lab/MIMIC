module real_jpeg_30270_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_0),
.Y(n_405)
);

BUFx12f_ASAP7_75t_L g540 ( 
.A(n_0),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_1),
.B(n_61),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_1),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_1),
.B(n_290),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_1),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_1),
.B(n_403),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_2),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_3),
.B(n_333),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_3),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_3),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_3),
.B(n_353),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_3),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_3),
.B(n_403),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_4),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_4),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g413 ( 
.A(n_4),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_4),
.B(n_154),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_4),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_186),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_5),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_5),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_5),
.B(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_6),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_8),
.Y(n_543)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_9),
.Y(n_291)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_9),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g277 ( 
.A(n_10),
.B(n_278),
.Y(n_277)
);

NAND2x1_ASAP7_75t_L g337 ( 
.A(n_10),
.B(n_31),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_10),
.B(n_365),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_10),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_10),
.B(n_506),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_10),
.B(n_542),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_10),
.B(n_549),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_11),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_11),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_11),
.B(n_162),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_11),
.B(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_11),
.B(n_174),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_11),
.B(n_555),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_11),
.B(n_563),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_12),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_12),
.B(n_89),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_13),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_13),
.B(n_198),
.Y(n_197)
);

NAND2x1_ASAP7_75t_SL g222 ( 
.A(n_13),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_158),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_14),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_15),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_15),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_15),
.B(n_131),
.Y(n_130)
);

NAND2x1_ASAP7_75t_L g153 ( 
.A(n_15),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_15),
.B(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_16),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_16),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_17),
.B(n_203),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g263 ( 
.A(n_17),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_17),
.B(n_293),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_17),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_17),
.B(n_468),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_17),
.B(n_511),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_17),
.B(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_17),
.B(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_19),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_19),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_19),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_19),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_19),
.B(n_198),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_19),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_19),
.B(n_403),
.Y(n_402)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_91),
.B(n_593),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_88),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_22),
.B(n_89),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_86),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI221xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.C(n_56),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.C(n_50),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_32),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_32),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_32),
.Y(n_265)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_32),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_39),
.Y(n_180)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_44),
.B1(n_60),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_64),
.C(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_53),
.Y(n_166)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_53),
.Y(n_357)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_83),
.C(n_84),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_57),
.B(n_83),
.CI(n_84),
.CON(n_141),
.SN(n_141)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_70),
.C(n_76),
.Y(n_57)
);

XNOR2x1_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_60),
.A2(n_77),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_62),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_63),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_77),
.C(n_80),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_76),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_123),
.C(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_77),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_77),
.A2(n_129),
.B1(n_130),
.B2(n_139),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_79),
.Y(n_270)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_91),
.A2(n_594),
.B(n_595),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_142),
.B(n_592),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_141),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_94),
.B(n_141),
.Y(n_592)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_119),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_95),
.B(n_97),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_111),
.C(n_115),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.C(n_106),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_99),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_107),
.Y(n_233)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_105),
.Y(n_365)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_109),
.Y(n_472)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_110),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.Y(n_121)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_119),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_135),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g306 ( 
.A(n_120),
.B(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_122),
.A2(n_136),
.B1(n_137),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_122),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_212),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_129),
.B(n_207),
.C(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_129),
.A2(n_130),
.B1(n_153),
.B2(n_207),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_134),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g596 ( 
.A(n_141),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_316),
.B(n_587),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_312),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_300),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_244),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_SL g589 ( 
.A(n_146),
.B(n_244),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_209),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_147),
.B(n_210),
.C(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_167),
.C(n_181),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_150),
.B(n_167),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_152),
.B(n_161),
.C(n_165),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_157),
.B1(n_201),
.B2(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_155),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_155),
.Y(n_491)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_155),
.Y(n_519)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_157),
.A2(n_197),
.B1(n_201),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_168),
.C(n_176),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_161),
.B(n_177),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_164),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_168),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_169),
.B(n_170),
.Y(n_274)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_173),
.B(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_182),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.C(n_205),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_183),
.B(n_196),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_188),
.C(n_191),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_187),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_193),
.B(n_340),
.Y(n_487)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_195),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.C(n_202),
.Y(n_196)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_200),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_205),
.B(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_230),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_211),
.B(n_214),
.C(n_217),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_226),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_235),
.B(n_236),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_235),
.B(n_236),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_237),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_R g244 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_248),
.Y(n_377)
);

XNOR2x2_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_252),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_275),
.C(n_297),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.C(n_273),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_254),
.B(n_258),
.C(n_273),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_258),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_266),
.B(n_271),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_263),
.B(n_272),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_266),
.Y(n_418)
);

INVx3_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_273),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_298),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_286),
.B(n_296),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.C(n_284),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_SL g370 ( 
.A(n_277),
.B(n_281),
.C(n_284),
.Y(n_370)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_281),
.A2(n_284),
.B1(n_285),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_292),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_287),
.B(n_292),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_287),
.B(n_292),
.Y(n_371)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_291),
.Y(n_416)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_291),
.Y(n_512)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_300),
.A2(n_589),
.B(n_590),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_301),
.B(n_303),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.C(n_309),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_312),
.A2(n_588),
.B(n_591),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_313),
.B(n_314),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_426),
.B(n_584),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_378),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_318),
.A2(n_585),
.B(n_586),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_375),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g586 ( 
.A(n_319),
.B(n_375),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.C(n_373),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_321),
.B(n_373),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_324),
.B(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_348),
.C(n_366),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_382),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.C(n_342),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_327),
.B(n_329),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_330),
.A2(n_331),
.B1(n_342),
.B2(n_343),
.Y(n_453)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_335),
.B(n_338),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_393),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_SL g338 ( 
.A1(n_333),
.A2(n_339),
.B(n_341),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_335),
.A2(n_336),
.B1(n_341),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OA21x2_ASAP7_75t_SL g437 ( 
.A1(n_343),
.A2(n_344),
.B(n_347),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_367),
.B1(n_368),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_359),
.C(n_363),
.Y(n_349)
);

XOR2x1_ASAP7_75t_L g422 ( 
.A(n_350),
.B(n_423),
.Y(n_422)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.C(n_358),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_351),
.A2(n_352),
.B1(n_358),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_354),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_356),
.B(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_359),
.A2(n_360),
.B1(n_363),
.B2(n_364),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_424),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_379),
.B(n_424),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.C(n_389),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_381),
.B(n_385),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_417),
.C(n_420),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_390),
.A2(n_391),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.C(n_406),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_392),
.B(n_476),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_395),
.A2(n_406),
.B1(n_407),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_396),
.A2(n_397),
.B1(n_401),
.B2(n_402),
.Y(n_473)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_412),
.C(n_413),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_408),
.A2(n_409),
.B1(n_413),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_412),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_417),
.A2(n_421),
.B1(n_422),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_480),
.B(n_582),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_454),
.B(n_457),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_428),
.B(n_454),
.C(n_583),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_433),
.C(n_450),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_429),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_451),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.C(n_438),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_437),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_460),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_444),
.C(n_446),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_439),
.B(n_496),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_440),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_486)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_444),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_496)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_449),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_478),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_458),
.B(n_478),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.C(n_474),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_498),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_475),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.C(n_473),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_473),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.C(n_470),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_466),
.B(n_470),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_467),
.B(n_531),
.Y(n_530)
);

INVx3_ASAP7_75t_SL g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_472),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_499),
.B(n_581),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_497),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_482),
.B(n_497),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.C(n_495),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_483),
.B(n_579),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_485),
.B(n_495),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.C(n_488),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_486),
.B(n_487),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_488),
.B(n_525),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_492),
.Y(n_488)
);

AO22x1_ASAP7_75t_L g521 ( 
.A1(n_489),
.A2(n_490),
.B1(n_492),
.B2(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_576),
.B(n_580),
.Y(n_499)
);

OAI21x1_ASAP7_75t_SL g500 ( 
.A1(n_501),
.A2(n_533),
.B(n_575),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_522),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_522),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_515),
.C(n_521),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_503),
.A2(n_504),
.B1(n_571),
.B2(n_573),
.Y(n_570)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_509),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_528),
.C(n_529),
.Y(n_527)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_513),
.Y(n_509)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_510),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_513),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_515),
.A2(n_516),
.B1(n_521),
.B2(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_520),
.Y(n_551)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_521),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_523),
.A2(n_524),
.B1(n_526),
.B2(n_532),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_523),
.B(n_527),
.C(n_530),
.Y(n_577)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_526),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_534),
.A2(n_568),
.B(n_574),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_535),
.A2(n_552),
.B(n_567),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_544),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_536),
.B(n_544),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_537),
.B(n_541),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_541),
.Y(n_560)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_541),
.B(n_562),
.Y(n_561)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_551),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_546),
.A2(n_547),
.B1(n_548),
.B2(n_550),
.Y(n_545)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_546),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_547),
.B(n_550),
.C(n_551),
.Y(n_569)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_553),
.A2(n_561),
.B(n_566),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_560),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_560),
.Y(n_566)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx3_ASAP7_75t_SL g563 ( 
.A(n_564),
.Y(n_563)
);

INVx8_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_570),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_569),
.B(n_570),
.Y(n_574)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_571),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g576 ( 
.A(n_577),
.B(n_578),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_577),
.B(n_578),
.Y(n_580)
);


endmodule