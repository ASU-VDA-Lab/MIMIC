module fake_ariane_2398_n_68 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_68);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_68;

wire n_66;
wire n_56;
wire n_60;
wire n_24;
wire n_22;
wire n_43;
wire n_49;
wire n_27;
wire n_20;
wire n_48;
wire n_29;
wire n_64;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_62;
wire n_47;
wire n_18;
wire n_32;
wire n_28;
wire n_58;
wire n_37;
wire n_65;
wire n_51;
wire n_67;
wire n_45;
wire n_34;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_33;
wire n_44;
wire n_19;
wire n_30;
wire n_40;
wire n_39;
wire n_59;
wire n_31;
wire n_42;
wire n_57;
wire n_63;
wire n_53;
wire n_21;
wire n_23;
wire n_61;
wire n_35;
wire n_54;
wire n_25;

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_7),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_5),
.B1(n_1),
.B2(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AND2x6_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_18),
.B(n_24),
.Y(n_38)
);

AO31x2_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_20),
.A3(n_21),
.B(n_30),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_30),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_27),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_32),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AO21x2_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_28),
.B(n_23),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_26),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_39),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_39),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_43),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_43),
.Y(n_54)
);

OAI31xp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_36),
.A3(n_43),
.B(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_50),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_22),
.B1(n_25),
.B2(n_19),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_37),
.Y(n_61)
);

OAI211xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_2),
.B(n_4),
.C(n_6),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_59),
.B(n_57),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_19),
.C(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_64),
.B1(n_62),
.B2(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_37),
.B1(n_14),
.B2(n_16),
.Y(n_68)
);


endmodule