module fake_jpeg_1092_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_544;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_8),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_22),
.C(n_30),
.Y(n_138)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_28),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_109),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_9),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_33),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_101),
.B(n_117),
.Y(n_144)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_33),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_112),
.Y(n_141)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_16),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_38),
.B(n_16),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_34),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

BUFx12f_ASAP7_75t_SL g117 ( 
.A(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_38),
.B(n_15),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_32),
.Y(n_152)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_124),
.A2(n_21),
.B(n_48),
.Y(n_191)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_57),
.B1(n_40),
.B2(n_59),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_127),
.A2(n_173),
.B1(n_182),
.B2(n_200),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_138),
.B(n_10),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_63),
.A2(n_22),
.B1(n_30),
.B2(n_32),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_140),
.A2(n_201),
.B1(n_179),
.B2(n_185),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_150),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_152),
.B(n_160),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_109),
.B(n_35),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_159),
.B(n_89),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_28),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_61),
.B(n_35),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_175),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_92),
.A2(n_57),
.B1(n_59),
.B2(n_39),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_56),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_75),
.B(n_55),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_178),
.B(n_181),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_69),
.B(n_56),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_64),
.A2(n_48),
.B1(n_55),
.B2(n_36),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_93),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_65),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_197),
.B(n_0),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_122),
.B(n_36),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

HAxp5_ASAP7_75t_SL g197 ( 
.A(n_117),
.B(n_21),
.CON(n_197),
.SN(n_197)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_125),
.B(n_59),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_67),
.A2(n_78),
.B1(n_116),
.B2(n_113),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_105),
.A2(n_31),
.B1(n_57),
.B2(n_21),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_102),
.A2(n_57),
.B1(n_31),
.B2(n_10),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_204),
.B1(n_106),
.B2(n_96),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_84),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_209),
.Y(n_295)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_153),
.B1(n_108),
.B2(n_119),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_213),
.Y(n_332)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_215),
.Y(n_310)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_216),
.Y(n_315)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_218),
.Y(n_328)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_220),
.Y(n_335)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_145),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_221),
.Y(n_343)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_222),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_227),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_228),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_133),
.A2(n_94),
.B1(n_120),
.B2(n_121),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_226),
.A2(n_229),
.B(n_249),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_169),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_180),
.B(n_80),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_230),
.A2(n_242),
.B1(n_272),
.B2(n_283),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_180),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_232),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_141),
.B(n_122),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_144),
.B(n_74),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_234),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_192),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_235),
.B(n_236),
.Y(n_317)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_238),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_182),
.A2(n_114),
.B(n_97),
.C(n_107),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g313 ( 
.A1(n_240),
.A2(n_148),
.B1(n_158),
.B2(n_2),
.Y(n_313)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_123),
.B1(n_103),
.B2(n_98),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_129),
.B1(n_202),
.B2(n_127),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_243),
.A2(n_245),
.B1(n_268),
.B2(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_130),
.Y(n_244)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_140),
.A2(n_91),
.B1(n_90),
.B2(n_86),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

AND2x4_ASAP7_75t_SL g249 ( 
.A(n_198),
.B(n_0),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_157),
.Y(n_252)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_259),
.Y(n_320)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_136),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_260),
.B(n_265),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_161),
.Y(n_261)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_139),
.Y(n_262)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_186),
.Y(n_263)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_172),
.Y(n_264)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_151),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_170),
.B(n_13),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_270),
.Y(n_341)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_126),
.Y(n_267)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_168),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_134),
.B(n_13),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_132),
.Y(n_271)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_155),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_143),
.Y(n_274)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_135),
.B(n_0),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_275),
.B(n_276),
.Y(n_345)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_168),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_136),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_277),
.B(n_278),
.Y(n_342)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_149),
.A2(n_15),
.B1(n_11),
.B2(n_2),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_281),
.Y(n_347)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_156),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_142),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_282),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_173),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_210),
.B(n_250),
.C(n_234),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_284),
.B(n_297),
.C(n_300),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_219),
.A2(n_205),
.B1(n_147),
.B2(n_148),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_285),
.A2(n_293),
.B1(n_306),
.B2(n_337),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_147),
.B1(n_187),
.B2(n_176),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_137),
.C(n_165),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_165),
.C(n_205),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_228),
.A2(n_223),
.B1(n_249),
.B2(n_239),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_187),
.B1(n_176),
.B2(n_167),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_164),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_308),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_167),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_158),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_327),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_240),
.B(n_276),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g323 ( 
.A1(n_226),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_323),
.A2(n_309),
.B1(n_306),
.B2(n_285),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_236),
.B(n_1),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_225),
.B(n_3),
.C(n_4),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_262),
.C(n_241),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_249),
.B(n_225),
.CI(n_233),
.CON(n_334),
.SN(n_334)
);

MAJIxp5_ASAP7_75t_SL g356 ( 
.A(n_334),
.B(n_302),
.C(n_287),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_279),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_229),
.A2(n_3),
.B(n_5),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_347),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_353),
.Y(n_400)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_341),
.B(n_217),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_350),
.B(n_372),
.Y(n_399)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_351),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_352),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_329),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_214),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_385),
.C(n_286),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_304),
.Y(n_420)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

AOI21x1_ASAP7_75t_L g360 ( 
.A1(n_303),
.A2(n_271),
.B(n_267),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_360),
.A2(n_310),
.B(n_325),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_376),
.B1(n_389),
.B2(n_393),
.Y(n_412)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_289),
.Y(n_362)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_365),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_320),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_292),
.B(n_312),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_366),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_280),
.B1(n_278),
.B2(n_238),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_369),
.B1(n_386),
.B2(n_388),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_332),
.A2(n_237),
.B1(n_222),
.B2(n_216),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_290),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_319),
.B(n_317),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_379),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_375),
.B(n_374),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_301),
.A2(n_212),
.B1(n_256),
.B2(n_246),
.Y(n_376)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_377),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_336),
.A2(n_264),
.B1(n_211),
.B2(n_221),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_378),
.A2(n_391),
.B1(n_394),
.B2(n_397),
.Y(n_432)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_296),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_387),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_311),
.B(n_248),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_381),
.B(n_383),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_302),
.B(n_327),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_302),
.B(n_258),
.C(n_209),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_345),
.A2(n_220),
.B1(n_218),
.B2(n_263),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_208),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_345),
.A2(n_259),
.B1(n_257),
.B2(n_277),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_307),
.A2(n_269),
.B1(n_255),
.B2(n_6),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_326),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_392),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_308),
.A2(n_215),
.B1(n_5),
.B2(n_6),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_345),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_303),
.A2(n_313),
.B1(n_334),
.B2(n_291),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_323),
.A2(n_300),
.B1(n_313),
.B2(n_297),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_396),
.Y(n_404)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_313),
.A2(n_286),
.B1(n_346),
.B2(n_342),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_349),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_401),
.B(n_422),
.C(n_439),
.Y(n_480)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_340),
.B(n_334),
.C(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_407),
.B(n_385),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_409),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_364),
.A2(n_304),
.B(n_305),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_410),
.A2(n_417),
.B(n_433),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_364),
.A2(n_360),
.B(n_395),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_393),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_423),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_420),
.B(n_430),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_318),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_425),
.Y(n_467)
);

BUFx24_ASAP7_75t_SL g423 ( 
.A(n_350),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_318),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_377),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_441),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_354),
.B(n_339),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_374),
.B(n_322),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_352),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_348),
.A2(n_316),
.B(n_305),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_353),
.A2(n_383),
.B(n_375),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_388),
.B(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_368),
.B(n_325),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_436),
.B(n_380),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_368),
.B(n_316),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_440),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_338),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_299),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_373),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_396),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_351),
.Y(n_465)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_444),
.A2(n_427),
.B(n_418),
.C(n_443),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_445),
.B(n_448),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_437),
.B(n_421),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_446),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_425),
.B(n_379),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_473),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_440),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_450),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_408),
.A2(n_355),
.B1(n_389),
.B2(n_367),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_452),
.A2(n_461),
.B1(n_471),
.B2(n_472),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_438),
.B(n_392),
.Y(n_454)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_414),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_456),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_411),
.A2(n_358),
.B1(n_370),
.B2(n_357),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_457),
.A2(n_343),
.B1(n_328),
.B2(n_321),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_414),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_459),
.Y(n_509)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_460),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_408),
.A2(n_404),
.B1(n_417),
.B2(n_412),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_404),
.A2(n_369),
.B1(n_386),
.B2(n_390),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_462),
.A2(n_475),
.B1(n_478),
.B2(n_411),
.Y(n_489)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_464),
.Y(n_498)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_469),
.B(n_470),
.Y(n_512)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_428),
.A2(n_363),
.B1(n_362),
.B2(n_344),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_398),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_422),
.B(n_299),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_431),
.C(n_401),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_400),
.B(n_294),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_474),
.B(n_479),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_432),
.A2(n_288),
.B1(n_371),
.B2(n_290),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_424),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_476),
.A2(n_477),
.B1(n_429),
.B2(n_441),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_412),
.A2(n_371),
.B1(n_288),
.B2(n_344),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_419),
.A2(n_335),
.B1(n_298),
.B2(n_295),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_399),
.B(n_335),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_493),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_484),
.B(n_466),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_461),
.A2(n_434),
.B1(n_400),
.B2(n_428),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_487),
.A2(n_508),
.B1(n_513),
.B2(n_509),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_489),
.A2(n_499),
.B1(n_501),
.B2(n_510),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_439),
.C(n_420),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_490),
.B(n_503),
.C(n_504),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_430),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_407),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_502),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_458),
.A2(n_433),
.B1(n_407),
.B2(n_403),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_458),
.A2(n_403),
.B1(n_424),
.B2(n_435),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_449),
.B(n_410),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_409),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_416),
.C(n_402),
.Y(n_504)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_450),
.A2(n_402),
.B1(n_416),
.B2(n_405),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_451),
.A2(n_399),
.B1(n_418),
.B2(n_405),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_454),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_445),
.A2(n_415),
.B1(n_413),
.B2(n_298),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_466),
.B(n_415),
.C(n_413),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_444),
.C(n_460),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_451),
.A2(n_294),
.B1(n_295),
.B2(n_328),
.Y(n_515)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_515),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_517),
.A2(n_457),
.B(n_453),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_518),
.A2(n_537),
.B1(n_548),
.B2(n_486),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_512),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_522),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_497),
.A2(n_481),
.B(n_447),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_521),
.A2(n_542),
.B(n_544),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_487),
.B(n_476),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_523),
.B(n_546),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_525),
.B(n_503),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_500),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_527),
.B(n_529),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_507),
.B(n_474),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_494),
.Y(n_530)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_530),
.Y(n_559)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_494),
.Y(n_531)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_531),
.Y(n_562)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_496),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_532),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_448),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_533),
.Y(n_551)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_496),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_534),
.Y(n_555)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_492),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_541),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_504),
.B(n_446),
.Y(n_539)
);

NOR3xp33_ASAP7_75t_SL g549 ( 
.A(n_539),
.B(n_485),
.C(n_467),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_483),
.C(n_490),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_540),
.B(n_543),
.C(n_501),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_484),
.B(n_463),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_491),
.B(n_479),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_514),
.B(n_455),
.C(n_468),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_516),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_545),
.A2(n_453),
.B1(n_508),
.B2(n_498),
.Y(n_570)
);

FAx1_ASAP7_75t_SL g546 ( 
.A(n_495),
.B(n_467),
.CI(n_468),
.CON(n_546),
.SN(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_455),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_547),
.B(n_471),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_509),
.B(n_469),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_554),
.Y(n_575)
);

MAJx2_ASAP7_75t_L g586 ( 
.A(n_552),
.B(n_561),
.C(n_569),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_544),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_528),
.B(n_540),
.C(n_524),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_556),
.B(n_558),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_511),
.C(n_499),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_524),
.B(n_488),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_520),
.A2(n_518),
.B1(n_536),
.B2(n_489),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_563),
.A2(n_475),
.B1(n_459),
.B2(n_477),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_505),
.C(n_486),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_564),
.B(n_566),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_541),
.B(n_505),
.C(n_456),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_568),
.B(n_573),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_492),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_570),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_535),
.B(n_525),
.C(n_547),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_482),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_535),
.B(n_485),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_526),
.B1(n_537),
.B2(n_533),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_574),
.B(n_584),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_SL g576 ( 
.A(n_552),
.B(n_523),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_576),
.B(n_589),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_L g577 ( 
.A(n_550),
.B(n_534),
.C(n_532),
.Y(n_577)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_577),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_551),
.A2(n_526),
.B1(n_521),
.B2(n_519),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_578),
.B(n_583),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_579),
.B(n_593),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_558),
.A2(n_545),
.B(n_513),
.Y(n_582)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_582),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_557),
.A2(n_564),
.B1(n_561),
.B2(n_566),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_498),
.C(n_545),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_590),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_554),
.B(n_472),
.C(n_465),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_565),
.B(n_546),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_570),
.A2(n_546),
.B1(n_452),
.B2(n_462),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_565),
.B(n_464),
.C(n_470),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_573),
.B(n_516),
.C(n_478),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_591),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_569),
.C(n_571),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_SL g620 ( 
.A(n_595),
.B(n_597),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_585),
.B(n_568),
.C(n_567),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_588),
.B(n_559),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_599),
.B(n_610),
.Y(n_613)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_600),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_592),
.B(n_567),
.C(n_560),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_602),
.B(n_333),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_586),
.B(n_591),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_606),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_560),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_578),
.A2(n_555),
.B(n_549),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_607),
.A2(n_600),
.B1(n_609),
.B2(n_605),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_575),
.B(n_562),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_583),
.Y(n_612)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_612),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_598),
.B(n_580),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_616),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_595),
.B(n_579),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_603),
.A2(n_581),
.B(n_590),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_617),
.A2(n_607),
.B(n_605),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_603),
.A2(n_576),
.B1(n_589),
.B2(n_594),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_618),
.B(n_621),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_606),
.B(n_343),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_602),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_622),
.B(n_597),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_624),
.A2(n_596),
.B(n_608),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_613),
.B(n_601),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_625),
.B(n_632),
.Y(n_635)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_627),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_628),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_629),
.B(n_623),
.C(n_622),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_620),
.A2(n_618),
.B(n_614),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_630),
.A2(n_612),
.B(n_623),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_616),
.B(n_604),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g641 ( 
.A1(n_634),
.A2(n_639),
.B(n_631),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_636),
.A2(n_629),
.B(n_633),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_619),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_640),
.B(n_641),
.C(n_642),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_637),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_642),
.B(n_635),
.C(n_638),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_633),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_645),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_646),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_643),
.Y(n_648)
);


endmodule