module fake_jpeg_13383_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_24),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_25),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_16),
.B1(n_13),
.B2(n_10),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_16),
.B1(n_13),
.B2(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_1),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_7),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_32),
.B1(n_34),
.B2(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_34),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_14),
.B1(n_15),
.B2(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_14),
.B1(n_26),
.B2(n_25),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_2),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_2),
.C(n_3),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_45),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_43),
.B(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_21),
.B1(n_6),
.B2(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_21),
.B1(n_6),
.B2(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_5),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B(n_28),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_29),
.B1(n_32),
.B2(n_22),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_52),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_51),
.C(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_39),
.B1(n_45),
.B2(n_51),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_54),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_57),
.B(n_56),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_57),
.Y(n_62)
);


endmodule