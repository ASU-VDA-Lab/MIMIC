module fake_jpeg_30877_n_455 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_455);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_74),
.Y(n_93)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_32),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_26),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_96),
.B(n_32),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_34),
.C(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_110),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_63),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_34),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_40),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_38),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_63),
.A2(n_34),
.B1(n_40),
.B2(n_30),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_40),
.B1(n_30),
.B2(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_142),
.B1(n_135),
.B2(n_31),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_28),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_28),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_159),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_93),
.B(n_26),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_53),
.B1(n_48),
.B2(n_51),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_71),
.B1(n_114),
.B2(n_118),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_95),
.A2(n_64),
.B1(n_76),
.B2(n_82),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_169),
.B1(n_37),
.B2(n_30),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_93),
.B(n_25),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_28),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_174),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx4f_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_140),
.B(n_126),
.C(n_134),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_168),
.B(n_24),
.CI(n_116),
.CON(n_207),
.SN(n_207)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_38),
.B1(n_32),
.B2(n_46),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx6_ASAP7_75t_SL g172 ( 
.A(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_23),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_23),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_136),
.A3(n_45),
.B1(n_31),
.B2(n_35),
.Y(n_184)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_176),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_37),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_101),
.B1(n_103),
.B2(n_131),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_20),
.B1(n_135),
.B2(n_31),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_180),
.A2(n_183),
.B1(n_185),
.B2(n_160),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_181),
.B(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_166),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_114),
.B1(n_102),
.B2(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_62),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_139),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_176),
.B(n_24),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_214),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_168),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_195),
.B1(n_206),
.B2(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_145),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_221),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_146),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_175),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_158),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_171),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_143),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_227),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.Y(n_247)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_143),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_188),
.B(n_150),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_230),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_195),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_148),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_192),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_172),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_101),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_233),
.A2(n_123),
.B1(n_120),
.B2(n_106),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_185),
.B1(n_183),
.B2(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_236),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_211),
.B1(n_223),
.B2(n_220),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_184),
.B1(n_197),
.B2(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_251),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_206),
.B(n_208),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_201),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_189),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_230),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_242),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_195),
.B(n_186),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_253),
.B(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_163),
.B1(n_199),
.B2(n_167),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_258),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_209),
.A2(n_194),
.B1(n_189),
.B2(n_205),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_192),
.C(n_187),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_229),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_256),
.A2(n_232),
.B1(n_194),
.B2(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_241),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_216),
.B(n_14),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_260),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_274),
.B1(n_279),
.B2(n_243),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_286),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_233),
.B1(n_212),
.B2(n_213),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_238),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_283),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_214),
.B1(n_219),
.B2(n_225),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_147),
.B(n_109),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_237),
.A2(n_224),
.B1(n_221),
.B2(n_205),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_244),
.B(n_249),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_203),
.B1(n_199),
.B2(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_201),
.Y(n_281)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_252),
.B(n_240),
.Y(n_282)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_240),
.B1(n_236),
.B2(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_215),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_285),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_215),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_250),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_250),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_248),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_303),
.B(n_278),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_249),
.C(n_246),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_290),
.B(n_304),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_240),
.C(n_254),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_295),
.C(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_240),
.C(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_238),
.B(n_240),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_268),
.A2(n_239),
.B1(n_246),
.B2(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_307),
.A2(n_280),
.B1(n_265),
.B2(n_284),
.Y(n_329)
);

NAND2xp33_ASAP7_75t_R g308 ( 
.A(n_269),
.B(n_239),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_308),
.A2(n_317),
.B(n_277),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_182),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_164),
.C(n_149),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_313),
.C(n_261),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_286),
.B(n_149),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_311),
.B(n_316),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_182),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_266),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_282),
.Y(n_313)
);

HAxp5_ASAP7_75t_SL g317 ( 
.A(n_272),
.B(n_119),
.CON(n_317),
.SN(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_287),
.Y(n_318)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_327),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_321),
.B(n_288),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_283),
.B1(n_274),
.B2(n_262),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_323),
.A2(n_315),
.B1(n_310),
.B2(n_300),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_271),
.B1(n_267),
.B2(n_260),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_324),
.A2(n_329),
.B1(n_332),
.B2(n_336),
.Y(n_343)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_294),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_288),
.A2(n_271),
.B(n_282),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_328),
.A2(n_312),
.B(n_290),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_320),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_273),
.B1(n_279),
.B2(n_263),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_335),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_299),
.A2(n_285),
.B1(n_281),
.B2(n_162),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_152),
.C(n_138),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_341),
.C(n_288),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_15),
.Y(n_340)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_156),
.C(n_130),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_349),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_334),
.A2(n_289),
.B1(n_305),
.B2(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_348),
.B(n_358),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_338),
.A2(n_303),
.B1(n_295),
.B2(n_306),
.Y(n_350)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_364),
.C(n_341),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_338),
.A2(n_315),
.B1(n_313),
.B2(n_296),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_353),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_327),
.B(n_316),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_334),
.B(n_309),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_360),
.Y(n_371)
);

AOI21x1_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_328),
.B(n_322),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_326),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_157),
.B1(n_178),
.B2(n_141),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_322),
.A2(n_325),
.B1(n_321),
.B2(n_331),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_156),
.C(n_115),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_336),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_375),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_326),
.C(n_329),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_375),
.C(n_372),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_347),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_373),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_339),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_345),
.B(n_319),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_377),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_350),
.B(n_348),
.Y(n_375)
);

BUFx12f_ASAP7_75t_SL g376 ( 
.A(n_355),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_332),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_380),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_360),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_362),
.B(n_361),
.Y(n_383)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_342),
.B(n_330),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_385),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_154),
.B(n_35),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_386),
.B1(n_382),
.B2(n_356),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_392),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_372),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_366),
.B1(n_343),
.B2(n_365),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_376),
.A2(n_351),
.B(n_364),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_394),
.A2(n_395),
.B(n_397),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_368),
.A2(n_343),
.B(n_359),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_141),
.B1(n_129),
.B2(n_67),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_154),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_SL g400 ( 
.A(n_371),
.B(n_14),
.C(n_16),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_13),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_401),
.B(n_378),
.C(n_367),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_407),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_410),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_369),
.C(n_379),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_411),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_390),
.A2(n_121),
.B1(n_72),
.B2(n_70),
.Y(n_409)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_409),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_12),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_11),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_403),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_412),
.A2(n_16),
.B(n_14),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_393),
.B1(n_402),
.B2(n_400),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_414),
.B(n_35),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_11),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_415),
.B(n_416),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_408),
.A2(n_389),
.B(n_388),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_421),
.B(n_423),
.Y(n_438)
);

NOR2x1_ASAP7_75t_L g420 ( 
.A(n_413),
.B(n_392),
.Y(n_420)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_397),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_399),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_0),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_427),
.B(n_428),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_404),
.A2(n_13),
.B(n_1),
.Y(n_428)
);

HAxp5_ASAP7_75t_SL g429 ( 
.A(n_420),
.B(n_409),
.CON(n_429),
.SN(n_429)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_423),
.C(n_4),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_69),
.C(n_59),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_432),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_425),
.A2(n_0),
.B(n_1),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_431),
.A2(n_437),
.B(n_424),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_419),
.A2(n_45),
.B1(n_2),
.B2(n_3),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_436),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_436)
);

NAND5xp2_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_2),
.C(n_4),
.D(n_5),
.E(n_6),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_426),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_441),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_442),
.A2(n_444),
.B1(n_433),
.B2(n_432),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_434),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_39),
.C(n_5),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_445),
.A2(n_437),
.B(n_5),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_447),
.C(n_2),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_429),
.C(n_39),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_443),
.B(n_6),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_450),
.A2(n_451),
.B(n_449),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_7),
.B(n_39),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_7),
.B(n_318),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_7),
.Y(n_455)
);


endmodule