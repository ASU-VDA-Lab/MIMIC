module fake_jpeg_21149_n_185 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_29),
.B(n_26),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_71),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_7),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_74),
.B(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_17),
.B1(n_20),
.B2(n_3),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_14),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_14),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_42),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_9),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_30),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_85),
.C(n_87),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_35),
.C(n_42),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_86),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_45),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_89),
.Y(n_110)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_42),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_92),
.B(n_107),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_30),
.B(n_22),
.Y(n_92)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_42),
.B(n_21),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_85),
.B1(n_65),
.B2(n_78),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_102),
.B1(n_105),
.B2(n_113),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_96),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

OR2x4_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_5),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_13),
.B(n_9),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_11),
.B(n_13),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_105),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_79),
.B1(n_64),
.B2(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_87),
.B1(n_80),
.B2(n_83),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_100),
.B1(n_117),
.B2(n_92),
.Y(n_141)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_126),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_112),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_130),
.B(n_93),
.C(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_65),
.B1(n_78),
.B2(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_104),
.C(n_101),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_122),
.C(n_129),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_93),
.B1(n_104),
.B2(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_117),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_144),
.B(n_141),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_98),
.B(n_108),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_120),
.B(n_116),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_137),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_147),
.B(n_143),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_127),
.C(n_120),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.C(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_125),
.C(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_133),
.B1(n_136),
.B2(n_132),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_155),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_126),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_163),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_162),
.C(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_148),
.B(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_132),
.B1(n_102),
.B2(n_93),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_178),
.B(n_170),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_156),
.A3(n_131),
.B1(n_121),
.B2(n_123),
.C1(n_169),
.C2(n_171),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_182),
.B(n_156),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_169),
.Y(n_185)
);


endmodule