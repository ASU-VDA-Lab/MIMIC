module fake_jpeg_10495_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_48),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_55),
.B1(n_65),
.B2(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_63),
.B1(n_26),
.B2(n_20),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_15),
.B1(n_18),
.B2(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_23),
.Y(n_84)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_38),
.A3(n_41),
.B1(n_23),
.B2(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_75),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_21),
.B(n_36),
.C(n_37),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_60),
.B1(n_53),
.B2(n_46),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_102),
.Y(n_118)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_47),
.B1(n_46),
.B2(n_50),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_85),
.B1(n_56),
.B2(n_76),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_47),
.B1(n_60),
.B2(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_41),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_126),
.Y(n_142)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_114),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_77),
.B1(n_70),
.B2(n_87),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_132),
.B1(n_135),
.B2(n_99),
.Y(n_138)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_130),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_0),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_101),
.B(n_17),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_125),
.Y(n_155)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_131),
.Y(n_149)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_100),
.B1(n_90),
.B2(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_66),
.B1(n_87),
.B2(n_36),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_78),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_140),
.B1(n_113),
.B2(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_97),
.B1(n_108),
.B2(n_105),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_133),
.C(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_158),
.C(n_121),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_124),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_161),
.B(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_8),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_85),
.C(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_14),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_176),
.B1(n_178),
.B2(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_177),
.C(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_172),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_147),
.B(n_141),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_17),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_157),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_181),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_127),
.B1(n_126),
.B2(n_122),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_76),
.C(n_111),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_95),
.B1(n_129),
.B2(n_111),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_32),
.C(n_34),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_185),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_34),
.C(n_35),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_186),
.C(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_34),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_159),
.B1(n_160),
.B2(n_152),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_187),
.A2(n_62),
.B1(n_37),
.B2(n_57),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_154),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_195),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_190),
.B(n_197),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_196),
.C(n_199),
.Y(n_210)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_162),
.C(n_156),
.Y(n_193)
);

OAI322xp33_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_165),
.A3(n_179),
.B1(n_168),
.B2(n_178),
.C1(n_4),
.C2(n_5),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_203),
.B(n_56),
.Y(n_221)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_194),
.C(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_62),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_170),
.C(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_217),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_182),
.C(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_R g235 ( 
.A(n_218),
.B(n_8),
.C(n_1),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_179),
.B1(n_155),
.B2(n_144),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_187),
.B1(n_198),
.B2(n_205),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_144),
.C(n_35),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_35),
.C(n_83),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_62),
.B1(n_37),
.B2(n_57),
.Y(n_234)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_9),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_196),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_210),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_200),
.Y(n_230)
);

AO32x1_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_231),
.A3(n_235),
.B1(n_223),
.B2(n_2),
.Y(n_248)
);

AND2x4_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_237),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_212),
.B1(n_214),
.B2(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_9),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_251),
.B1(n_230),
.B2(n_233),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_245),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_220),
.B1(n_211),
.B2(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_248),
.B1(n_236),
.B2(n_239),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_235),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_227),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_11),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_247),
.A2(n_0),
.B(n_4),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_249),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_250),
.B1(n_247),
.B2(n_10),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_13),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_5),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_57),
.C(n_61),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_61),
.C(n_6),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_61),
.C(n_6),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_267),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_5),
.B(n_6),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_14),
.B(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_261),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_272),
.B(n_273),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_259),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_262),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_264),
.B(n_267),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_275),
.B(n_274),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_278),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_14),
.Y(n_280)
);


endmodule