module fake_jpeg_18223_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_58),
.B1(n_46),
.B2(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_49),
.B1(n_59),
.B2(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_3),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_54),
.B1(n_47),
.B2(n_48),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_44),
.B(n_49),
.C(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_88),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_41),
.B1(n_55),
.B2(n_45),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_42),
.B1(n_39),
.B2(n_5),
.Y(n_96)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_92),
.Y(n_102)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_2),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_4),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_112),
.B1(n_93),
.B2(n_94),
.Y(n_116)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_111),
.B1(n_101),
.B2(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_8),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_117),
.C(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_113),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_110),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_115),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_118),
.B1(n_115),
.B2(n_17),
.C(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_15),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_16),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_20),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_23),
.C(n_24),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_25),
.Y(n_128)
);


endmodule