module real_aes_4169_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_713;
wire n_147;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_649;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_639;
wire n_546;
wire n_151;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_0), .A2(n_15), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_0), .Y(n_131) );
INVx1_ASAP7_75t_L g604 ( .A(n_1), .Y(n_604) );
INVx1_ASAP7_75t_L g313 ( .A(n_2), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_3), .A2(n_19), .B1(n_220), .B2(n_263), .Y(n_283) );
INVx2_ASAP7_75t_L g170 ( .A(n_4), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_5), .B(n_617), .Y(n_715) );
INVx1_ASAP7_75t_SL g232 ( .A(n_6), .Y(n_232) );
BUFx2_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
INVxp67_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g557 ( .A(n_7), .Y(n_557) );
INVx1_ASAP7_75t_L g562 ( .A(n_7), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_8), .B(n_209), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_9), .A2(n_40), .B1(n_616), .B2(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_10), .A2(n_46), .B1(n_261), .B2(n_596), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_11), .A2(n_68), .B1(n_578), .B2(n_579), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_12), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_13), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g599 ( .A(n_14), .Y(n_599) );
INVx1_ASAP7_75t_L g130 ( .A(n_15), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_16), .A2(n_56), .B1(n_208), .B2(n_209), .Y(n_207) );
INVx1_ASAP7_75t_L g602 ( .A(n_17), .Y(n_602) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_18), .A2(n_72), .B(n_150), .Y(n_149) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_18), .A2(n_72), .B(n_150), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_20), .A2(n_70), .B1(n_578), .B2(n_579), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_21), .B(n_166), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_22), .A2(n_82), .B1(n_153), .B2(n_156), .Y(n_152) );
INVx2_ASAP7_75t_L g267 ( .A(n_23), .Y(n_267) );
INVx1_ASAP7_75t_L g595 ( .A(n_24), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_25), .A2(n_29), .B1(n_192), .B2(n_231), .Y(n_284) );
BUFx3_ASAP7_75t_L g115 ( .A(n_26), .Y(n_115) );
O2A1O1Ixp5_ASAP7_75t_L g260 ( .A1(n_27), .A2(n_190), .B(n_261), .C(n_262), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_28), .A2(n_65), .B1(n_163), .B2(n_165), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_30), .Y(n_194) );
AO22x1_ASAP7_75t_L g712 ( .A1(n_31), .A2(n_80), .B1(n_237), .B2(n_713), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_32), .Y(n_620) );
AND2x2_ASAP7_75t_L g630 ( .A(n_33), .B(n_596), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_34), .B(n_237), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_35), .A2(n_83), .B1(n_217), .B2(n_219), .Y(n_216) );
INVx1_ASAP7_75t_L g105 ( .A(n_36), .Y(n_105) );
INVx1_ASAP7_75t_L g256 ( .A(n_37), .Y(n_256) );
AOI22x1_ASAP7_75t_L g652 ( .A1(n_38), .A2(n_97), .B1(n_578), .B2(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_39), .B(n_655), .Y(n_668) );
AND2x2_ASAP7_75t_L g111 ( .A(n_41), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_42), .B(n_252), .Y(n_308) );
INVx2_ASAP7_75t_L g264 ( .A(n_43), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_44), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_45), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g272 ( .A(n_47), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_48), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g236 ( .A(n_49), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_50), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_51), .B(n_231), .Y(n_684) );
INVx1_ASAP7_75t_L g186 ( .A(n_52), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_53), .B(n_258), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_54), .Y(n_956) );
INVx1_ASAP7_75t_L g150 ( .A(n_55), .Y(n_150) );
AND2x4_ASAP7_75t_L g144 ( .A(n_57), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g181 ( .A(n_57), .B(n_145), .Y(n_181) );
INVx1_ASAP7_75t_L g241 ( .A(n_58), .Y(n_241) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_59), .Y(n_161) );
INVx2_ASAP7_75t_L g581 ( .A(n_60), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_61), .A2(n_75), .B1(n_616), .B2(n_653), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_62), .Y(n_548) );
CKINVDCx14_ASAP7_75t_R g718 ( .A(n_63), .Y(n_718) );
AND2x2_ASAP7_75t_L g636 ( .A(n_64), .B(n_237), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_66), .B(n_234), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_67), .B(n_306), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_69), .B(n_300), .Y(n_678) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_71), .B(n_583), .Y(n_640) );
CKINVDCx14_ASAP7_75t_R g657 ( .A(n_73), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_74), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_76), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_77), .B(n_617), .Y(n_682) );
INVx1_ASAP7_75t_L g108 ( .A(n_78), .Y(n_108) );
OR2x6_ASAP7_75t_L g124 ( .A(n_78), .B(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_79), .B(n_157), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_81), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g112 ( .A(n_84), .Y(n_112) );
INVx1_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_85), .Y(n_158) );
BUFx5_ASAP7_75t_L g193 ( .A(n_85), .Y(n_193) );
INVx2_ASAP7_75t_L g606 ( .A(n_86), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_87), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g963 ( .A(n_88), .B(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g275 ( .A(n_89), .Y(n_275) );
INVx1_ASAP7_75t_L g279 ( .A(n_90), .Y(n_279) );
NAND2xp33_ASAP7_75t_L g632 ( .A(n_91), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g200 ( .A(n_92), .Y(n_200) );
INVx2_ASAP7_75t_SL g145 ( .A(n_93), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_94), .B(n_183), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_95), .B(n_639), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_96), .B(n_300), .Y(n_299) );
AO32x2_ASAP7_75t_L g281 ( .A1(n_98), .A2(n_265), .A3(n_282), .B1(n_286), .B2(n_287), .Y(n_281) );
AO22x2_ASAP7_75t_L g318 ( .A1(n_98), .A2(n_282), .B1(n_319), .B2(n_321), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_99), .B(n_627), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_113), .B(n_963), .Y(n_100) );
BUFx2_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
BUFx16f_ASAP7_75t_R g965 ( .A(n_102), .Y(n_965) );
AND2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_105), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .C(n_111), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_116), .B(n_551), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
CKINVDCx6p67_ASAP7_75t_R g962 ( .A(n_115), .Y(n_962) );
OAI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_127), .B(n_547), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx4f_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_119), .Y(n_550) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OR2x6_ASAP7_75t_L g561 ( .A(n_123), .B(n_562), .Y(n_561) );
INVx8_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g556 ( .A(n_124), .B(n_557), .Y(n_556) );
OR2x6_ASAP7_75t_L g958 ( .A(n_124), .B(n_557), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_132), .B2(n_546), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
XNOR2x1_ASAP7_75t_L g558 ( .A(n_131), .B(n_134), .Y(n_558) );
INVx1_ASAP7_75t_L g546 ( .A(n_132), .Y(n_546) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_470), .Y(n_134) );
NOR2xp67_ASAP7_75t_L g135 ( .A(n_136), .B(n_392), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_334), .C(n_371), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_242), .B(n_288), .Y(n_137) );
OAI31xp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_172), .A3(n_203), .B(n_223), .Y(n_138) );
INVx1_ASAP7_75t_L g529 ( .A(n_139), .Y(n_529) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g366 ( .A(n_140), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g398 ( .A(n_140), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_140), .B(n_325), .Y(n_412) );
AND2x2_ASAP7_75t_L g516 ( .A(n_140), .B(n_502), .Y(n_516) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g390 ( .A(n_141), .B(n_346), .Y(n_390) );
AND2x2_ASAP7_75t_L g429 ( .A(n_141), .B(n_326), .Y(n_429) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_141), .Y(n_463) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g343 ( .A(n_142), .Y(n_343) );
INVx1_ASAP7_75t_L g362 ( .A(n_142), .Y(n_362) );
AOI21x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_151), .B(n_169), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx3_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_144), .Y(n_286) );
AND2x2_ASAP7_75t_L g319 ( .A(n_144), .B(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g576 ( .A(n_144), .Y(n_576) );
INVx1_ASAP7_75t_L g591 ( .A(n_144), .Y(n_591) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_146), .A2(n_575), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_147), .B(n_212), .Y(n_228) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g583 ( .A(n_148), .Y(n_583) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
BUFx3_ASAP7_75t_L g198 ( .A(n_149), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_159), .B1(n_162), .B2(n_167), .Y(n_151) );
INVx2_ASAP7_75t_L g713 ( .A(n_153), .Y(n_713) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
INVx1_ASAP7_75t_L g579 ( .A(n_156), .Y(n_579) );
INVx1_ASAP7_75t_L g667 ( .A(n_156), .Y(n_667) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
INVx2_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
INVx1_ASAP7_75t_L g304 ( .A(n_157), .Y(n_304) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx6_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
INVx2_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx2_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
AOI21x1_ASAP7_75t_L g711 ( .A1(n_159), .A2(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_160), .B(n_211), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_160), .A2(n_230), .B(n_232), .C(n_233), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_160), .A2(n_178), .B(n_275), .C(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g285 ( .A(n_160), .Y(n_285) );
INVxp67_ASAP7_75t_L g625 ( .A(n_160), .Y(n_625) );
INVx2_ASAP7_75t_SL g642 ( .A(n_160), .Y(n_642) );
INVx1_ASAP7_75t_L g686 ( .A(n_160), .Y(n_686) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_161), .Y(n_190) );
INVx1_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
INVx4_ASAP7_75t_L g253 ( .A(n_161), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_161), .B(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_161), .B(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_L g634 ( .A(n_161), .Y(n_634) );
INVx3_ASAP7_75t_L g261 ( .A(n_163), .Y(n_261) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
INVx1_ASAP7_75t_L g271 ( .A(n_165), .Y(n_271) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
INVx2_ASAP7_75t_L g250 ( .A(n_166), .Y(n_250) );
INVx2_ASAP7_75t_SL g263 ( .A(n_166), .Y(n_263) );
INVx1_ASAP7_75t_L g633 ( .A(n_166), .Y(n_633) );
INVx1_ASAP7_75t_L g639 ( .A(n_166), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_167), .B(n_180), .Y(n_179) );
NOR3xp33_ASAP7_75t_L g185 ( .A(n_167), .B(n_180), .C(n_186), .Y(n_185) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_167), .B(n_574), .C(n_575), .Y(n_585) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_168), .A2(n_236), .B(n_237), .C(n_238), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_168), .A2(n_271), .B(n_272), .C(n_273), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
BUFx3_ASAP7_75t_L g265 ( .A(n_171), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_171), .B(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g300 ( .A(n_171), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_171), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g353 ( .A(n_172), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_172), .B(n_354), .Y(n_446) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g226 ( .A(n_173), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g331 ( .A(n_173), .Y(n_331) );
AND2x2_ASAP7_75t_L g464 ( .A(n_173), .B(n_367), .Y(n_464) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_197), .B(n_199), .Y(n_173) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_174), .A2(n_199), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_187), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B1(n_182), .B2(n_185), .Y(n_175) );
NOR2xp67_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_180), .B(n_189), .Y(n_188) );
AOI221x1_ASAP7_75t_L g247 ( .A1(n_180), .A2(n_248), .B1(n_251), .B2(n_255), .C(n_257), .Y(n_247) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g218 ( .A(n_184), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_191), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_189), .B(n_619), .Y(n_618) );
OAI22x1_ASAP7_75t_L g649 ( .A1(n_189), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_190), .A2(n_283), .B1(n_284), .B2(n_285), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_190), .A2(n_303), .B(n_305), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_190), .A2(n_616), .B1(n_618), .B2(n_621), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_190), .B(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_190), .A2(n_681), .B(n_682), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g208 ( .A(n_193), .Y(n_208) );
INVx2_ASAP7_75t_L g237 ( .A(n_193), .Y(n_237) );
INVx2_ASAP7_75t_L g306 ( .A(n_193), .Y(n_306) );
INVx1_ASAP7_75t_L g310 ( .A(n_193), .Y(n_310) );
INVx2_ASAP7_75t_L g617 ( .A(n_193), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_195), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g596 ( .A(n_195), .Y(n_596) );
NOR2xp67_ASAP7_75t_SL g656 ( .A(n_197), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g717 ( .A(n_197), .B(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OA21x2_ASAP7_75t_L g613 ( .A1(n_198), .A2(n_614), .B(n_626), .Y(n_613) );
OA21x2_ASAP7_75t_L g704 ( .A1(n_198), .A2(n_614), .B(n_626), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g287 ( .A(n_201), .Y(n_287) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp67_ASAP7_75t_L g211 ( .A(n_202), .B(n_212), .Y(n_211) );
BUFx3_ASAP7_75t_L g214 ( .A(n_202), .Y(n_214) );
INVx1_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_202), .B(n_212), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_202), .B(n_212), .Y(n_314) );
INVx1_ASAP7_75t_L g320 ( .A(n_202), .Y(n_320) );
INVx2_ASAP7_75t_L g574 ( .A(n_202), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_202), .B(n_212), .Y(n_662) );
BUFx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g494 ( .A(n_204), .B(n_405), .Y(n_494) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g225 ( .A(n_205), .Y(n_225) );
INVx2_ASAP7_75t_L g330 ( .A(n_205), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_205), .B(n_298), .Y(n_349) );
AND2x2_ASAP7_75t_L g354 ( .A(n_205), .B(n_355), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_206), .B(n_215), .Y(n_205) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_206), .B(n_215), .Y(n_293) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_210), .B(n_213), .Y(n_206) );
INVx2_ASAP7_75t_L g578 ( .A(n_208), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_211), .B(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_221), .Y(n_215) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
INVx1_ASAP7_75t_L g651 ( .A(n_222), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_222), .B(n_662), .Y(n_665) );
INVx2_ASAP7_75t_L g508 ( .A(n_223), .Y(n_508) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
AND2x4_ASAP7_75t_L g433 ( .A(n_224), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g448 ( .A(n_225), .B(n_332), .Y(n_448) );
INVx2_ASAP7_75t_L g410 ( .A(n_226), .Y(n_410) );
INVx1_ASAP7_75t_L g315 ( .A(n_227), .Y(n_315) );
INVx2_ASAP7_75t_L g333 ( .A(n_227), .Y(n_333) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_227), .Y(n_348) );
INVx2_ASAP7_75t_L g367 ( .A(n_227), .Y(n_367) );
AND2x2_ASAP7_75t_L g381 ( .A(n_227), .B(n_294), .Y(n_381) );
INVx1_ASAP7_75t_L g406 ( .A(n_227), .Y(n_406) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .A3(n_235), .B(n_239), .Y(n_227) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_237), .A2(n_258), .B1(n_601), .B2(n_603), .Y(n_600) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_240), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g655 ( .A(n_240), .Y(n_655) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_244), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_280), .Y(n_244) );
AND2x2_ASAP7_75t_L g337 ( .A(n_245), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g365 ( .A(n_245), .Y(n_365) );
INVx2_ASAP7_75t_L g423 ( .A(n_245), .Y(n_423) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_268), .Y(n_245) );
INVx2_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_246), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g397 ( .A(n_246), .B(n_343), .Y(n_397) );
INVx1_ASAP7_75t_L g438 ( .A(n_246), .Y(n_438) );
AND2x2_ASAP7_75t_L g502 ( .A(n_246), .B(n_346), .Y(n_502) );
AO31x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_259), .A3(n_265), .B(n_266), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g255 ( .A(n_252), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_253), .B(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_SL g573 ( .A(n_253), .B(n_574), .C(n_575), .Y(n_573) );
NOR2xp33_ASAP7_75t_SL g601 ( .A(n_253), .B(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_253), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_258), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g321 ( .A(n_265), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_268), .Y(n_322) );
INVx2_ASAP7_75t_L g346 ( .A(n_268), .Y(n_346) );
AND2x4_ASAP7_75t_L g358 ( .A(n_268), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g400 ( .A(n_268), .Y(n_400) );
AND2x4_ASAP7_75t_L g437 ( .A(n_268), .B(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .A3(n_277), .B(n_278), .Y(n_269) );
INVx1_ASAP7_75t_L g413 ( .A(n_280), .Y(n_413) );
INVx2_ASAP7_75t_L g415 ( .A(n_280), .Y(n_415) );
AND2x4_ASAP7_75t_L g444 ( .A(n_280), .B(n_429), .Y(n_444) );
AND2x2_ASAP7_75t_L g510 ( .A(n_280), .B(n_511), .Y(n_510) );
BUFx8_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g359 ( .A(n_281), .Y(n_359) );
AND2x2_ASAP7_75t_L g374 ( .A(n_281), .B(n_375), .Y(n_374) );
OAI21x1_ASAP7_75t_L g614 ( .A1(n_286), .A2(n_615), .B(n_622), .Y(n_614) );
AO31x2_ASAP7_75t_L g648 ( .A1(n_286), .A2(n_649), .A3(n_654), .B(n_656), .Y(n_648) );
AO31x2_ASAP7_75t_L g692 ( .A1(n_286), .A2(n_649), .A3(n_654), .B(n_656), .Y(n_692) );
INVxp67_ASAP7_75t_L g295 ( .A(n_287), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_316), .B1(n_323), .B2(n_327), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_289), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI211xp5_ASAP7_75t_L g489 ( .A1(n_290), .A2(n_372), .B(n_490), .C(n_496), .Y(n_489) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_296), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NOR2xp67_ASAP7_75t_SL g483 ( .A(n_292), .B(n_385), .Y(n_483) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g418 ( .A(n_293), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g425 ( .A(n_293), .B(n_419), .Y(n_425) );
INVx1_ASAP7_75t_L g531 ( .A(n_293), .Y(n_531) );
OR2x2_ASAP7_75t_L g370 ( .A(n_294), .B(n_355), .Y(n_370) );
AND2x2_ASAP7_75t_L g377 ( .A(n_294), .B(n_330), .Y(n_377) );
AND2x2_ASAP7_75t_L g495 ( .A(n_294), .B(n_297), .Y(n_495) );
AND2x2_ASAP7_75t_L g454 ( .A(n_296), .B(n_377), .Y(n_454) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_315), .Y(n_296) );
OR2x2_ASAP7_75t_L g385 ( .A(n_297), .B(n_331), .Y(n_385) );
INVx1_ASAP7_75t_L g479 ( .A(n_297), .Y(n_479) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g332 ( .A(n_298), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
INVx1_ASAP7_75t_L g419 ( .A(n_298), .Y(n_419) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_300), .B(n_576), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_307), .B(n_314), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B(n_311), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_L g391 ( .A(n_315), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_315), .B(n_505), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_316), .A2(n_411), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
INVx1_ASAP7_75t_L g338 ( .A(n_318), .Y(n_338) );
AND2x4_ASAP7_75t_L g345 ( .A(n_318), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
AND2x2_ASAP7_75t_L g519 ( .A(n_318), .B(n_343), .Y(n_519) );
INVx2_ASAP7_75t_SL g395 ( .A(n_322), .Y(n_395) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_324), .B(n_395), .Y(n_467) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g386 ( .A(n_325), .B(n_359), .Y(n_386) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g373 ( .A(n_326), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_326), .B(n_359), .Y(n_388) );
BUFx3_ASAP7_75t_L g486 ( .A(n_326), .Y(n_486) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g383 ( .A1(n_329), .A2(n_384), .B1(n_386), .B2(n_387), .Y(n_383) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_330), .Y(n_458) );
BUFx2_ASAP7_75t_L g505 ( .A(n_330), .Y(n_505) );
AND2x4_ASAP7_75t_L g442 ( .A(n_331), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g376 ( .A(n_332), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g443 ( .A(n_333), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_347), .B(n_350), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_337), .B(n_529), .Y(n_534) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
OAI21xp33_ASAP7_75t_SL g378 ( .A1(n_341), .A2(n_344), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g474 ( .A(n_341), .Y(n_474) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g511 ( .A(n_342), .Y(n_511) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_343), .Y(n_542) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_345), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g380 ( .A(n_349), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g461 ( .A(n_349), .Y(n_461) );
AND2x2_ASAP7_75t_L g509 ( .A(n_349), .B(n_464), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_356), .B1(n_363), .B2(n_368), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_353), .B(n_536), .Y(n_535) );
NAND2xp67_ASAP7_75t_L g409 ( .A(n_354), .B(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g431 ( .A(n_354), .Y(n_431) );
AND2x2_ASAP7_75t_L g539 ( .A(n_354), .B(n_442), .Y(n_539) );
AND2x2_ASAP7_75t_L g545 ( .A(n_354), .B(n_381), .Y(n_545) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_358), .B(n_361), .Y(n_379) );
INVx2_ASAP7_75t_L g491 ( .A(n_358), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_359), .B(n_375), .Y(n_453) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_SL g426 ( .A(n_361), .Y(n_426) );
AND2x2_ASAP7_75t_L g527 ( .A(n_361), .B(n_437), .Y(n_527) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g375 ( .A(n_362), .Y(n_375) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NOR2xp67_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_367), .Y(n_469) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g514 ( .A(n_369), .B(n_494), .Y(n_514) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g434 ( .A(n_370), .Y(n_434) );
OR2x6_ASAP7_75t_L g468 ( .A(n_370), .B(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_370), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B1(n_378), .B2(n_380), .C(n_382), .Y(n_371) );
AND2x4_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g498 ( .A(n_374), .Y(n_498) );
AND2x4_ASAP7_75t_L g403 ( .A(n_377), .B(n_404), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_389), .C(n_391), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g541 ( .A(n_388), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g485 ( .A(n_390), .B(n_486), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_420), .C(n_436), .D(n_449), .Y(n_392) );
O2A1O1Ixp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_398), .B(n_402), .C(n_408), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g460 ( .A(n_395), .Y(n_460) );
OAI32xp33_ASAP7_75t_L g528 ( .A1(n_395), .A2(n_416), .A3(n_497), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g414 ( .A(n_397), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g523 ( .A(n_397), .Y(n_523) );
INVx1_ASAP7_75t_L g459 ( .A(n_399), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_399), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g544 ( .A(n_399), .B(n_486), .Y(n_544) );
AND2x4_ASAP7_75t_SL g399 ( .A(n_400), .B(n_401), .Y(n_399) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_405), .Y(n_417) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI32xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .A3(n_413), .B1(n_414), .B2(n_416), .Y(n_408) );
AND2x2_ASAP7_75t_L g424 ( .A(n_410), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g475 ( .A(n_414), .Y(n_475) );
AND2x2_ASAP7_75t_L g501 ( .A(n_415), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g536 ( .A(n_418), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_426), .B(n_427), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_423), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_423), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g441 ( .A(n_425), .B(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_432), .B2(n_435), .Y(n_427) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_429), .B(n_452), .Y(n_466) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_435), .A2(n_491), .B(n_492), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_444), .B2(n_445), .Y(n_436) );
INVx2_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_437), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g478 ( .A(n_442), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g504 ( .A(n_442), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI221xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_454), .B1(n_455), .B2(n_462), .C(n_465), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_457), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g487 ( .A(n_458), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx2_ASAP7_75t_L g526 ( .A(n_464), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_464), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_468), .Y(n_465) );
NOR2x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_506), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .C(n_489), .Y(n_471) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .B(n_476), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_483), .A2(n_521), .B1(n_524), .B2(n_527), .C(n_528), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_500), .B(n_503), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g525 ( .A(n_505), .Y(n_525) );
NAND3xp33_ASAP7_75t_SL g506 ( .A(n_507), .B(n_520), .C(n_532), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_510), .C(n_512), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_515), .B1(n_517), .B2(n_518), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2x1p5_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B(n_537), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .B(n_543), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NOR2xp33_ASAP7_75t_R g944 ( .A(n_548), .B(n_549), .Y(n_944) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_945), .B(n_959), .Y(n_551) );
AOI21xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_943), .B(n_944), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_558), .B(n_559), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_555), .Y(n_554) );
BUFx8_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_556), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g947 ( .A1(n_558), .A2(n_948), .B(n_951), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g954 ( .A(n_561), .Y(n_954) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_565), .B(n_952), .Y(n_951) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_566), .B(n_817), .Y(n_565) );
NOR4xp75_ASAP7_75t_L g566 ( .A(n_567), .B(n_730), .C(n_748), .D(n_774), .Y(n_566) );
AO21x1_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_607), .B(n_698), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_570), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g738 ( .A(n_570), .B(n_708), .Y(n_738) );
INVx2_ASAP7_75t_L g800 ( .A(n_570), .Y(n_800) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_587), .Y(n_570) );
INVx1_ASAP7_75t_L g672 ( .A(n_571), .Y(n_672) );
INVx1_ASAP7_75t_L g697 ( .A(n_571), .Y(n_697) );
AND2x2_ASAP7_75t_L g720 ( .A(n_571), .B(n_588), .Y(n_720) );
INVx1_ASAP7_75t_L g751 ( .A(n_571), .Y(n_751) );
INVx2_ASAP7_75t_L g783 ( .A(n_571), .Y(n_783) );
NOR2x1_ASAP7_75t_L g825 ( .A(n_571), .B(n_826), .Y(n_825) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_571), .Y(n_840) );
AND2x2_ASAP7_75t_L g889 ( .A(n_571), .B(n_676), .Y(n_889) );
OR2x6_ASAP7_75t_L g571 ( .A(n_572), .B(n_584), .Y(n_571) );
OAI21x1_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B(n_580), .Y(n_572) );
INVx1_ASAP7_75t_L g590 ( .A(n_574), .Y(n_590) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g627 ( .A(n_582), .Y(n_627) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AND2x2_ASAP7_75t_L g782 ( .A(n_587), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g787 ( .A(n_588), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g807 ( .A(n_588), .Y(n_807) );
INVx1_ASAP7_75t_L g826 ( .A(n_588), .Y(n_826) );
AND2x2_ASAP7_75t_L g888 ( .A(n_588), .B(n_753), .Y(n_888) );
INVxp67_ASAP7_75t_L g918 ( .A(n_588), .Y(n_918) );
AO21x2_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B(n_605), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OR2x2_ASAP7_75t_L g710 ( .A(n_591), .B(n_627), .Y(n_710) );
NAND3xp33_ASAP7_75t_SL g592 ( .A(n_593), .B(n_597), .C(n_600), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_669), .B1(n_688), .B2(n_695), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_610), .B(n_645), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g859 ( .A(n_611), .Y(n_859) );
OR2x2_ASAP7_75t_L g941 ( .A(n_611), .B(n_773), .Y(n_941) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g772 ( .A(n_612), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_628), .Y(n_612) );
AND2x2_ASAP7_75t_L g689 ( .A(n_613), .B(n_690), .Y(n_689) );
NAND2x1_ASAP7_75t_L g734 ( .A(n_613), .B(n_647), .Y(n_734) );
AND2x2_ASAP7_75t_L g869 ( .A(n_613), .B(n_659), .Y(n_869) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g699 ( .A(n_628), .B(n_692), .Y(n_699) );
AND2x4_ASAP7_75t_L g723 ( .A(n_628), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g842 ( .A(n_628), .B(n_692), .Y(n_842) );
AO21x2_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_635), .B(n_643), .Y(n_628) );
AO21x2_ASAP7_75t_L g694 ( .A1(n_629), .A2(n_635), .B(n_643), .Y(n_694) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g653 ( .A(n_633), .Y(n_653) );
OAI21x1_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_637), .B(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_640), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_640), .Y(n_644) );
AOI21x1_ASAP7_75t_L g714 ( .A1(n_642), .A2(n_715), .B(n_716), .Y(n_714) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_658), .Y(n_645) );
INVx2_ASAP7_75t_L g725 ( .A(n_646), .Y(n_725) );
INVx1_ASAP7_75t_L g757 ( .A(n_646), .Y(n_757) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g747 ( .A(n_647), .B(n_694), .Y(n_747) );
INVx1_ASAP7_75t_L g761 ( .A(n_647), .Y(n_761) );
AND2x2_ASAP7_75t_L g901 ( .A(n_647), .B(n_705), .Y(n_901) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g773 ( .A(n_658), .Y(n_773) );
OR2x2_ASAP7_75t_L g885 ( .A(n_658), .B(n_734), .Y(n_885) );
INVx2_ASAP7_75t_L g893 ( .A(n_658), .Y(n_893) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_660), .B(n_664), .Y(n_690) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
OA21x2_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g808 ( .A(n_672), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g833 ( .A(n_674), .B(n_793), .Y(n_833) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g767 ( .A(n_675), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g708 ( .A(n_676), .B(n_709), .Y(n_708) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g729 ( .A(n_677), .Y(n_729) );
AND2x2_ASAP7_75t_L g752 ( .A(n_677), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g764 ( .A(n_677), .B(n_709), .Y(n_764) );
AND2x4_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B(n_687), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B(n_686), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g789 ( .A(n_689), .B(n_733), .Y(n_789) );
INVx1_ASAP7_75t_L g902 ( .A(n_689), .Y(n_902) );
AND2x2_ASAP7_75t_L g934 ( .A(n_689), .B(n_761), .Y(n_934) );
INVx2_ASAP7_75t_L g705 ( .A(n_690), .Y(n_705) );
AND2x2_ASAP7_75t_L g744 ( .A(n_690), .B(n_703), .Y(n_744) );
INVx1_ASAP7_75t_L g794 ( .A(n_690), .Y(n_794) );
INVx1_ASAP7_75t_L g846 ( .A(n_690), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_690), .B(n_813), .Y(n_854) );
BUFx3_ASAP7_75t_L g741 ( .A(n_691), .Y(n_741) );
NOR2xp67_ASAP7_75t_L g861 ( .A(n_691), .B(n_743), .Y(n_861) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g771 ( .A(n_692), .Y(n_771) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g733 ( .A(n_694), .Y(n_733) );
INVx1_ASAP7_75t_L g813 ( .A(n_694), .Y(n_813) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g763 ( .A(n_696), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g766 ( .A(n_696), .B(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_696), .Y(n_795) );
OR2x2_ASAP7_75t_L g922 ( .A(n_696), .B(n_799), .Y(n_922) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g785 ( .A(n_697), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_697), .B(n_851), .Y(n_850) );
OAI32xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .A3(n_706), .B1(n_721), .B2(n_726), .Y(n_698) );
INVx2_ASAP7_75t_L g857 ( .A(n_699), .Y(n_857) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g884 ( .A(n_701), .Y(n_884) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g804 ( .A(n_702), .Y(n_804) );
OR2x2_ASAP7_75t_L g811 ( .A(n_702), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g896 ( .A(n_703), .Y(n_896) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g724 ( .A(n_704), .Y(n_724) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_704), .Y(n_852) );
INVx1_ASAP7_75t_L g746 ( .A(n_705), .Y(n_746) );
INVx2_ASAP7_75t_L g736 ( .A(n_706), .Y(n_736) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_719), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g824 ( .A(n_708), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g911 ( .A(n_708), .B(n_782), .Y(n_911) );
INVx2_ASAP7_75t_SL g753 ( .A(n_709), .Y(n_753) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_717), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_710), .A2(n_711), .B(n_717), .Y(n_788) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g860 ( .A(n_720), .B(n_764), .Y(n_860) );
NAND2x1_ASAP7_75t_SL g882 ( .A(n_720), .B(n_752), .Y(n_882) );
AND2x2_ASAP7_75t_L g891 ( .A(n_720), .B(n_780), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_720), .B(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g935 ( .A(n_722), .B(n_793), .Y(n_935) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
AND2x4_ASAP7_75t_SL g760 ( .A(n_723), .B(n_761), .Y(n_760) );
BUFx3_ASAP7_75t_L g836 ( .A(n_723), .Y(n_836) );
INVxp67_ASAP7_75t_SL g829 ( .A(n_724), .Y(n_829) );
INVx1_ASAP7_75t_L g862 ( .A(n_726), .Y(n_862) );
AOI211xp5_ASAP7_75t_SL g849 ( .A1(n_727), .A2(n_761), .B(n_850), .C(n_852), .Y(n_849) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g806 ( .A(n_728), .B(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g864 ( .A(n_728), .B(n_865), .Y(n_864) );
AND2x2_ASAP7_75t_L g931 ( .A(n_728), .B(n_782), .Y(n_931) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g815 ( .A(n_729), .B(n_751), .Y(n_815) );
OR2x2_ASAP7_75t_L g830 ( .A(n_729), .B(n_787), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g917 ( .A(n_729), .B(n_918), .Y(n_917) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_735), .B1(n_737), .B2(n_739), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_733), .Y(n_828) );
AND3x2_ASAP7_75t_L g908 ( .A(n_733), .B(n_893), .C(n_896), .Y(n_908) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OA21x2_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_742), .B(n_745), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g927 ( .A(n_742), .Y(n_927) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g758 ( .A(n_744), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
BUFx3_ASAP7_75t_L g822 ( .A(n_747), .Y(n_822) );
AND2x2_ASAP7_75t_L g892 ( .A(n_747), .B(n_893), .Y(n_892) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_754), .B(n_762), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
AND2x2_ASAP7_75t_L g872 ( .A(n_752), .B(n_782), .Y(n_872) );
INVx2_ASAP7_75t_L g880 ( .A(n_752), .Y(n_880) );
INVx1_ASAP7_75t_L g768 ( .A(n_753), .Y(n_768) );
INVx1_ASAP7_75t_L g797 ( .A(n_753), .Y(n_797) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_756), .B(n_759), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_756), .A2(n_777), .B1(n_792), .B2(n_798), .Y(n_791) );
OR2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
OR2x2_ASAP7_75t_L g867 ( .A(n_757), .B(n_868), .Y(n_867) );
INVx2_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g777 ( .A(n_760), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_765), .B(n_769), .Y(n_762) );
INVx2_ASAP7_75t_L g799 ( .A(n_764), .Y(n_799) );
AND2x2_ASAP7_75t_L g844 ( .A(n_764), .B(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_766), .A2(n_867), .B1(n_895), .B2(n_897), .Y(n_894) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_768), .Y(n_780) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_770), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_770), .B(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND3x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_790), .C(n_801), .Y(n_774) );
AOI21x1_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B(n_784), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_779), .A2(n_864), .B1(n_941), .B2(n_942), .Y(n_940) );
OR2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_789), .Y(n_784) );
INVx1_ASAP7_75t_L g834 ( .A(n_786), .Y(n_834) );
AND2x2_ASAP7_75t_L g914 ( .A(n_786), .B(n_840), .Y(n_914) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g816 ( .A(n_787), .Y(n_816) );
BUFx2_ASAP7_75t_L g809 ( .A(n_788), .Y(n_809) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .C(n_796), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g848 ( .A(n_797), .B(n_807), .Y(n_848) );
OR2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVxp67_ASAP7_75t_L g838 ( .A(n_800), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_805), .B1(n_810), .B2(n_814), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND3xp33_ASAP7_75t_SL g856 ( .A(n_803), .B(n_857), .C(n_858), .Y(n_856) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_808), .Y(n_805) );
AND2x2_ASAP7_75t_L g916 ( .A(n_808), .B(n_917), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_808), .B(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g851 ( .A(n_809), .Y(n_851) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_812), .B(n_846), .Y(n_942) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_813), .A2(n_838), .B1(n_839), .B2(n_841), .Y(n_837) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
NAND2x2_ASAP7_75t_L g925 ( .A(n_815), .B(n_926), .Y(n_925) );
NOR2x1_ASAP7_75t_L g817 ( .A(n_818), .B(n_903), .Y(n_817) );
NAND4xp25_ASAP7_75t_L g818 ( .A(n_819), .B(n_855), .C(n_870), .D(n_890), .Y(n_818) );
NOR2xp67_ASAP7_75t_L g819 ( .A(n_820), .B(n_831), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B1(n_827), .B2(n_830), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AOI21xp33_ASAP7_75t_L g912 ( .A1(n_823), .A2(n_835), .B(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g865 ( .A(n_825), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
OAI211xp5_ASAP7_75t_SL g847 ( .A1(n_829), .A2(n_848), .B(n_849), .C(n_853), .Y(n_847) );
INVx1_ASAP7_75t_L g874 ( .A(n_829), .Y(n_874) );
AOI21xp33_ASAP7_75t_L g899 ( .A1(n_830), .A2(n_900), .B(n_902), .Y(n_899) );
OAI321xp33_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_834), .A3(n_835), .B1(n_837), .B2(n_843), .C(n_847), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
OR2x2_ASAP7_75t_L g897 ( .A(n_834), .B(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_836), .B(n_877), .Y(n_876) );
NOR2x1_ASAP7_75t_R g919 ( .A(n_836), .B(n_900), .Y(n_919) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g920 ( .A(n_841), .B(n_869), .Y(n_920) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
OR2x2_ASAP7_75t_L g895 ( .A(n_842), .B(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g907 ( .A(n_842), .Y(n_907) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g877 ( .A(n_846), .Y(n_877) );
INVxp67_ASAP7_75t_L g933 ( .A(n_851), .Y(n_933) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI222xp33_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_860), .B1(n_861), .B2(n_862), .C1(n_863), .C2(n_866), .Y(n_855) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g924 ( .A(n_859), .Y(n_924) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
OR2x2_ASAP7_75t_L g879 ( .A(n_865), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AOI221x1_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_873), .B1(n_875), .B2(n_878), .C(n_881), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp33_ASAP7_75t_SL g881 ( .A1(n_882), .A2(n_883), .B1(n_885), .B2(n_886), .Y(n_881) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
BUFx3_ASAP7_75t_L g926 ( .A(n_888), .Y(n_926) );
INVx2_ASAP7_75t_L g898 ( .A(n_889), .Y(n_898) );
AOI211xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B(n_894), .C(n_899), .Y(n_890) );
NAND2x1_ASAP7_75t_L g906 ( .A(n_893), .B(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_SL g923 ( .A1(n_897), .A2(n_924), .B1(n_925), .B2(n_927), .Y(n_923) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NAND3xp33_ASAP7_75t_SL g903 ( .A(n_904), .B(n_915), .C(n_928), .Y(n_903) );
O2A1O1Ixp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_908), .B(n_909), .C(n_912), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_919), .B1(n_920), .B2(n_921), .C(n_923), .Y(n_915) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_918), .Y(n_939) );
INVxp67_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_934), .B1(n_935), .B2(n_936), .C(n_940), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_932), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_943), .B(n_947), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_955), .Y(n_945) );
INVx1_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
BUFx12f_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
CKINVDCx11_ASAP7_75t_R g953 ( .A(n_954), .Y(n_953) );
NOR2xp67_ASAP7_75t_R g955 ( .A(n_956), .B(n_957), .Y(n_955) );
BUFx3_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_SL g959 ( .A(n_960), .Y(n_959) );
BUFx4_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
CKINVDCx11_ASAP7_75t_R g964 ( .A(n_965), .Y(n_964) );
endmodule