module fake_netlist_5_342_n_33 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_33);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_33;

wire n_29;
wire n_16;
wire n_12;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_10;
wire n_28;
wire n_24;
wire n_21;
wire n_32;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_26;
wire n_30;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;

BUFx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_2),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_1),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_5),
.B(n_8),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_13),
.C(n_11),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_R g24 ( 
.A(n_22),
.B(n_16),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

AND2x4_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_18),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_29),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_33)
);


endmodule