module real_jpeg_6242_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_1),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_1),
.Y(n_435)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_1),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_2),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_2),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_2),
.B(n_87),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_4),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_4),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_4),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_4),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_4),
.B(n_92),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_4),
.B(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_5),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_5),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_5),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_5),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_5),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_6),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_6),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_6),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_6),
.B(n_70),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_6),
.Y(n_436)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_8),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_8),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_8),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_9),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_9),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_9),
.B(n_76),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_9),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_9),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_9),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_9),
.B(n_384),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_11),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_11),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_11),
.B(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_14),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_14),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_14),
.B(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_15),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_16),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_16),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_16),
.B(n_76),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_16),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_16),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_16),
.B(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_17),
.Y(n_179)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_17),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_17),
.Y(n_384)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_507),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_485),
.B(n_506),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_426),
.B(n_482),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_276),
.B(n_311),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_234),
.B(n_275),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_207),
.B(n_233),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_30),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_162),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_31),
.B(n_162),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_110),
.C(n_146),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_32),
.B(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g521 ( 
.A(n_32),
.Y(n_521)
);

FAx1_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_72),
.CI(n_89),
.CON(n_32),
.SN(n_32)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_33),
.B(n_72),
.C(n_89),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_48),
.C(n_63),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_34),
.B(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_36),
.B(n_40),
.C(n_44),
.Y(n_161)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_39),
.Y(n_226)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_46),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_47),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_48),
.A2(n_63),
.B1(n_64),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_48),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_60),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_49),
.A2(n_60),
.B1(n_184),
.B2(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_49),
.A2(n_216),
.B1(n_224),
.B2(n_255),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_49),
.A2(n_112),
.B1(n_113),
.B2(n_216),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_49),
.B(n_224),
.C(n_282),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_75),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g170 ( 
.A(n_50),
.B(n_171),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_50),
.B(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_51),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_52),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_53),
.B(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_58),
.Y(n_326)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_59),
.Y(n_177)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_59),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_60),
.A2(n_184),
.B1(n_185),
.B2(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_60),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_60),
.B(n_185),
.C(n_190),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g321 ( 
.A(n_62),
.Y(n_321)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_227)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_73),
.A2(n_74),
.B1(n_112),
.B2(n_113),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_73),
.B(n_113),
.C(n_466),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_73),
.A2(n_74),
.B1(n_169),
.B2(n_170),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_73),
.B(n_170),
.C(n_297),
.Y(n_513)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_74),
.B(n_81),
.C(n_86),
.Y(n_198)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_78),
.Y(n_339)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_81),
.A2(n_88),
.B1(n_132),
.B2(n_133),
.Y(n_344)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_91),
.B(n_96),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_90),
.B(n_101),
.C(n_108),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_98),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_99),
.B(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_108),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_105),
.Y(n_360)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_106),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_109),
.B(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_109),
.B(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_109),
.B(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_110),
.B(n_146),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_127),
.C(n_129),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_111),
.A2(n_127),
.B1(n_128),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_126),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_116),
.C(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_113),
.B(n_216),
.C(n_448),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_114),
.Y(n_343)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_121),
.A2(n_122),
.B1(n_242),
.B2(n_247),
.Y(n_241)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_122),
.B(n_243),
.C(n_244),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_129),
.B(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.C(n_142),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_130),
.A2(n_131),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_143),
.Y(n_414)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_161),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_149),
.C(n_161),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_157),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_151),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_151),
.Y(n_296)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_165),
.C(n_206),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_193),
.B1(n_205),
.B2(n_206),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_181),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_167),
.B(n_168),
.C(n_181),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_180),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_169),
.A2(n_170),
.B1(n_251),
.B2(n_252),
.Y(n_515)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_170),
.B(n_272),
.C(n_273),
.Y(n_271)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_174),
.Y(n_272)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_178),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_189),
.B2(n_190),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_185),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_185),
.A2(n_188),
.B1(n_224),
.B2(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_185),
.B(n_224),
.C(n_252),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_185),
.A2(n_188),
.B1(n_336),
.B2(n_337),
.Y(n_354)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_188),
.B(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_189),
.A2(n_190),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_190),
.B(n_433),
.C(n_439),
.Y(n_461)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_192),
.Y(n_294)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_200),
.B(n_202),
.C(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_204),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_231),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_208),
.B(n_231),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.C(n_228),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_209),
.A2(n_210),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_213),
.B(n_228),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.C(n_227),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_214),
.B(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_217),
.B(n_227),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_224),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_333)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_224),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_224),
.A2(n_255),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_235),
.B(n_276),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_277),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_237),
.B(n_277),
.Y(n_425)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_257),
.CI(n_274),
.CON(n_237),
.SN(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_250),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_248),
.B2(n_249),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_249),
.C(n_250),
.Y(n_301)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_256),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_260),
.C(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_271),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_269),
.C(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_270),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_267),
.A2(n_270),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_267),
.B(n_459),
.C(n_461),
.Y(n_489)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_268),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_270),
.B(n_306),
.C(n_309),
.Y(n_444)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_278),
.B(n_280),
.C(n_299),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_299),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_281),
.B(n_289),
.C(n_290),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_297),
.B2(n_298),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_293),
.B(n_296),
.C(n_297),
.Y(n_453)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_297),
.A2(n_298),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_310),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_300),
.B(n_303),
.C(n_305),
.Y(n_478)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

OAI31xp33_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_422),
.A3(n_423),
.B(n_425),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_416),
.B(n_421),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_401),
.B(n_415),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_355),
.B(n_400),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_345),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_316),
.B(n_345),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_334),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_331),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_318),
.B(n_331),
.C(n_334),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.C(n_327),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_347)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_327),
.B(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_340),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_335),
.B(n_410),
.C(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_344),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.C(n_354),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_354),
.B1(n_392),
.B2(n_398),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_394),
.B(n_399),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_380),
.B(n_393),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_365),
.B(n_379),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_376),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_376),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_371),
.B(n_375),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_371),
.Y(n_375)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_375),
.A2(n_382),
.B1(n_387),
.B2(n_388),
.Y(n_381)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_389),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_389),
.Y(n_393)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_383),
.A2(n_385),
.B(n_387),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_391),
.B(n_392),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_396),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_403),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_407),
.B2(n_408),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_409),
.C(n_412),
.Y(n_417)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.Y(n_408)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_418),
.Y(n_421)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_419),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_479),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_427),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_471),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_471),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g524 ( 
.A(n_428),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_445),
.CI(n_455),
.CON(n_428),
.SN(n_428)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_429),
.B(n_445),
.C(n_455),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.C(n_444),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_430),
.A2(n_431),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_444),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_437),
.B1(n_438),
.B2(n_443),
.Y(n_432)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_433),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_433),
.A2(n_443),
.B1(n_515),
.B2(n_516),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

INVx8_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_439),
.Y(n_442)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_453),
.C(n_454),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_446),
.A2(n_447),
.B1(n_476),
.B2(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_452),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_454),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_457),
.B1(n_462),
.B2(n_470),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_463),
.C(n_464),
.Y(n_504)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.C(n_478),
.Y(n_471)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_472),
.B(n_475),
.CI(n_478),
.CON(n_481),
.SN(n_481)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_473),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_481),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_481),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_505),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_505),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_504),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_490),
.C(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_492),
.A2(n_493),
.B1(n_500),
.B2(n_501),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_494),
.Y(n_498)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_497),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_498),
.C(n_500),
.Y(n_511)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_503),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_520),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_519),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_519),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_517),
.B2(n_518),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_513),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_515),
.Y(n_516)
);


endmodule