module fake_aes_10637_n_1169 (n_303, n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_304, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_302, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1169);
input n_303;
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_304;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_302;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1169;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_1128;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_971;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_434;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_599;
wire n_461;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1078;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1024;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_1042;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1160;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1063;
wire n_767;
wire n_828;
wire n_1014;
wire n_1138;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_601;
wire n_439;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_420;
wire n_621;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_716;
wire n_357;
wire n_653;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_947;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_1125;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_1159;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_1069;
wire n_1021;
wire n_972;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_912;
wire n_841;
wire n_1043;
wire n_924;
wire n_1141;
wire n_582;
wire n_378;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1112;
wire n_1075;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_631;
wire n_453;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
INVx1_ASAP7_75t_L g305 ( .A(n_36), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_260), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_27), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_126), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_164), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_34), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_2), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_92), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_31), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_103), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_254), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_87), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_184), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_193), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_45), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_163), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_261), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_152), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_180), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_69), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_145), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_43), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_113), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_223), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_79), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_230), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_233), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_54), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_5), .Y(n_334) );
INVxp33_ASAP7_75t_SL g335 ( .A(n_226), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_243), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_66), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_13), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_210), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_122), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_151), .Y(n_341) );
BUFx2_ASAP7_75t_SL g342 ( .A(n_301), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_253), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_19), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_62), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_120), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_222), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_130), .Y(n_348) );
BUFx2_ASAP7_75t_SL g349 ( .A(n_155), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_192), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_197), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_279), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_201), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_105), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_270), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_304), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_269), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_4), .Y(n_359) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_282), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_121), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_142), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_58), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_189), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_244), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_298), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_76), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_71), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_194), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_131), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_48), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_208), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_81), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_18), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_129), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_23), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_288), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_143), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_206), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_258), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_119), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_157), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_175), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_4), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_118), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_147), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_99), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_7), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_272), .Y(n_389) );
INVxp33_ASAP7_75t_L g390 ( .A(n_198), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_280), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_171), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_196), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_78), .Y(n_394) );
BUFx5_ASAP7_75t_L g395 ( .A(n_271), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_165), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_281), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_75), .Y(n_398) );
INVx4_ASAP7_75t_R g399 ( .A(n_292), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_77), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_265), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_255), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_85), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_297), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_276), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_274), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_273), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_53), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_203), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_228), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_191), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_291), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_286), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_14), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_246), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_278), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_202), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_61), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_225), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_127), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_56), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_283), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_52), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_285), .Y(n_424) );
BUFx2_ASAP7_75t_SL g425 ( .A(n_59), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_290), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_117), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_37), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_153), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_13), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_141), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_159), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_123), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_295), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_186), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_235), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_11), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_72), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_213), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_293), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_289), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_90), .B(n_68), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_104), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_238), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_231), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_88), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_241), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_30), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_181), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_124), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_114), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_190), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_107), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_176), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_220), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_1), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_232), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_252), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_284), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_144), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_110), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_275), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_89), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_287), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_93), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_172), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_95), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_148), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_41), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_299), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_277), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_0), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_239), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_240), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_219), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_374), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_352), .Y(n_477) );
OAI22x1_ASAP7_75t_R g478 ( .A1(n_312), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_478) );
OAI21x1_ASAP7_75t_L g479 ( .A1(n_352), .A2(n_26), .B(n_25), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_458), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_423), .B(n_3), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_448), .B(n_3), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_390), .B(n_315), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_448), .B(n_5), .Y(n_484) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_331), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_472), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_454), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_331), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_454), .B(n_6), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_306), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_414), .B(n_6), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_311), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_395), .Y(n_493) );
INVx6_ASAP7_75t_L g494 ( .A(n_395), .Y(n_494) );
BUFx8_ASAP7_75t_SL g495 ( .A(n_313), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_430), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_348), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_338), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_498) );
NAND2xp33_ASAP7_75t_L g499 ( .A(n_395), .B(n_302), .Y(n_499) );
OAI22x1_ASAP7_75t_L g500 ( .A1(n_334), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_376), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_309), .B(n_12), .Y(n_502) );
OAI22x1_ASAP7_75t_SL g503 ( .A1(n_384), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_344), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_308), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_331), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_495), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_485), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_484), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_493), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_484), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_485), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_487), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_485), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_483), .B(n_400), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_476), .B(n_437), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_477), .B(n_316), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_494), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_480), .Y(n_519) );
INVxp33_ASAP7_75t_L g520 ( .A(n_492), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_488), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_477), .B(n_456), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_504), .B(n_395), .Y(n_524) );
INVx6_ASAP7_75t_L g525 ( .A(n_490), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_505), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_490), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_489), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_486), .B(n_359), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_489), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_496), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_481), .A2(n_388), .B1(n_335), .B2(n_366), .Y(n_532) );
INVx4_ASAP7_75t_L g533 ( .A(n_525), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_525), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_520), .B(n_502), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_510), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_509), .B(n_498), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_523), .A2(n_499), .B(n_479), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_517), .B(n_494), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_520), .B(n_497), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_511), .B(n_527), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_516), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_511), .B(n_491), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_513), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_517), .B(n_491), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_528), .B(n_482), .C(n_498), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_531), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_526), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_526), .Y(n_549) );
O2A1O1Ixp5_ASAP7_75t_L g550 ( .A1(n_524), .A2(n_392), .B(n_360), .C(n_307), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_515), .B(n_501), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_525), .B(n_310), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_530), .A2(n_500), .B1(n_349), .B2(n_425), .Y(n_554) );
NOR2xp33_ASAP7_75t_SL g555 ( .A(n_507), .B(n_393), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_519), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_529), .B(n_314), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_518), .B(n_317), .Y(n_558) );
INVxp33_ASAP7_75t_L g559 ( .A(n_532), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_518), .B(n_318), .Y(n_560) );
NOR2xp33_ASAP7_75t_SL g561 ( .A(n_512), .B(n_405), .Y(n_561) );
INVx8_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_512), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_514), .B(n_501), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_514), .A2(n_342), .B1(n_322), .B2(n_324), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_521), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_521), .B(n_319), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_522), .Y(n_568) );
BUFx2_ASAP7_75t_L g569 ( .A(n_522), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_548), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_545), .B(n_410), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_535), .B(n_428), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_543), .A2(n_327), .B(n_328), .C(n_305), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_559), .B(n_503), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_540), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_548), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_538), .A2(n_347), .B(n_345), .Y(n_577) );
OR2x6_ASAP7_75t_L g578 ( .A(n_552), .B(n_478), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_547), .B(n_460), .Y(n_579) );
BUFx3_ASAP7_75t_L g580 ( .A(n_548), .Y(n_580) );
BUFx2_ASAP7_75t_SL g581 ( .A(n_556), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_542), .B(n_467), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_564), .B(n_330), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_539), .A2(n_358), .B(n_353), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_533), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_564), .B(n_463), .Y(n_586) );
NOR3xp33_ASAP7_75t_L g587 ( .A(n_546), .B(n_363), .C(n_351), .Y(n_587) );
AO21x1_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_362), .B(n_361), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_537), .B(n_15), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_537), .A2(n_442), .B1(n_367), .B2(n_373), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_546), .B(n_365), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_550), .A2(n_382), .B(n_375), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_536), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_551), .A2(n_396), .B(n_391), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_557), .A2(n_401), .B(n_398), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_552), .B(n_370), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_541), .A2(n_411), .B(n_404), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_554), .A2(n_565), .B1(n_534), .B2(n_533), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_553), .A2(n_415), .B(n_413), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_560), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_558), .B(n_444), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_534), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_562), .A2(n_421), .B(n_420), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_563), .A2(n_426), .B(n_424), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_561), .A2(n_431), .B1(n_434), .B2(n_429), .Y(n_606) );
BUFx3_ASAP7_75t_L g607 ( .A(n_569), .Y(n_607) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_561), .B(n_326), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_567), .B(n_445), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_562), .B(n_320), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_562), .A2(n_449), .B(n_447), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_583), .B(n_555), .Y(n_612) );
AO31x2_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_455), .A3(n_459), .B(n_451), .Y(n_613) );
AO31x2_ASAP7_75t_L g614 ( .A1(n_588), .A2(n_466), .A3(n_468), .B(n_462), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_607), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g616 ( .A(n_574), .B(n_582), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_591), .A2(n_566), .B(n_568), .Y(n_617) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_573), .A2(n_475), .A3(n_470), .B(n_364), .Y(n_618) );
AO31x2_ASAP7_75t_L g619 ( .A1(n_595), .A2(n_368), .A3(n_394), .B(n_339), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_575), .B(n_16), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_578), .Y(n_621) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_605), .A2(n_419), .B(n_408), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_570), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_578), .Y(n_624) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_594), .A2(n_469), .B(n_427), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_584), .A2(n_323), .B(n_321), .Y(n_626) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_592), .A2(n_395), .B(n_355), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_601), .A2(n_332), .B(n_325), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_570), .Y(n_629) );
OAI21x1_ASAP7_75t_SL g630 ( .A1(n_604), .A2(n_611), .B(n_606), .Y(n_630) );
OAI21x1_ASAP7_75t_L g631 ( .A1(n_600), .A2(n_355), .B(n_336), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_581), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_586), .B(n_333), .Y(n_633) );
OA21x2_ASAP7_75t_L g634 ( .A1(n_596), .A2(n_587), .B(n_598), .Y(n_634) );
O2A1O1Ixp5_ASAP7_75t_L g635 ( .A1(n_599), .A2(n_399), .B(n_343), .C(n_379), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_571), .B(n_337), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_589), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_579), .A2(n_340), .B1(n_346), .B2(n_341), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_597), .B(n_350), .Y(n_639) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_593), .A2(n_355), .B(n_336), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_572), .B(n_590), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_593), .Y(n_642) );
AND2x6_ASAP7_75t_L g643 ( .A(n_580), .B(n_329), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_609), .B(n_354), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_608), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_602), .B(n_356), .Y(n_646) );
OR2x6_ASAP7_75t_L g647 ( .A(n_585), .B(n_416), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_609), .B(n_387), .C(n_336), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_603), .A2(n_443), .B(n_432), .C(n_438), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_610), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_585), .B(n_357), .Y(n_651) );
OAI21x1_ASAP7_75t_SL g652 ( .A1(n_576), .A2(n_17), .B(n_18), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_585), .B(n_369), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_589), .Y(n_654) );
AOI211x1_ASAP7_75t_L g655 ( .A1(n_588), .A2(n_20), .B(n_17), .C(n_19), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_589), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_589), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_577), .A2(n_432), .B(n_387), .Y(n_658) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_577), .A2(n_432), .B(n_387), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_621), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_641), .A2(n_433), .B1(n_372), .B2(n_377), .C(n_474), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_624), .A2(n_378), .B1(n_380), .B2(n_371), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_650), .A2(n_457), .B1(n_471), .B2(n_438), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_632), .A2(n_383), .B1(n_385), .B2(n_381), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_642), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_637), .B(n_20), .Y(n_666) );
OAI21x1_ASAP7_75t_L g667 ( .A1(n_640), .A2(n_457), .B(n_438), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_655), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_652), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_623), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_615), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_654), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_622), .A2(n_389), .B(n_386), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_656), .Y(n_675) );
AO21x2_ASAP7_75t_L g676 ( .A1(n_617), .A2(n_506), .B(n_488), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_647), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_625), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g679 ( .A1(n_620), .A2(n_441), .A3(n_402), .B1(n_403), .B2(n_406), .Y(n_679) );
OAI21x1_ASAP7_75t_L g680 ( .A1(n_627), .A2(n_471), .B(n_457), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_657), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_612), .B(n_21), .Y(n_682) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_658), .A2(n_471), .B(n_506), .Y(n_683) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_651), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_659), .A2(n_506), .B(n_29), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_647), .Y(n_686) );
OAI21x1_ASAP7_75t_L g687 ( .A1(n_631), .A2(n_32), .B(n_28), .Y(n_687) );
OAI21x1_ASAP7_75t_SL g688 ( .A1(n_630), .A2(n_21), .B(n_22), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_614), .Y(n_689) );
AO31x2_ASAP7_75t_L g690 ( .A1(n_649), .A2(n_22), .A3(n_23), .B(n_24), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_614), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_635), .A2(n_634), .B(n_648), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_645), .B(n_24), .Y(n_693) );
BUFx3_ASAP7_75t_L g694 ( .A(n_643), .Y(n_694) );
OAI21x1_ASAP7_75t_L g695 ( .A1(n_629), .A2(n_33), .B(n_35), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_619), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_616), .A2(n_439), .B1(n_473), .B2(n_465), .Y(n_697) );
OA21x2_ASAP7_75t_L g698 ( .A1(n_626), .A2(n_407), .B(n_397), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_613), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_634), .B(n_409), .Y(n_700) );
OAI21x1_ASAP7_75t_L g701 ( .A1(n_653), .A2(n_38), .B(n_39), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_646), .A2(n_440), .B(n_464), .C(n_461), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_643), .Y(n_703) );
OA21x2_ASAP7_75t_L g704 ( .A1(n_628), .A2(n_417), .B(n_412), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_613), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_643), .Y(n_706) );
OAI21x1_ASAP7_75t_L g707 ( .A1(n_636), .A2(n_40), .B(n_42), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_638), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_618), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_618), .Y(n_710) );
AO21x2_ASAP7_75t_L g711 ( .A1(n_633), .A2(n_508), .B(n_44), .Y(n_711) );
INVx2_ASAP7_75t_SL g712 ( .A(n_644), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_639), .A2(n_422), .B(n_418), .Y(n_713) );
OR2x6_ASAP7_75t_L g714 ( .A(n_624), .B(n_508), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_650), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_641), .B(n_435), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_650), .Y(n_717) );
OAI21x1_ASAP7_75t_L g718 ( .A1(n_640), .A2(n_46), .B(n_47), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_621), .Y(n_719) );
OAI21x1_ASAP7_75t_SL g720 ( .A1(n_630), .A2(n_49), .B(n_50), .Y(n_720) );
NOR2x1_ASAP7_75t_SL g721 ( .A(n_647), .B(n_51), .Y(n_721) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_640), .A2(n_55), .B(n_57), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_694), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_699), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_715), .B(n_436), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_665), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_677), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_705), .Y(n_728) );
OR2x6_ASAP7_75t_L g729 ( .A(n_693), .B(n_60), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_689), .Y(n_730) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_668), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_691), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_673), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_717), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_675), .Y(n_735) );
BUFx2_ASAP7_75t_SL g736 ( .A(n_703), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_681), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_693), .B(n_446), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_668), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_672), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_671), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_666), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_712), .B(n_450), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_706), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_669), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_682), .Y(n_746) );
INVx3_ASAP7_75t_L g747 ( .A(n_714), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_684), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_708), .B(n_452), .Y(n_749) );
BUFx3_ASAP7_75t_L g750 ( .A(n_660), .Y(n_750) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_692), .A2(n_453), .B(n_508), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_686), .B(n_63), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_688), .Y(n_753) );
BUFx6f_ASAP7_75t_L g754 ( .A(n_714), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_709), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_716), .B(n_64), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_710), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_696), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_721), .Y(n_759) );
AO31x2_ASAP7_75t_L g760 ( .A1(n_700), .A2(n_65), .A3(n_67), .B(n_70), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_690), .Y(n_761) );
INVx4_ASAP7_75t_L g762 ( .A(n_719), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_679), .B(n_73), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_690), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_690), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_670), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_714), .B(n_74), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_704), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_704), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_698), .Y(n_770) );
OAI21x1_ASAP7_75t_L g771 ( .A1(n_680), .A2(n_80), .B(n_82), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_678), .Y(n_772) );
HB1xp67_ASAP7_75t_SL g773 ( .A(n_661), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_674), .A2(n_83), .B(n_84), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_695), .Y(n_775) );
AO21x1_ASAP7_75t_L g776 ( .A1(n_674), .A2(n_86), .B(n_91), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_662), .B(n_94), .Y(n_777) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_698), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_720), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_701), .Y(n_780) );
INVx3_ASAP7_75t_L g781 ( .A(n_722), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_718), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_713), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_707), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_687), .Y(n_785) );
AO21x2_ASAP7_75t_L g786 ( .A1(n_692), .A2(n_96), .B(n_97), .Y(n_786) );
BUFx10_ASAP7_75t_L g787 ( .A(n_679), .Y(n_787) );
INVx8_ASAP7_75t_L g788 ( .A(n_664), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_711), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_676), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_676), .Y(n_791) );
AO21x2_ASAP7_75t_L g792 ( .A1(n_711), .A2(n_98), .B(n_100), .Y(n_792) );
INVx3_ASAP7_75t_L g793 ( .A(n_685), .Y(n_793) );
OAI21xp5_ASAP7_75t_L g794 ( .A1(n_663), .A2(n_101), .B(n_102), .Y(n_794) );
BUFx3_ASAP7_75t_L g795 ( .A(n_683), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_702), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_697), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_677), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_699), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_715), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_660), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_715), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_715), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_694), .B(n_106), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_715), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_677), .Y(n_806) );
INVx4_ASAP7_75t_SL g807 ( .A(n_694), .Y(n_807) );
CKINVDCx6p67_ASAP7_75t_R g808 ( .A(n_694), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_715), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_699), .Y(n_810) );
INVx4_ASAP7_75t_L g811 ( .A(n_706), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_667), .A2(n_108), .B(n_109), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_672), .Y(n_813) );
INVx5_ASAP7_75t_L g814 ( .A(n_694), .Y(n_814) );
AOI21xp33_ASAP7_75t_L g815 ( .A1(n_779), .A2(n_111), .B(n_112), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_726), .Y(n_816) );
BUFx3_ASAP7_75t_L g817 ( .A(n_750), .Y(n_817) );
INVx2_ASAP7_75t_SL g818 ( .A(n_727), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_748), .B(n_115), .Y(n_819) );
OR2x2_ASAP7_75t_L g820 ( .A(n_740), .B(n_300), .Y(n_820) );
INVx4_ASAP7_75t_L g821 ( .A(n_729), .Y(n_821) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_754), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_734), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_800), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_802), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_803), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_805), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_733), .B(n_116), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_809), .B(n_125), .Y(n_829) );
BUFx2_ASAP7_75t_L g830 ( .A(n_813), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_735), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_737), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_729), .B(n_128), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_787), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_745), .B(n_135), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_758), .Y(n_836) );
INVxp67_ASAP7_75t_L g837 ( .A(n_778), .Y(n_837) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_724), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_724), .B(n_136), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_787), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_725), .B(n_140), .Y(n_841) );
BUFx3_ASAP7_75t_L g842 ( .A(n_798), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_728), .Y(n_843) );
INVxp33_ASAP7_75t_L g844 ( .A(n_806), .Y(n_844) );
INVx2_ASAP7_75t_R g845 ( .A(n_795), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_728), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_799), .Y(n_847) );
NOR2x1_ASAP7_75t_L g848 ( .A(n_759), .B(n_146), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_797), .B(n_149), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_799), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_738), .B(n_150), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_743), .B(n_154), .Y(n_852) );
INVx1_ASAP7_75t_SL g853 ( .A(n_736), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_746), .B(n_156), .Y(n_854) );
BUFx2_ASAP7_75t_L g855 ( .A(n_731), .Y(n_855) );
INVx1_ASAP7_75t_SL g856 ( .A(n_736), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_810), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_810), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_730), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_730), .B(n_158), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_732), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_742), .B(n_160), .Y(n_862) );
INVx3_ASAP7_75t_L g863 ( .A(n_767), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_752), .B(n_161), .Y(n_864) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_772), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_755), .B(n_162), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_741), .B(n_166), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_741), .B(n_167), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_783), .B(n_168), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_757), .Y(n_870) );
BUFx2_ASAP7_75t_L g871 ( .A(n_731), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_766), .Y(n_872) );
OR2x2_ASAP7_75t_L g873 ( .A(n_739), .B(n_169), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_749), .B(n_170), .Y(n_874) );
CKINVDCx6p67_ASAP7_75t_R g875 ( .A(n_762), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_739), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_753), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_768), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_747), .B(n_173), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_744), .B(n_174), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_723), .B(n_177), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_769), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_761), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_723), .B(n_178), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_808), .B(n_179), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_765), .B(n_182), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_773), .B(n_183), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_796), .B(n_185), .Y(n_888) );
NOR2x1_ASAP7_75t_L g889 ( .A(n_811), .B(n_187), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_770), .B(n_188), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_767), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_764), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_762), .B(n_195), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_747), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_760), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_754), .Y(n_896) );
INVx1_ASAP7_75t_SL g897 ( .A(n_754), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_756), .B(n_199), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_804), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_807), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_807), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_811), .B(n_200), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_790), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_779), .Y(n_904) );
AND2x4_ASAP7_75t_L g905 ( .A(n_814), .B(n_204), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_763), .B(n_205), .Y(n_906) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_790), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_801), .B(n_296), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_814), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_781), .Y(n_910) );
BUFx3_ASAP7_75t_L g911 ( .A(n_814), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_788), .B(n_207), .Y(n_912) );
INVxp67_ASAP7_75t_SL g913 ( .A(n_791), .Y(n_913) );
INVx4_ASAP7_75t_L g914 ( .A(n_788), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_777), .B(n_209), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_776), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_SL g917 ( .A1(n_774), .A2(n_789), .B(n_793), .C(n_782), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_784), .B(n_211), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_751), .B(n_212), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_836), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_830), .B(n_791), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_836), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_823), .B(n_751), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_824), .B(n_780), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_816), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_825), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_826), .B(n_792), .Y(n_927) );
NAND2xp33_ASAP7_75t_R g928 ( .A(n_863), .B(n_789), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_872), .B(n_785), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_827), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_831), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_832), .B(n_786), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_870), .Y(n_933) );
INVx3_ASAP7_75t_L g934 ( .A(n_853), .Y(n_934) );
OR2x2_ASAP7_75t_L g935 ( .A(n_838), .B(n_775), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_838), .B(n_794), .Y(n_936) );
INVx2_ASAP7_75t_SL g937 ( .A(n_817), .Y(n_937) );
BUFx3_ASAP7_75t_L g938 ( .A(n_911), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_853), .B(n_214), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_883), .Y(n_940) );
NOR2x1_ASAP7_75t_L g941 ( .A(n_821), .B(n_771), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_861), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_903), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_850), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_856), .B(n_215), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_861), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_856), .B(n_216), .Y(n_947) );
INVx1_ASAP7_75t_SL g948 ( .A(n_855), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_843), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_857), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_896), .B(n_217), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_903), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_846), .Y(n_953) );
NOR2xp67_ASAP7_75t_L g954 ( .A(n_821), .B(n_218), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_847), .Y(n_955) );
NAND3xp33_ASAP7_75t_L g956 ( .A(n_887), .B(n_812), .C(n_221), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_858), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_859), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_877), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_914), .B(n_224), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_907), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_914), .B(n_227), .Y(n_962) );
INVxp67_ASAP7_75t_SL g963 ( .A(n_865), .Y(n_963) );
INVx3_ASAP7_75t_L g964 ( .A(n_863), .Y(n_964) );
INVx3_ASAP7_75t_L g965 ( .A(n_822), .Y(n_965) );
AND2x4_ASAP7_75t_L g966 ( .A(n_904), .B(n_229), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_878), .B(n_234), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_899), .B(n_236), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_897), .B(n_842), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_882), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_894), .B(n_237), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_907), .B(n_242), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_839), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_876), .Y(n_974) );
INVx2_ASAP7_75t_SL g975 ( .A(n_875), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_891), .B(n_245), .Y(n_976) );
BUFx2_ASAP7_75t_L g977 ( .A(n_871), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_839), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_844), .B(n_247), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_833), .A2(n_248), .B1(n_249), .B2(n_250), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_860), .Y(n_981) );
HB1xp67_ASAP7_75t_L g982 ( .A(n_837), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_837), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_892), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_913), .B(n_251), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_819), .B(n_256), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_822), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_869), .B(n_257), .Y(n_988) );
INVx1_ASAP7_75t_SL g989 ( .A(n_909), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_849), .B(n_259), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_913), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_860), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_912), .B(n_262), .Y(n_993) );
INVx2_ASAP7_75t_L g994 ( .A(n_910), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_818), .B(n_263), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_829), .B(n_264), .Y(n_996) );
AND2x4_ASAP7_75t_L g997 ( .A(n_900), .B(n_266), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_866), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_820), .B(n_267), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_828), .B(n_268), .Y(n_1000) );
INVxp67_ASAP7_75t_L g1001 ( .A(n_920), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_920), .B(n_901), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_933), .B(n_916), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_969), .B(n_845), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_937), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_989), .B(n_880), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_922), .B(n_886), .Y(n_1007) );
AND2x4_ASAP7_75t_SL g1008 ( .A(n_975), .B(n_885), .Y(n_1008) );
INVxp67_ASAP7_75t_L g1009 ( .A(n_922), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_950), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_948), .B(n_895), .Y(n_1011) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_964), .B(n_905), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_950), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_926), .B(n_886), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_977), .B(n_902), .Y(n_1015) );
NAND2xp67_ASAP7_75t_L g1016 ( .A(n_960), .B(n_915), .Y(n_1016) );
INVx4_ASAP7_75t_L g1017 ( .A(n_938), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_934), .B(n_879), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_921), .B(n_918), .Y(n_1019) );
INVxp67_ASAP7_75t_SL g1020 ( .A(n_963), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_934), .B(n_879), .Y(n_1021) );
INVx4_ASAP7_75t_L g1022 ( .A(n_938), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_982), .B(n_851), .Y(n_1023) );
BUFx2_ASAP7_75t_SL g1024 ( .A(n_954), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_982), .B(n_862), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_983), .B(n_918), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_991), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_983), .B(n_854), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_930), .B(n_874), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_970), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_931), .B(n_868), .Y(n_1031) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_995), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_974), .B(n_867), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_963), .B(n_866), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_953), .B(n_835), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_940), .Y(n_1036) );
INVxp67_ASAP7_75t_L g1037 ( .A(n_943), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_958), .B(n_835), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_959), .B(n_906), .Y(n_1039) );
NAND2x1p5_ASAP7_75t_L g1040 ( .A(n_962), .B(n_905), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_944), .B(n_881), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_943), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_940), .Y(n_1043) );
AND2x4_ASAP7_75t_SL g1044 ( .A(n_997), .B(n_893), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_925), .B(n_884), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_964), .B(n_919), .Y(n_1046) );
NOR2x1_ASAP7_75t_L g1047 ( .A(n_941), .B(n_889), .Y(n_1047) );
OA211x2_ASAP7_75t_L g1048 ( .A1(n_979), .A2(n_840), .B(n_834), .C(n_908), .Y(n_1048) );
NAND2x1p5_ASAP7_75t_L g1049 ( .A(n_954), .B(n_864), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_949), .B(n_852), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_942), .B(n_890), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_955), .Y(n_1052) );
NAND4xp25_ASAP7_75t_L g1053 ( .A(n_956), .B(n_840), .C(n_834), .D(n_841), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_957), .B(n_890), .Y(n_1054) );
AND2x4_ASAP7_75t_SL g1055 ( .A(n_997), .B(n_898), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_952), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1030), .Y(n_1057) );
OAI21xp33_ASAP7_75t_L g1058 ( .A1(n_1016), .A2(n_1053), .B(n_1020), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_1042), .B(n_952), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1004), .B(n_961), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1030), .Y(n_1061) );
OAI21xp33_ASAP7_75t_L g1062 ( .A1(n_1053), .A2(n_980), .B(n_956), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1015), .B(n_923), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1001), .B(n_946), .Y(n_1064) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_1009), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1052), .Y(n_1066) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_1005), .Y(n_1067) );
INVx1_ASAP7_75t_SL g1068 ( .A(n_1017), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1002), .B(n_927), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1056), .Y(n_1070) );
NAND2xp5_ASAP7_75t_SL g1071 ( .A(n_1017), .B(n_936), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1052), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1003), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1037), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1002), .B(n_932), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1036), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_1026), .B(n_929), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1036), .Y(n_1078) );
INVxp67_ASAP7_75t_L g1079 ( .A(n_1006), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_1034), .B(n_984), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1023), .B(n_994), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_1048), .A2(n_973), .B1(n_981), .B2(n_992), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1043), .Y(n_1083) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_1022), .Y(n_1084) );
INVxp67_ASAP7_75t_SL g1085 ( .A(n_1022), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_1007), .B(n_935), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_1008), .B(n_1055), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_1011), .B(n_924), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1050), .B(n_998), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1027), .Y(n_1090) );
INVx2_ASAP7_75t_SL g1091 ( .A(n_1068), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1068), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1088), .B(n_1018), .Y(n_1093) );
OAI322xp33_ASAP7_75t_L g1094 ( .A1(n_1079), .A2(n_1039), .A3(n_1019), .B1(n_1051), .B2(n_1054), .C1(n_1038), .C2(n_1035), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1059), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_1077), .B(n_1043), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1076), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1098 ( .A(n_1085), .B(n_1012), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1057), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1084), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1084), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1061), .Y(n_1102) );
INVxp67_ASAP7_75t_L g1103 ( .A(n_1065), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1066), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1072), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1086), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1064), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1078), .Y(n_1108) );
NOR2x1p5_ASAP7_75t_SL g1109 ( .A(n_1074), .B(n_1010), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1088), .B(n_1021), .Y(n_1110) );
AOI32xp33_ASAP7_75t_L g1111 ( .A1(n_1058), .A2(n_1044), .A3(n_1047), .B1(n_1012), .B2(n_1032), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_1103), .A2(n_1058), .B1(n_1062), .B2(n_1082), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_1094), .B(n_1087), .Y(n_1113) );
AOI21xp5_ASAP7_75t_L g1114 ( .A1(n_1111), .A2(n_1062), .B(n_1071), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1097), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1096), .B(n_1080), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1097), .Y(n_1117) );
NAND2x1_ASAP7_75t_L g1118 ( .A(n_1098), .B(n_1047), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_1098), .A2(n_1067), .B1(n_1040), .B2(n_1049), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1108), .Y(n_1120) );
OAI21xp5_ASAP7_75t_SL g1121 ( .A1(n_1091), .A2(n_980), .B(n_993), .Y(n_1121) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_1092), .Y(n_1122) );
OAI322xp33_ASAP7_75t_L g1123 ( .A1(n_1107), .A2(n_1073), .A3(n_1089), .B1(n_1083), .B2(n_1070), .C1(n_979), .C2(n_1063), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1108), .Y(n_1124) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_1093), .B(n_1069), .Y(n_1125) );
O2A1O1Ixp33_ASAP7_75t_L g1126 ( .A1(n_1114), .A2(n_1101), .B(n_1100), .C(n_1095), .Y(n_1126) );
NOR3xp33_ASAP7_75t_L g1127 ( .A(n_1113), .B(n_848), .C(n_972), .Y(n_1127) );
NAND2xp5_ASAP7_75t_SL g1128 ( .A(n_1112), .B(n_1090), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_1123), .A2(n_1106), .B1(n_1105), .B2(n_1104), .C(n_1102), .Y(n_1129) );
NAND3xp33_ASAP7_75t_L g1130 ( .A(n_1121), .B(n_1099), .C(n_972), .Y(n_1130) );
A2O1A1Ixp33_ASAP7_75t_L g1131 ( .A1(n_1118), .A2(n_1109), .B(n_1110), .C(n_1075), .Y(n_1131) );
OAI221xp5_ASAP7_75t_SL g1132 ( .A1(n_1122), .A2(n_1029), .B1(n_1028), .B2(n_1025), .C(n_1048), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1119), .A2(n_1024), .B1(n_1081), .B2(n_1060), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1115), .Y(n_1134) );
AOI322xp5_ASAP7_75t_L g1135 ( .A1(n_1125), .A2(n_1031), .A3(n_1046), .B1(n_978), .B2(n_1041), .C1(n_1045), .C2(n_1014), .Y(n_1135) );
NOR3xp33_ASAP7_75t_L g1136 ( .A(n_1132), .B(n_1126), .C(n_1127), .Y(n_1136) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_1129), .B(n_1124), .C(n_1120), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1134), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1135), .B(n_1117), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1128), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1130), .Y(n_1141) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_1133), .B(n_1116), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1141), .B(n_1131), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1142), .B(n_1033), .Y(n_1144) );
NOR3x1_ASAP7_75t_L g1145 ( .A(n_1140), .B(n_986), .C(n_917), .Y(n_1145) );
NOR2xp67_ASAP7_75t_L g1146 ( .A(n_1137), .B(n_965), .Y(n_1146) );
AND4x2_ASAP7_75t_L g1147 ( .A(n_1136), .B(n_928), .C(n_999), .D(n_988), .Y(n_1147) );
NOR3xp33_ASAP7_75t_L g1148 ( .A(n_1143), .B(n_1139), .C(n_1138), .Y(n_1148) );
NOR2x1_ASAP7_75t_L g1149 ( .A(n_1146), .B(n_939), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1150 ( .A(n_1144), .B(n_1013), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1145), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1150), .Y(n_1152) );
CKINVDCx20_ASAP7_75t_R g1153 ( .A(n_1151), .Y(n_1153) );
NOR2x1_ASAP7_75t_L g1154 ( .A(n_1149), .B(n_1147), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1152), .Y(n_1155) );
XOR2xp5_ASAP7_75t_L g1156 ( .A(n_1153), .B(n_1148), .Y(n_1156) );
AOI222xp33_ASAP7_75t_L g1157 ( .A1(n_1154), .A2(n_945), .B1(n_947), .B2(n_966), .C1(n_985), .C2(n_951), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1155), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1156), .B(n_1013), .Y(n_1159) );
XOR2xp5_ASAP7_75t_L g1160 ( .A(n_1157), .B(n_990), .Y(n_1160) );
AOI21xp5_ASAP7_75t_L g1161 ( .A1(n_1158), .A2(n_971), .B(n_967), .Y(n_1161) );
AOI22xp5_ASAP7_75t_L g1162 ( .A1(n_1159), .A2(n_996), .B1(n_968), .B2(n_1000), .Y(n_1162) );
AOI21xp5_ASAP7_75t_L g1163 ( .A1(n_1160), .A2(n_971), .B(n_967), .Y(n_1163) );
AOI21xp33_ASAP7_75t_SL g1164 ( .A1(n_1162), .A2(n_1163), .B(n_1161), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_1163), .A2(n_965), .B1(n_976), .B2(n_987), .Y(n_1165) );
INVxp33_ASAP7_75t_L g1166 ( .A(n_1164), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1166), .B(n_1165), .Y(n_1167) );
OA21x2_ASAP7_75t_L g1168 ( .A1(n_1167), .A2(n_815), .B(n_985), .Y(n_1168) );
AOI21xp5_ASAP7_75t_L g1169 ( .A1(n_1168), .A2(n_873), .B(n_888), .Y(n_1169) );
endmodule