module real_jpeg_7114_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_1),
.A2(n_91),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_1),
.A2(n_91),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_3),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_4),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_113),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_5),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_5),
.A2(n_86),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_5),
.A2(n_86),
.B1(n_251),
.B2(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_5),
.A2(n_86),
.B1(n_161),
.B2(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_7),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_7),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_8),
.A2(n_46),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_8),
.B(n_253),
.C(n_257),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_8),
.B(n_71),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_8),
.B(n_209),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_8),
.B(n_96),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_8),
.B(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_11),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_12),
.A2(n_188),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_13),
.A2(n_158),
.B1(n_159),
.B2(n_163),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_13),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_13),
.A2(n_163),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_14),
.Y(n_127)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_14),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_15),
.A2(n_52),
.B1(n_116),
.B2(n_121),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_15),
.A2(n_52),
.B1(n_142),
.B2(n_182),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_15),
.A2(n_52),
.B1(n_171),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_232),
.B1(n_233),
.B2(n_357),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_18),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_231),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_193),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_20),
.B(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_131),
.C(n_177),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_21),
.B(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_56),
.B2(n_130),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_22),
.B(n_57),
.C(n_94),
.Y(n_210)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_41),
.B(n_49),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_24),
.B(n_51),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_27),
.Y(n_139)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_32),
.B(n_46),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_32)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_33),
.Y(n_141)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_36),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_36),
.Y(n_143)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_42),
.Y(n_138)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_46),
.A2(n_146),
.B(n_267),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_46),
.A2(n_92),
.B(n_321),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_47),
.A2(n_135),
.A3(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_55),
.Y(n_225)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_94),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_81),
.B1(n_87),
.B2(n_88),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_58),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_71),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_64),
.Y(n_323)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_70),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_71),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_77),
.B2(n_80),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_73),
.Y(n_335)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_76),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_76),
.Y(n_251)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_79),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_79),
.Y(n_276)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_79),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_79),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_81),
.A2(n_87),
.B(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_82),
.Y(n_331)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_87),
.B(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_88),
.Y(n_229)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_107),
.B(n_114),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_95),
.A2(n_107),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_95),
.A2(n_197),
.B1(n_273),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_96),
.B(n_115),
.Y(n_247)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_97),
.A2(n_114),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_103),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_103),
.Y(n_269)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_104),
.Y(n_284)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVx5_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_111),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_123),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_127),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_131),
.A2(n_132),
.B1(n_177),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_144),
.B2(n_145),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_134),
.B(n_144),
.Y(n_214)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_156),
.B1(n_164),
.B2(n_167),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_146),
.A2(n_262),
.B(n_267),
.Y(n_261)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_157),
.B1(n_185),
.B2(n_189),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_168),
.B1(n_203),
.B2(n_208),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_147),
.B(n_268),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_147),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_158),
.Y(n_266)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_165),
.B(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_172),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_177),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.C(n_192),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_178),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_183),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_183),
.A2(n_230),
.B(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_184),
.B(n_192),
.Y(n_348)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_185),
.Y(n_326)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_190),
.A2(n_289),
.B(n_292),
.Y(n_288)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_213),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_240),
.B(n_247),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_197),
.A2(n_247),
.B(n_313),
.Y(n_345)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_227),
.B2(n_228),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_225),
.B(n_226),
.Y(n_217)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_351),
.B(n_356),
.Y(n_233)
);

AO21x1_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_340),
.B(n_350),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_307),
.B(n_339),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_279),
.B(n_306),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_260),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_238),
.B(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_248),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_239),
.A2(n_248),
.B1(n_249),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_239),
.Y(n_304)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_270),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_271),
.C(n_278),
.Y(n_308)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_277),
.B2(n_278),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_295),
.B(n_305),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_287),
.B(n_294),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_293),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_303),
.Y(n_305)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_309),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_324),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_318),
.B2(n_319),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_318),
.C(n_324),
.Y(n_341)
);

INVx3_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI32xp33_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_331),
.A3(n_332),
.B1(n_334),
.B2(n_336),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_330),
.Y(n_346)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_341),
.B(n_342),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_349),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_346),
.C(n_349),
.Y(n_352)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_352),
.B(n_353),
.Y(n_356)
);


endmodule