module fake_jpeg_27564_n_241 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx12f_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_0),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_61),
.B(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_25),
.B(n_32),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_20),
.B(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_70),
.Y(n_105)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_26),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_26),
.B1(n_19),
.B2(n_31),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_80),
.B1(n_83),
.B2(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_79),
.Y(n_110)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_30),
.B1(n_27),
.B2(n_34),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_113),
.B(n_0),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_73),
.B1(n_65),
.B2(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_141)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_65),
.B1(n_75),
.B2(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_117),
.B1(n_25),
.B2(n_1),
.Y(n_118)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_102),
.Y(n_121)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_106),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_38),
.C(n_18),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_34),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_114),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_38),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_81),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_53),
.B1(n_21),
.B2(n_25),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_118),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_129),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_136),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_2),
.B(n_3),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_134),
.B(n_13),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_11),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_11),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_100),
.B1(n_117),
.B2(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_154),
.B1(n_162),
.B2(n_166),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_158),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_106),
.C(n_89),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_157),
.C(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_153),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_93),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_109),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_113),
.C(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_110),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_107),
.B1(n_88),
.B2(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_165),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_170),
.C(n_176),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_122),
.C(n_129),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_136),
.C(n_126),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_151),
.C(n_146),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_182),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_178),
.B1(n_144),
.B2(n_156),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_134),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_118),
.B1(n_138),
.B2(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_143),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_113),
.C(n_140),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_188),
.B(n_167),
.C(n_144),
.D(n_146),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_152),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_201),
.B(n_203),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_153),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_164),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_114),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_215),
.C(n_193),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_184),
.B(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_174),
.B1(n_187),
.B2(n_177),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_212),
.B1(n_191),
.B2(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_187),
.B1(n_177),
.B2(n_183),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_170),
.B(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_172),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_204),
.C(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_210),
.C(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_195),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_205),
.C(n_213),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_95),
.Y(n_222)
);

NAND2x1_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_14),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_228),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_222),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_223),
.B1(n_226),
.B2(n_213),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_224),
.B(n_115),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_228),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_237),
.A2(n_231),
.B(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_238),
.C(n_236),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_127),
.Y(n_241)
);


endmodule