module fake_jpeg_12787_n_410 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_72),
.Y(n_116)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_60),
.B(n_62),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_63),
.B(n_74),
.Y(n_114)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_65),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_0),
.CON(n_66),
.SN(n_66)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_100),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_109),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_8),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_8),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_77),
.B(n_96),
.Y(n_125)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_33),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_92),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_31),
.B(n_0),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_86),
.B(n_102),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_87),
.Y(n_179)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_1),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_104),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_28),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_26),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_107),
.Y(n_138)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_28),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_110),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_1),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_42),
.B1(n_44),
.B2(n_30),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_115),
.A2(n_131),
.B1(n_140),
.B2(n_141),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_54),
.A2(n_42),
.B1(n_44),
.B2(n_32),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_117),
.A2(n_132),
.B1(n_146),
.B2(n_161),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_51),
.B1(n_49),
.B2(n_38),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_128),
.A2(n_153),
.B1(n_160),
.B2(n_177),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_133),
.B(n_118),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_50),
.B1(n_41),
.B2(n_52),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_52),
.B1(n_35),
.B2(n_22),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_114),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_45),
.B1(n_2),
.B2(n_3),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_112),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_94),
.B1(n_79),
.B2(n_68),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_169),
.B1(n_180),
.B2(n_157),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_67),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_73),
.B(n_83),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_66),
.A2(n_3),
.B1(n_6),
.B2(n_89),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_81),
.B(n_6),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_103),
.A2(n_6),
.B1(n_104),
.B2(n_109),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_71),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_170),
.B(n_176),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_58),
.A2(n_27),
.B1(n_53),
.B2(n_47),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_178),
.B1(n_169),
.B2(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_60),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_54),
.A2(n_59),
.B1(n_17),
.B2(n_36),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_58),
.A2(n_27),
.B1(n_53),
.B2(n_47),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_125),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_181),
.B(n_192),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_162),
.B(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_182),
.B(n_187),
.C(n_215),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_183),
.B(n_201),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_166),
.C(n_116),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_202),
.Y(n_240)
);

OR2x2_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_133),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_186),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_189),
.A2(n_212),
.B1(n_213),
.B2(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_123),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_194),
.B(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_147),
.B(n_160),
.C(n_153),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_196),
.A2(n_218),
.B(n_210),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_138),
.A2(n_119),
.B(n_121),
.C(n_168),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_197),
.A2(n_221),
.B(n_232),
.C(n_225),
.Y(n_272)
);

NAND2x1_ASAP7_75t_SL g198 ( 
.A(n_147),
.B(n_113),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_198),
.Y(n_243)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_199),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_136),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_229),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_113),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_205),
.B(n_207),
.Y(n_249)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_143),
.B(n_165),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_214),
.Y(n_275)
);

BUFx12_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_172),
.B1(n_157),
.B2(n_135),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_134),
.A2(n_167),
.B1(n_165),
.B2(n_129),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_122),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_127),
.C(n_120),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_137),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_226),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_135),
.A2(n_129),
.B1(n_122),
.B2(n_151),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

BUFx24_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_163),
.B(n_120),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_220),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_127),
.B(n_163),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_126),
.B(n_151),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_231),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_124),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_206),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_124),
.A2(n_169),
.B1(n_180),
.B2(n_59),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_234),
.A2(n_238),
.B1(n_228),
.B2(n_223),
.Y(n_276)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_149),
.B(n_162),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_186),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_114),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_169),
.A2(n_180),
.B1(n_54),
.B2(n_59),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_230),
.B1(n_208),
.B2(n_196),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_239),
.A2(n_253),
.B1(n_265),
.B2(n_267),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_222),
.B(n_188),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_246),
.A2(n_254),
.B(n_270),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_194),
.B(n_182),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_209),
.B(n_193),
.C(n_211),
.D(n_191),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_187),
.A2(n_218),
.B1(n_182),
.B2(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_187),
.A2(n_236),
.B1(n_229),
.B2(n_204),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_185),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_269),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_215),
.B1(n_181),
.B2(n_203),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_197),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_213),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_235),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_195),
.B1(n_224),
.B2(n_219),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_221),
.B(n_214),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_280),
.A2(n_291),
.B(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_286),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_199),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_256),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_290),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_190),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_248),
.B1(n_278),
.B2(n_261),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_264),
.B(n_233),
.CI(n_209),
.CON(n_290),
.SN(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_271),
.B(n_241),
.C(n_245),
.D(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_277),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_298),
.B(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_269),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_241),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_275),
.B(n_244),
.C(n_240),
.D(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_265),
.B(n_267),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_249),
.A2(n_272),
.B(n_243),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_SL g301 ( 
.A(n_254),
.B(n_246),
.C(n_270),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_276),
.C(n_257),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_239),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_305),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_279),
.B(n_243),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_270),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_251),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_248),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_274),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_301),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_268),
.C(n_261),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_331),
.C(n_285),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_323),
.Y(n_337)
);

AO22x1_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_260),
.B1(n_273),
.B2(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_258),
.B1(n_259),
.B2(n_263),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_299),
.A2(n_259),
.B1(n_262),
.B2(n_251),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_287),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_285),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_293),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_334),
.B(n_336),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_316),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_335),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_288),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_339),
.B(n_321),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_347),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_280),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_342),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_294),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_344),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_307),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_346),
.A2(n_330),
.B1(n_311),
.B2(n_326),
.Y(n_364)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_350),
.C(n_327),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_323),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_349),
.B(n_351),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_305),
.C(n_283),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_284),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_314),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_357),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_321),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_362),
.C(n_363),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_351),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_312),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_328),
.Y(n_366)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_352),
.A2(n_342),
.B(n_330),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_374),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_363),
.B(n_351),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_356),
.Y(n_379)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_358),
.Y(n_370)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_335),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_372),
.B(n_375),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_303),
.B(n_340),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_SL g375 ( 
.A1(n_355),
.A2(n_311),
.A3(n_292),
.B1(n_298),
.B2(n_282),
.C1(n_290),
.C2(n_308),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_358),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_377),
.Y(n_385)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_365),
.B(n_366),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_376),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_361),
.C(n_362),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_387),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_371),
.A2(n_360),
.B(n_342),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_383),
.A2(n_369),
.B1(n_370),
.B2(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_390),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_283),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_380),
.A2(n_381),
.B1(n_369),
.B2(n_365),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_378),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_391),
.A2(n_385),
.B(n_353),
.Y(n_396)
);

AOI21xp33_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_367),
.B(n_368),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_393),
.A2(n_309),
.B(n_338),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_381),
.Y(n_395)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_396),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_376),
.C(n_357),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_392),
.C(n_389),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_400),
.Y(n_403)
);

AOI322xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_402),
.A3(n_404),
.B1(n_403),
.B2(n_395),
.C1(n_398),
.C2(n_391),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_SL g407 ( 
.A(n_405),
.B(n_406),
.C(n_337),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_388),
.A3(n_359),
.B1(n_347),
.B2(n_345),
.C1(n_341),
.C2(n_313),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_332),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_319),
.Y(n_410)
);


endmodule