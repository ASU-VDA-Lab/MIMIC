module fake_jpeg_5729_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_28),
.B1(n_31),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_59),
.B1(n_42),
.B2(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_37),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_28),
.B1(n_25),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_65),
.B1(n_33),
.B2(n_29),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_72),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_68),
.Y(n_96)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_70),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_29),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_77),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_76),
.A2(n_41),
.B1(n_39),
.B2(n_45),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_31),
.B1(n_33),
.B2(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_51),
.B1(n_48),
.B2(n_67),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_39),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_80),
.B(n_86),
.C(n_92),
.Y(n_126)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_100),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_25),
.B(n_21),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_44),
.B1(n_41),
.B2(n_39),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_61),
.B1(n_50),
.B2(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NAND2xp67_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_17),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_63),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_50),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_43),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_112),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_62),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_79),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_108),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_124),
.B1(n_125),
.B2(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_83),
.B1(n_98),
.B2(n_88),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_119),
.Y(n_143)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_116),
.Y(n_156)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_56),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_122),
.B(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_64),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_92),
.B1(n_95),
.B2(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_77),
.C(n_93),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_139),
.C(n_155),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_154),
.B1(n_111),
.B2(n_152),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_89),
.B1(n_76),
.B2(n_91),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_141),
.B1(n_107),
.B2(n_109),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_151),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_110),
.C(n_122),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_93),
.B1(n_79),
.B2(n_87),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_86),
.B(n_88),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_147),
.B(n_105),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_93),
.B(n_83),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_41),
.B1(n_39),
.B2(n_94),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_41),
.B1(n_94),
.B2(n_68),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_123),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_75),
.B1(n_27),
.B2(n_18),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_75),
.C(n_73),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_126),
.B(n_101),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_160),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_179),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_180),
.B1(n_181),
.B2(n_18),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_118),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_108),
.B(n_106),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_137),
.Y(n_172)
);

BUFx4f_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_153),
.B(n_155),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_183),
.B1(n_148),
.B2(n_142),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_134),
.B1(n_132),
.B2(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_127),
.B1(n_114),
.B2(n_128),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_127),
.B(n_27),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_147),
.C(n_145),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_127),
.B1(n_116),
.B2(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_176),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_203),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_132),
.B1(n_151),
.B2(n_99),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_73),
.B1(n_40),
.B2(n_137),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_199),
.B1(n_204),
.B2(n_159),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_73),
.B1(n_40),
.B2(n_19),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_24),
.B1(n_19),
.B2(n_21),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_202),
.B(n_184),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_40),
.B1(n_19),
.B2(n_24),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_176),
.C(n_182),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_229),
.C(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_190),
.B(n_168),
.CI(n_157),
.CON(n_220),
.SN(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_235),
.B1(n_210),
.B2(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_163),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_189),
.B1(n_3),
.B2(n_4),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_170),
.C(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_24),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_34),
.B(n_24),
.C(n_23),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_232),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_202),
.A2(n_34),
.B(n_1),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_0),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_0),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_221),
.B1(n_215),
.B2(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_252),
.C(n_234),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_235),
.B1(n_222),
.B2(n_226),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_198),
.C(n_189),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_249),
.C(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_189),
.C(n_205),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_202),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_256),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_228),
.B(n_202),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_237),
.B1(n_215),
.B2(n_212),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_11),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_1),
.C(n_4),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_272),
.Y(n_290)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_276),
.C(n_256),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_227),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_219),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_270),
.B(n_244),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_213),
.B(n_223),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_278),
.B(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_219),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_243),
.A2(n_220),
.B1(n_232),
.B2(n_214),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_216),
.C(n_225),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_220),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_281),
.B(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_238),
.C(n_250),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_245),
.C(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_271),
.C(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_252),
.C(n_241),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_293),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_241),
.B(n_242),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_225),
.B(n_233),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_264),
.B(n_254),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_254),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_274),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_251),
.B(n_270),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_308),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_274),
.B1(n_236),
.B2(n_6),
.Y(n_300)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_284),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_303)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_295),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_11),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_307),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_12),
.Y(n_307)
);

OAI21x1_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_12),
.B(n_15),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_290),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_313),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_289),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_294),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_281),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_315),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_13),
.C(n_14),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_10),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_306),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_299),
.B(n_301),
.Y(n_321)
);

AOI321xp33_ASAP7_75t_SL g333 ( 
.A1(n_321),
.A2(n_13),
.A3(n_16),
.B1(n_6),
.B2(n_4),
.C(n_5),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_317),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_302),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_328),
.B(n_13),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_320),
.A2(n_298),
.B1(n_10),
.B2(n_8),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.C(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_16),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_312),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_327),
.B(n_331),
.Y(n_336)
);

OAI321xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.A3(n_321),
.B1(n_334),
.B2(n_332),
.C(n_16),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_5),
.Y(n_339)
);


endmodule