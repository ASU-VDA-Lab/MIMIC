module real_jpeg_25990_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_295;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_51),
.B1(n_67),
.B2(n_68),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_67),
.B1(n_68),
.B2(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_81),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_4),
.A2(n_54),
.B1(n_67),
.B2(n_68),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_4),
.A2(n_33),
.B1(n_54),
.B2(n_123),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_42),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_8),
.A2(n_39),
.B1(n_67),
.B2(n_68),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_110),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_110),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_110),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_10),
.B(n_43),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_10),
.B(n_67),
.C(n_75),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_107),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_70),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_12),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_159),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_159),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_12),
.A2(n_67),
.B1(n_68),
.B2(n_159),
.Y(n_229)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_15),
.Y(n_222)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_15),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_138),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_19),
.B(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_92),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_20),
.B(n_83),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_57),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_44),
.C(n_82),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_40),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_24),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_24),
.A2(n_26),
.B1(n_157),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_25),
.A2(n_38),
.B1(n_43),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_25),
.A2(n_43),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_27),
.A2(n_30),
.B(n_154),
.C(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_28),
.B(n_29),
.C(n_123),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_29),
.A2(n_30),
.B1(n_46),
.B2(n_49),
.Y(n_56)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g247 ( 
.A(n_30),
.B(n_155),
.CON(n_247),
.SN(n_247)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_30),
.B(n_47),
.C(n_49),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_35),
.Y(n_162)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_36),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_41),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_43),
.B(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_50),
.B(n_52),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_45),
.A2(n_105),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_46),
.A2(n_48),
.B(n_247),
.C(n_248),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_48),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_48),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_50),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_53),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_107),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_55),
.A2(n_107),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_55),
.A2(n_107),
.B1(n_187),
.B2(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_72),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_58),
.A2(n_59),
.B1(n_72),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_69),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_61),
.A2(n_70),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_62),
.A2(n_69),
.B(n_174),
.Y(n_192)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_71),
.Y(n_97)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_67),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_70),
.B(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_66),
.A2(n_97),
.B(n_218),
.Y(n_249)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_68),
.B1(n_75),
.B2(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_68),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_70),
.A2(n_95),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_70),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_70),
.A2(n_175),
.B1(n_220),
.B2(n_229),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_72),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_80),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_73),
.A2(n_88),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_73),
.A2(n_78),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_73),
.A2(n_78),
.B1(n_205),
.B2(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_73),
.A2(n_128),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_79),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_78),
.B(n_155),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_85),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_90),
.A2(n_100),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_92),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.C(n_108),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_93),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_94),
.B(n_98),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_101),
.A2(n_102),
.B1(n_108),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_104),
.B(n_107),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_105),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_108),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_109),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_135),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_125),
.B2(n_126),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_124),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_123),
.B(n_155),
.CON(n_154),
.SN(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_130),
.B(n_134),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_292),
.B(n_296),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_193),
.B(n_279),
.C(n_291),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_179),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_141),
.B(n_179),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_163),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_143),
.B(n_146),
.C(n_163),
.Y(n_280)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_171),
.B2(n_178),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_166),
.B(n_168),
.C(n_178),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_176),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_184),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_183),
.B(n_184),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_191),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_185),
.B(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_264)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_278),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_273),
.B(n_277),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_259),
.B(n_272),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_243),
.B(n_258),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_215),
.B(n_242),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_206),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_212),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_226),
.B(n_241),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_224),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_223),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_237),
.B(n_240),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_257),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_257),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_253),
.C(n_256),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_268),
.C(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);


endmodule