module fake_jpeg_8549_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_19),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_21),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_18),
.B1(n_22),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_30),
.B1(n_22),
.B2(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_25),
.CON(n_55),
.SN(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_63),
.B1(n_30),
.B2(n_18),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_41),
.C(n_39),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_44),
.C(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_78),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_84),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_81),
.B1(n_83),
.B2(n_16),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_26),
.B(n_16),
.C(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_58),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_61),
.B1(n_56),
.B2(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_90),
.B1(n_72),
.B2(n_17),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_98),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_61),
.B1(n_59),
.B2(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_102),
.B1(n_76),
.B2(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_60),
.B1(n_23),
.B2(n_56),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_67),
.C(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_53),
.B1(n_16),
.B2(n_19),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_24),
.B1(n_54),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_27),
.B1(n_25),
.B2(n_15),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_27),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_122),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2x1p5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_66),
.Y(n_114)
);

XOR2x2_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_101),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_65),
.B(n_77),
.C(n_17),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_121),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_72),
.B1(n_65),
.B2(n_66),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_123),
.B1(n_125),
.B2(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_1),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_102),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_106),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_137),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_142),
.B1(n_126),
.B2(n_107),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_99),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_147),
.C(n_108),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_94),
.B(n_91),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_116),
.B(n_86),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_109),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_115),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_118),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_121),
.C(n_114),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_157),
.B1(n_135),
.B2(n_136),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_111),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_86),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_109),
.C(n_69),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_143),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_159),
.A2(n_142),
.B(n_140),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_132),
.B1(n_134),
.B2(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_177),
.B1(n_176),
.B2(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_176),
.B1(n_168),
.B2(n_171),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_69),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_160),
.B1(n_152),
.B2(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_170),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_186),
.B(n_188),
.C(n_189),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_167),
.B1(n_1),
.B2(n_6),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_167),
.Y(n_188)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_185),
.B1(n_187),
.B2(n_190),
.C(n_188),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_191),
.A2(n_192),
.B1(n_7),
.B2(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_11),
.C(n_12),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_12),
.B(n_13),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_14),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);


endmodule