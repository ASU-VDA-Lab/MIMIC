module fake_jpeg_31106_n_180 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_31),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_1),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_1),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_53),
.B1(n_60),
.B2(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_58),
.B1(n_76),
.B2(n_29),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_72),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_73),
.Y(n_96)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_108),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_111),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_119),
.B(n_2),
.Y(n_125)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_52),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_65),
.B1(n_63),
.B2(n_66),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_76),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_74),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_60),
.B(n_68),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_33),
.B(n_46),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_121),
.Y(n_131)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_63),
.B1(n_62),
.B2(n_59),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_76),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_128),
.B1(n_132),
.B2(n_136),
.Y(n_143)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_131),
.B(n_124),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_35),
.C(n_45),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_122),
.C(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_11),
.B1(n_12),
.B2(n_20),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_22),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_44),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_40),
.B1(n_43),
.B2(n_130),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_150),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_125),
.CON(n_150),
.SN(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_156),
.B1(n_133),
.B2(n_143),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_158),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_150),
.B(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_164),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_146),
.B1(n_155),
.B2(n_147),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_146),
.B1(n_160),
.B2(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_167),
.C(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_155),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);

AOI21x1_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_172),
.B(n_166),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_157),
.Y(n_179)
);

NAND2x1_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_161),
.Y(n_180)
);


endmodule