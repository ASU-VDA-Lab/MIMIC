module real_jpeg_27971_n_17 (n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_34),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_0),
.A2(n_56),
.B1(n_98),
.B2(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_0),
.A2(n_56),
.B1(n_157),
.B2(n_163),
.Y(n_190)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_2),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_115),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_98),
.B1(n_99),
.B2(n_115),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_2),
.A2(n_115),
.B1(n_157),
.B2(n_163),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_3),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_5),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_34),
.B1(n_36),
.B2(n_197),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_5),
.A2(n_98),
.B1(n_99),
.B2(n_197),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_5),
.A2(n_157),
.B1(n_163),
.B2(n_197),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_45),
.B1(n_98),
.B2(n_99),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_45),
.B1(n_157),
.B2(n_163),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_8),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_216),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_8),
.A2(n_98),
.B1(n_99),
.B2(n_216),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_8),
.A2(n_157),
.B1(n_163),
.B2(n_216),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_9),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_9),
.A2(n_34),
.B1(n_36),
.B2(n_153),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_9),
.A2(n_98),
.B1(n_99),
.B2(n_153),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_9),
.A2(n_153),
.B1(n_157),
.B2(n_163),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_36),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_35),
.B(n_36),
.C(n_40),
.D(n_43),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_10),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_60),
.B(n_64),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_98),
.B(n_100),
.C(n_101),
.D(n_105),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_10),
.B(n_98),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_10),
.A2(n_99),
.B(n_133),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_10),
.A2(n_82),
.B1(n_157),
.B2(n_163),
.Y(n_164)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_11),
.A2(n_36),
.B(n_41),
.C(n_42),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_12),
.A2(n_34),
.B1(n_36),
.B2(n_136),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_12),
.A2(n_98),
.B1(n_99),
.B2(n_136),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_12),
.A2(n_136),
.B1(n_157),
.B2(n_163),
.Y(n_288)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_14),
.A2(n_34),
.B1(n_36),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_14),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_15),
.A2(n_34),
.B1(n_36),
.B2(n_63),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_15),
.A2(n_63),
.B1(n_98),
.B2(n_99),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_15),
.A2(n_63),
.B1(n_157),
.B2(n_163),
.Y(n_208)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_325),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_312),
.B(n_324),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_276),
.A3(n_305),
.B1(n_310),
.B2(n_311),
.C(n_333),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_226),
.A3(n_265),
.B1(n_270),
.B2(n_275),
.C(n_334),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_177),
.C(n_222),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_144),
.B(n_176),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_120),
.B(n_143),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_93),
.B(n_119),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_69),
.B(n_92),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_47),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_27),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_39),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_29),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_30),
.B(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_34),
.B(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_36),
.A2(n_99),
.A3(n_100),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_40),
.A2(n_42),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_40),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_40),
.A2(n_42),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_40),
.A2(n_42),
.B1(n_242),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_43),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_46),
.A2(n_57),
.B(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_46),
.A2(n_140),
.B1(n_175),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_46),
.A2(n_140),
.B1(n_199),
.B2(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_46),
.A2(n_140),
.B(n_251),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_59),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_54),
.C(n_59),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_51),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_51),
.A2(n_101),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_51),
.A2(n_101),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_51),
.A2(n_101),
.B1(n_254),
.B2(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_51),
.A2(n_101),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_55),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_68),
.B1(n_114),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_60),
.A2(n_68),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_60),
.A2(n_196),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_60),
.A2(n_77),
.B(n_215),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_74),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx5_ASAP7_75t_SL g214 ( 
.A(n_67),
.Y(n_214)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_82),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_79),
.B(n_91),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_77),
.B(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_85),
.B(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_90),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_82),
.B(n_130),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_82),
.A2(n_132),
.B(n_156),
.C(n_157),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_111),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_108),
.C(n_111),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_99),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_107),
.A2(n_126),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_107),
.A2(n_185),
.B1(n_211),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_107),
.A2(n_185),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_137),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_138),
.C(n_139),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_129),
.C(n_134),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_130),
.A2(n_189),
.B(n_191),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_130),
.A2(n_191),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_130),
.A2(n_233),
.B1(n_261),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_130),
.A2(n_233),
.B1(n_288),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_131),
.A2(n_161),
.B1(n_190),
.B2(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_131),
.A2(n_161),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_131),
.A2(n_161),
.B1(n_320),
.B2(n_329),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_133),
.B1(n_157),
.B2(n_163),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_135),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_146),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_159),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_148),
.B(n_149),
.C(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_154),
.B1(n_155),
.B2(n_158),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_157),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_170),
.C(n_173),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B(n_165),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_166),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_178),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_201),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_179),
.B(n_201),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_193),
.C(n_200),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_183),
.C(n_192),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_192),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B(n_187),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_200),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_198),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_212),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_203),
.B(n_212),
.C(n_221),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_217),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_224),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_246),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_246),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.C(n_245),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_238),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_237),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_235),
.C(n_237),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_244),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_244),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_244),
.A2(n_259),
.B(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_264),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_256),
.B1(n_257),
.B2(n_263),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_252),
.B(n_255),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_252),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_255),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_255),
.A2(n_278),
.B1(n_279),
.B2(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_256),
.B(n_263),
.C(n_264),
.Y(n_306)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_268),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_293),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_290),
.C(n_291),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_287),
.B2(n_289),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_282),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_286),
.C(n_287),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_283),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_284),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_286),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_297),
.C(n_301),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_289),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_296),
.C(n_304),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_292),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_304),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_298),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_318),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_316),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_322),
.C(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_330),
.Y(n_331)
);


endmodule