module fake_jpeg_14020_n_390 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_59),
.Y(n_104)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_58),
.Y(n_114)
);

CKINVDCx11_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_62),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_63),
.B(n_7),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_72),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_78),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_2),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

BUFx24_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_17),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_96),
.Y(n_106)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_92),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_33),
.Y(n_91)
);

CKINVDCx12_ASAP7_75t_R g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_7),
.Y(n_129)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_98),
.Y(n_155)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_99),
.B(n_102),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_86),
.Y(n_107)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_103),
.B(n_10),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_108),
.B(n_125),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_48),
.B1(n_52),
.B2(n_41),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_109),
.A2(n_119),
.B1(n_135),
.B2(n_124),
.Y(n_209)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_41),
.B1(n_52),
.B2(n_29),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_44),
.B1(n_51),
.B2(n_47),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_137),
.B1(n_153),
.B2(n_83),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_20),
.B1(n_19),
.B2(n_40),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_124),
.A2(n_135),
.B1(n_156),
.B2(n_162),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_53),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_129),
.B(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_46),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_19),
.B1(n_40),
.B2(n_44),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_51),
.B1(n_47),
.B2(n_44),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_35),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_150),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_35),
.C(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_36),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_75),
.A2(n_51),
.B1(n_47),
.B2(n_43),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_157),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_102),
.A2(n_43),
.B1(n_39),
.B2(n_50),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_92),
.B(n_43),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_68),
.B(n_49),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_163),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_57),
.A2(n_39),
.B1(n_49),
.B2(n_36),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_57),
.B(n_12),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_14),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_170),
.B(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_155),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_198),
.Y(n_229)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_175),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_76),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_184),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_93),
.B1(n_87),
.B2(n_82),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_179),
.A2(n_181),
.B1(n_195),
.B2(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_69),
.B1(n_60),
.B2(n_101),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_156),
.B1(n_162),
.B2(n_130),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g258 ( 
.A(n_183),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_14),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_106),
.B(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_16),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_191),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_117),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_193),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_104),
.B(n_16),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_119),
.B(n_18),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_200),
.C(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_18),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_22),
.B1(n_128),
.B2(n_142),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_22),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_161),
.B(n_22),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_138),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_204),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_119),
.A2(n_109),
.B(n_127),
.C(n_138),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_109),
.A2(n_127),
.B(n_136),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_207),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_149),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_114),
.B(n_22),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_205),
.B(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_161),
.B(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_210),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_121),
.B1(n_158),
.B2(n_115),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_105),
.B(n_122),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_128),
.B(n_147),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_148),
.A2(n_122),
.B1(n_147),
.B2(n_132),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_115),
.B(n_110),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_194),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_220),
.A2(n_245),
.B1(n_252),
.B2(n_256),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_221),
.A2(n_222),
.B1(n_246),
.B2(n_250),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_158),
.B1(n_113),
.B2(n_132),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_113),
.B(n_110),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_228),
.A2(n_244),
.B(n_198),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_180),
.A2(n_110),
.B(n_199),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_237),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_177),
.C(n_190),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_241),
.C(n_231),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_175),
.A2(n_200),
.B(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_172),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_257),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_186),
.B(n_182),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_188),
.A2(n_164),
.B(n_202),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_181),
.A2(n_176),
.B1(n_167),
.B2(n_166),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_171),
.A2(n_165),
.B1(n_169),
.B2(n_217),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_203),
.B1(n_207),
.B2(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_178),
.A2(n_174),
.B1(n_183),
.B2(n_187),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_178),
.A2(n_208),
.B1(n_202),
.B2(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_208),
.A2(n_192),
.B1(n_188),
.B2(n_180),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_269),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_228),
.B(n_251),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_284),
.B(n_286),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_204),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_283),
.C(n_291),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_245),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_SL g298 ( 
.A(n_271),
.B(n_274),
.C(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_272),
.B(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_225),
.B(n_239),
.C(n_230),
.D(n_235),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_224),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_229),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_287),
.Y(n_306)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_249),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_285),
.Y(n_293)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_251),
.C(n_241),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_251),
.B1(n_233),
.B2(n_221),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_252),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_244),
.A2(n_242),
.B(n_229),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_229),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_289),
.Y(n_312)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_222),
.B(n_236),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_250),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_220),
.B(n_234),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_302),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_240),
.B(n_219),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_298),
.B(n_313),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_270),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_243),
.B1(n_248),
.B2(n_258),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_314),
.B1(n_289),
.B2(n_265),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_301),
.B(n_316),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_240),
.C(n_243),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_253),
.B(n_254),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_264),
.A2(n_254),
.B1(n_258),
.B2(n_290),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_258),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_264),
.B1(n_285),
.B2(n_260),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_330),
.B1(n_314),
.B2(n_310),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_335),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_305),
.A2(n_279),
.B(n_268),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_322),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_292),
.B(n_296),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_325),
.B(n_311),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_323),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_261),
.B(n_286),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_272),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_283),
.C(n_278),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_277),
.C(n_280),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_277),
.C(n_271),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_331),
.C(n_335),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_275),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_274),
.C(n_275),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_336),
.A2(n_299),
.B1(n_307),
.B2(n_311),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_334),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

XNOR2x2_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_329),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_284),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_310),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_348),
.A2(n_332),
.B(n_339),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_295),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_340),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_299),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_323),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_327),
.C(n_333),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_353),
.C(n_345),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_321),
.C(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_355),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_359),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_357),
.A2(n_361),
.B1(n_348),
.B2(n_339),
.Y(n_367)
);

XOR2x2_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_325),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_362),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_360),
.B(n_338),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_346),
.A2(n_307),
.B1(n_298),
.B2(n_300),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_366),
.C(n_359),
.Y(n_372)
);

OA21x2_ASAP7_75t_SL g366 ( 
.A1(n_354),
.A2(n_343),
.B(n_338),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_361),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_352),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_347),
.C(n_349),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_371),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_347),
.B1(n_337),
.B2(n_303),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_SL g380 ( 
.A(n_372),
.B(n_377),
.Y(n_380)
);

OAI221xp5_ASAP7_75t_L g382 ( 
.A1(n_373),
.A2(n_363),
.B1(n_369),
.B2(n_365),
.C(n_315),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_371),
.A2(n_353),
.B(n_369),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_376),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_315),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_337),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_383),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_375),
.B(n_373),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_370),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_384),
.A2(n_386),
.B(n_377),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_380),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_387),
.B(n_388),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_385),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g390 ( 
.A(n_389),
.B(n_284),
.CI(n_303),
.CON(n_390),
.SN(n_390)
);


endmodule