module fake_jpeg_30248_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g126 ( 
.A(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_62),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_0),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_48),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_64),
.B(n_89),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_35),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_77),
.B(n_46),
.Y(n_163)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_81),
.B(n_82),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_84),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_1),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_39),
.B1(n_45),
.B2(n_29),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_35),
.B(n_3),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_102),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_36),
.B(n_4),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_47),
.Y(n_160)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_111),
.B(n_135),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_54),
.A2(n_50),
.B1(n_34),
.B2(n_28),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_112),
.A2(n_136),
.B1(n_66),
.B2(n_59),
.Y(n_215)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_115),
.Y(n_183)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_77),
.B(n_21),
.CON(n_129),
.SN(n_129)
);

OR2x4_ASAP7_75t_L g205 ( 
.A(n_129),
.B(n_44),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_102),
.B1(n_28),
.B2(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_131),
.A2(n_133),
.B1(n_44),
.B2(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_62),
.B(n_52),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_56),
.A2(n_43),
.B1(n_28),
.B2(n_32),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_45),
.B(n_52),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_84),
.B(n_44),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_148),
.B(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_58),
.B(n_49),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_49),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_155),
.B(n_162),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_160),
.B(n_163),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_29),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_60),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_179),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_172),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_39),
.B1(n_47),
.B2(n_76),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_177),
.B(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_120),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_142),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_181),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_95),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_182),
.B(n_190),
.Y(n_245)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_78),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_186),
.B(n_206),
.Y(n_239)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_92),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_115),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_129),
.A2(n_104),
.B1(n_72),
.B2(n_105),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_192),
.A2(n_214),
.B1(n_86),
.B2(n_94),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_194),
.A2(n_96),
.B(n_25),
.Y(n_261)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_201),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_23),
.B1(n_32),
.B2(n_100),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_199),
.A2(n_215),
.B1(n_222),
.B2(n_156),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_21),
.B(n_44),
.C(n_67),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_134),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_71),
.Y(n_202)
);

OR2x6_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_158),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_74),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_109),
.B(n_79),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_210),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_126),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_211),
.B(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_150),
.B(n_69),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_110),
.Y(n_216)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_218),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_144),
.B(n_99),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_53),
.C(n_25),
.Y(n_276)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_224),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_137),
.A2(n_23),
.B1(n_106),
.B2(n_98),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_108),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_112),
.B(n_158),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_228),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_227),
.A2(n_146),
.B1(n_158),
.B2(n_139),
.Y(n_234)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_131),
.B1(n_150),
.B2(n_117),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_235),
.A2(n_237),
.B1(n_249),
.B2(n_259),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_194),
.A2(n_176),
.B1(n_200),
.B2(n_205),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_236),
.B(n_248),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_178),
.A2(n_117),
.B1(n_57),
.B2(n_65),
.Y(n_237)
);

AO22x2_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_137),
.B1(n_151),
.B2(n_75),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_260),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_151),
.B1(n_165),
.B2(n_128),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_263),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_203),
.A2(n_146),
.B1(n_145),
.B2(n_166),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_257),
.A2(n_227),
.B1(n_183),
.B2(n_187),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_202),
.A2(n_165),
.B1(n_128),
.B2(n_130),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_138),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_220),
.B(n_206),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_206),
.A2(n_138),
.B1(n_141),
.B2(n_140),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_271),
.B1(n_235),
.B2(n_239),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_141),
.B1(n_140),
.B2(n_130),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_209),
.B(n_145),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_217),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_248),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_254),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_223),
.B(n_204),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_279),
.B(n_299),
.C(n_303),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_281),
.A2(n_282),
.B(n_244),
.Y(n_338)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_207),
.B(n_212),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_218),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_283),
.B(n_290),
.Y(n_339)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_183),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_295),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_252),
.A2(n_181),
.B1(n_175),
.B2(n_173),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_289),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_250),
.B(n_218),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_247),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_293),
.Y(n_319)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_298),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_233),
.A2(n_196),
.A3(n_195),
.B1(n_197),
.B2(n_183),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_297),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_183),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_233),
.B(n_20),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_232),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_302),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_230),
.B(n_184),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_241),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_267),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_314),
.Y(n_337)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_213),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_308),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_174),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_239),
.B(n_220),
.C(n_171),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_276),
.C(n_260),
.Y(n_326)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_315),
.Y(n_353)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_238),
.A2(n_198),
.B(n_53),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_281),
.B(n_263),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_20),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_292),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_286),
.B1(n_312),
.B2(n_316),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_243),
.B(n_236),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_320),
.A2(n_328),
.B(n_296),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_286),
.A2(n_253),
.B1(n_242),
.B2(n_244),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_343),
.B1(n_294),
.B2(n_291),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_288),
.A2(n_236),
.B(n_246),
.C(n_243),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g376 ( 
.A1(n_323),
.A2(n_325),
.B(n_332),
.C(n_345),
.Y(n_376)
);

NAND2x1p5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_246),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_352),
.C(n_354),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_350),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_300),
.A2(n_272),
.B(n_265),
.Y(n_328)
);

AO21x2_ASAP7_75t_L g332 ( 
.A1(n_297),
.A2(n_295),
.B(n_305),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_305),
.A2(n_259),
.B1(n_237),
.B2(n_246),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_334),
.A2(n_346),
.B1(n_277),
.B2(n_285),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_347),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_284),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_246),
.B1(n_264),
.B2(n_255),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_278),
.A2(n_252),
.B(n_251),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_344),
.A2(n_231),
.B(n_314),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_284),
.A2(n_282),
.B(n_305),
.C(n_312),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_299),
.A2(n_221),
.B1(n_266),
.B2(n_251),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_315),
.A2(n_264),
.B1(n_255),
.B2(n_266),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_303),
.A2(n_266),
.B1(n_273),
.B2(n_262),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_5),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_273),
.C(n_262),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_193),
.C(n_189),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_355),
.B(n_6),
.Y(n_389)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_357),
.A2(n_367),
.B(n_381),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_361),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_359),
.Y(n_398)
);

INVx11_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_337),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_298),
.C(n_293),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_372),
.C(n_379),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_377),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_366),
.A2(n_378),
.B1(n_343),
.B2(n_365),
.Y(n_395)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_340),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_371),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_301),
.C(n_306),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_319),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_374),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_337),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_375),
.Y(n_410)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_334),
.A2(n_277),
.B1(n_172),
.B2(n_188),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_382),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_309),
.C(n_313),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_335),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_348),
.B(n_349),
.C(n_333),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_320),
.A2(n_310),
.B(n_287),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_344),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_231),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_287),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_327),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_328),
.A2(n_5),
.B(n_6),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_389),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_388),
.A2(n_346),
.B1(n_341),
.B2(n_336),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_401),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_392),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_362),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_394),
.B(n_402),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_395),
.A2(n_377),
.B1(n_332),
.B2(n_386),
.Y(n_428)
);

AOI21xp33_ASAP7_75t_SL g397 ( 
.A1(n_385),
.A2(n_329),
.B(n_324),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_397),
.B(n_404),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_358),
.B(n_355),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_370),
.A2(n_321),
.B1(n_345),
.B2(n_332),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_405),
.A2(n_376),
.B1(n_375),
.B2(n_374),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_363),
.B(n_332),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_381),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_354),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_367),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_388),
.A2(n_348),
.B1(n_330),
.B2(n_345),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_412),
.A2(n_383),
.B1(n_357),
.B2(n_361),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_420),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_345),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_418),
.C(n_379),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_345),
.C(n_322),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g420 ( 
.A(n_370),
.B(n_325),
.CI(n_332),
.CON(n_420),
.SN(n_420)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_405),
.A2(n_357),
.B1(n_366),
.B2(n_356),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_421),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_422),
.A2(n_428),
.B1(n_443),
.B2(n_445),
.Y(n_450)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_402),
.A2(n_376),
.B1(n_368),
.B2(n_382),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_435),
.Y(n_448)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_427),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_437),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_390),
.Y(n_434)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_387),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_439),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_380),
.B1(n_323),
.B2(n_359),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_376),
.B1(n_325),
.B2(n_323),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_442),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_416),
.A2(n_323),
.B1(n_350),
.B2(n_369),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_410),
.A2(n_323),
.B1(n_349),
.B2(n_360),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_444),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_409),
.A2(n_399),
.B1(n_396),
.B2(n_406),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_7),
.C(n_8),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_392),
.C(n_419),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_447),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_451),
.B(n_463),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_430),
.A2(n_407),
.B(n_392),
.Y(n_452)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_414),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_437),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_394),
.C(n_417),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_458),
.C(n_446),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_418),
.C(n_391),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_428),
.A2(n_406),
.B1(n_413),
.B2(n_409),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_459),
.A2(n_467),
.B1(n_456),
.B2(n_461),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_438),
.B(n_419),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_413),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_442),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_427),
.A2(n_420),
.B1(n_415),
.B2(n_398),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_456),
.A2(n_430),
.B(n_431),
.C(n_434),
.Y(n_471)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_471),
.Y(n_491)
);

BUFx12_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_481),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_425),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_480),
.Y(n_492)
);

XNOR2x1_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_426),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_474),
.B(n_479),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_460),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_485),
.C(n_486),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_453),
.A2(n_421),
.B1(n_423),
.B2(n_443),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_435),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_454),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_467),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_482),
.A2(n_452),
.B1(n_465),
.B2(n_450),
.Y(n_488)
);

AO221x1_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_403),
.B1(n_441),
.B2(n_436),
.C(n_408),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_484),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_440),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_482),
.A2(n_450),
.B1(n_454),
.B2(n_461),
.Y(n_487)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_487),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_490),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_478),
.A2(n_459),
.B1(n_448),
.B2(n_449),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_455),
.C(n_462),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_499),
.C(n_474),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_480),
.A2(n_448),
.B1(n_464),
.B2(n_447),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_16),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_462),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_496),
.B(n_502),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_420),
.C(n_398),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_408),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_492),
.A2(n_478),
.B(n_471),
.Y(n_503)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_503),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_513),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_500),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_506),
.B(n_511),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_492),
.A2(n_493),
.B(n_494),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_508),
.B(n_509),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_493),
.A2(n_472),
.B(n_484),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_479),
.C(n_472),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_7),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_512),
.A2(n_514),
.B(n_9),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_9),
.C(n_10),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_491),
.A2(n_9),
.B(n_11),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_515),
.A2(n_497),
.B1(n_501),
.B2(n_487),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_517),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_518),
.B(n_11),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_499),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_522),
.C(n_524),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_504),
.A2(n_488),
.B1(n_490),
.B2(n_501),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_9),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_510),
.C(n_513),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_528),
.Y(n_532)
);

MAJx2_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_11),
.C(n_12),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_530),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_521),
.C(n_523),
.Y(n_531)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_523),
.A3(n_527),
.B1(n_519),
.B2(n_524),
.C1(n_13),
.C2(n_16),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_532),
.C(n_14),
.Y(n_535)
);

NAND2x1_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_534),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_536),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_13),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_16),
.B(n_492),
.Y(n_539)
);


endmodule