module real_jpeg_12447_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_3),
.A2(n_37),
.B1(n_39),
.B2(n_68),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_5),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_117),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_37),
.B1(n_39),
.B2(n_79),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_26),
.C(n_42),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g138 ( 
.A(n_5),
.B(n_63),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_100),
.B(n_144),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_5),
.A2(n_59),
.B(n_62),
.C(n_171),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_5),
.A2(n_60),
.B1(n_62),
.B2(n_79),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_37),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_46),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_65),
.B1(n_73),
.B2(n_74),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_37),
.B1(n_39),
.B2(n_65),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_65),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_53),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_53),
.B1(n_60),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_53),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_19),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_84),
.B2(n_85),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_23)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_24),
.A2(n_29),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_145),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_25),
.B(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_29),
.B(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_37),
.B(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_39),
.A2(n_58),
.B(n_79),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_40),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_40),
.A2(n_47),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_50),
.B(n_51),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_44),
.A2(n_51),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_44),
.B(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_47),
.B(n_52),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_69),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_49),
.B(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_67),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_55),
.A2(n_89),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_90),
.Y(n_114)
);

NOR2x1_ASAP7_75t_R g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_62),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_60),
.B(n_76),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_74),
.A3(n_77),
.B1(n_81),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_66),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_70),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_83)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_79),
.B(n_80),
.C(n_82),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_79),
.B(n_102),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_97),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_96),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_103),
.B1(n_104),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_150),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_102),
.A2(n_119),
.B(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_107),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_112),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.C(n_118),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_113),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_197),
.B(n_201),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_182),
.B(n_196),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_166),
.B(n_181),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_146),
.B(n_165),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B(n_132),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_131),
.A2(n_132),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_154),
.B(n_164),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_152),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_159),
.B(n_163),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_168),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_176),
.C(n_180),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_192),
.C(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);


endmodule