module real_aes_9048_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g515 ( .A(n_1), .Y(n_515) );
INVx1_ASAP7_75t_L g196 ( .A(n_2), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_3), .A2(n_38), .B1(n_158), .B2(n_457), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_4), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g137 ( .A1(n_5), .A2(n_138), .B(n_145), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_6), .B(n_131), .Y(n_506) );
AND2x6_ASAP7_75t_L g143 ( .A(n_7), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_8), .A2(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_9), .B(n_39), .Y(n_114) );
INVx1_ASAP7_75t_L g155 ( .A(n_10), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_11), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_13), .B(n_168), .Y(n_452) );
INVx1_ASAP7_75t_L g243 ( .A(n_14), .Y(n_243) );
INVx1_ASAP7_75t_L g510 ( .A(n_15), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_16), .B(n_132), .Y(n_491) );
AO32x2_ASAP7_75t_L g472 ( .A1(n_17), .A2(n_131), .A3(n_165), .B1(n_473), .B2(n_477), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_18), .B(n_158), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_19), .B(n_184), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_20), .B(n_132), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_21), .A2(n_50), .B1(n_158), .B2(n_457), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_22), .B(n_138), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_23), .A2(n_76), .B1(n_158), .B2(n_168), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_24), .B(n_158), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_25), .B(n_129), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_26), .A2(n_241), .B(n_242), .C(n_244), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_27), .A2(n_74), .B1(n_726), .B2(n_727), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_27), .Y(n_727) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_29), .B(n_161), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_30), .B(n_153), .Y(n_198) );
INVx1_ASAP7_75t_L g174 ( .A(n_31), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_32), .B(n_161), .Y(n_470) );
INVx2_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_34), .B(n_158), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_35), .B(n_161), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_36), .A2(n_62), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_36), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_37), .A2(n_143), .B(n_148), .C(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g172 ( .A(n_40), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_41), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_42), .B(n_153), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_43), .B(n_158), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_44), .A2(n_87), .B1(n_215), .B2(n_457), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_45), .B(n_158), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_46), .B(n_158), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_47), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_48), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_49), .B(n_138), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_51), .A2(n_60), .B1(n_158), .B2(n_168), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_52), .A2(n_148), .B1(n_168), .B2(n_170), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_53), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_54), .B(n_158), .Y(n_451) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_55), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_56), .B(n_158), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_57), .A2(n_152), .B(n_154), .C(n_157), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_58), .Y(n_261) );
INVx1_ASAP7_75t_L g146 ( .A(n_59), .Y(n_146) );
INVx1_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_62), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_63), .B(n_158), .Y(n_516) );
INVx1_ASAP7_75t_L g135 ( .A(n_64), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_65), .Y(n_738) );
AO32x2_ASAP7_75t_L g482 ( .A1(n_66), .A2(n_131), .A3(n_223), .B1(n_477), .B2(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g527 ( .A(n_67), .Y(n_527) );
INVx1_ASAP7_75t_L g465 ( .A(n_68), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_SL g183 ( .A1(n_69), .A2(n_157), .B(n_184), .C(n_185), .Y(n_183) );
INVxp67_ASAP7_75t_L g186 ( .A(n_70), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_71), .B(n_168), .Y(n_466) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_73), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_74), .Y(n_726) );
INVx1_ASAP7_75t_L g254 ( .A(n_75), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_77), .A2(n_102), .B1(n_115), .B2(n_755), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_78), .A2(n_143), .B(n_148), .C(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_79), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_80), .B(n_168), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_81), .B(n_197), .Y(n_211) );
INVx2_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_83), .B(n_184), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_84), .B(n_168), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_85), .A2(n_143), .B(n_148), .C(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
OR2x2_ASAP7_75t_L g121 ( .A(n_86), .B(n_112), .Y(n_121) );
OR2x2_ASAP7_75t_L g748 ( .A(n_86), .B(n_111), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_88), .A2(n_100), .B1(n_168), .B2(n_169), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_89), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_90), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_91), .A2(n_143), .B(n_148), .C(n_226), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_92), .Y(n_233) );
INVx1_ASAP7_75t_L g182 ( .A(n_93), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_94), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_95), .B(n_197), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_96), .B(n_168), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_97), .B(n_131), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_98), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_99), .A2(n_138), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g756 ( .A(n_105), .Y(n_756) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g734 ( .A(n_109), .Y(n_734) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g440 ( .A(n_110), .B(n_112), .Y(n_440) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AO221x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_736), .B1(n_739), .B2(n_749), .C(n_751), .Y(n_115) );
OAI222xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_724), .B1(n_725), .B2(n_728), .C1(n_732), .C2(n_735), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B1(n_439), .B2(n_441), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g729 ( .A(n_121), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_122), .A2(n_730), .B1(n_742), .B2(n_743), .Y(n_741) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g730 ( .A(n_123), .Y(n_730) );
AND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_361), .C(n_406), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_284), .C(n_325), .D(n_342), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_188), .B(n_204), .C(n_246), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_162), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_127), .B(n_189), .Y(n_188) );
NOR4xp25_ASAP7_75t_L g308 ( .A(n_127), .B(n_302), .C(n_309), .D(n_315), .Y(n_308) );
AND2x2_ASAP7_75t_L g381 ( .A(n_127), .B(n_270), .Y(n_381) );
AND2x2_ASAP7_75t_L g400 ( .A(n_127), .B(n_346), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_127), .B(n_395), .Y(n_409) );
AND2x2_ASAP7_75t_L g422 ( .A(n_127), .B(n_203), .Y(n_422) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_SL g267 ( .A(n_128), .Y(n_267) );
AND2x2_ASAP7_75t_L g274 ( .A(n_128), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g324 ( .A(n_128), .B(n_163), .Y(n_324) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_128), .B(n_270), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_128), .B(n_163), .Y(n_339) );
AND2x2_ASAP7_75t_L g348 ( .A(n_128), .B(n_273), .Y(n_348) );
BUFx2_ASAP7_75t_L g371 ( .A(n_128), .Y(n_371) );
AND2x2_ASAP7_75t_L g375 ( .A(n_128), .B(n_179), .Y(n_375) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_137), .B(n_160), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_SL g217 ( .A(n_130), .B(n_218), .Y(n_217) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_130), .B(n_477), .C(n_493), .Y(n_492) );
AO21x1_ASAP7_75t_L g530 ( .A1(n_130), .A2(n_493), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_131), .A2(n_180), .B(n_187), .Y(n_179) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_131), .A2(n_498), .B(n_506), .Y(n_497) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_133), .B(n_134), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx2_ASAP7_75t_L g237 ( .A(n_138), .Y(n_237) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_139), .B(n_143), .Y(n_176) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g505 ( .A(n_140), .Y(n_505) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
INVx1_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx1_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx4_ASAP7_75t_SL g159 ( .A(n_143), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_143), .A2(n_450), .B(n_454), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_143), .A2(n_464), .B(n_467), .Y(n_463) );
BUFx3_ASAP7_75t_L g477 ( .A(n_143), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_143), .A2(n_499), .B(n_502), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_143), .A2(n_509), .B(n_513), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_151), .C(n_159), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_147), .A2(n_159), .B(n_182), .C(n_183), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_147), .A2(n_159), .B(n_239), .C(n_240), .Y(n_238) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx3_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g457 ( .A(n_149), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_152), .A2(n_455), .B(n_456), .Y(n_454) );
O2A1O1Ixp5_ASAP7_75t_L g526 ( .A1(n_152), .A2(n_514), .B(n_527), .C(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g229 ( .A(n_153), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_153), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_153), .A2(n_156), .B1(n_484), .B2(n_485), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_153), .A2(n_475), .B1(n_494), .B2(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_156), .B(n_186), .Y(n_185) );
INVx5_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_SL g464 ( .A1(n_157), .A2(n_197), .B(n_465), .C(n_466), .Y(n_464) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_167), .B1(n_175), .B2(n_176), .Y(n_166) );
INVx1_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_161), .A2(n_236), .B(n_245), .Y(n_235) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_161), .A2(n_449), .B(n_458), .Y(n_448) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_161), .A2(n_463), .B(n_470), .Y(n_462) );
OR2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_179), .Y(n_162) );
AND2x2_ASAP7_75t_L g203 ( .A(n_163), .B(n_179), .Y(n_203) );
BUFx2_ASAP7_75t_L g277 ( .A(n_163), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_163), .A2(n_310), .B1(n_312), .B2(n_313), .Y(n_309) );
OR2x2_ASAP7_75t_L g331 ( .A(n_163), .B(n_191), .Y(n_331) );
AND2x2_ASAP7_75t_L g395 ( .A(n_163), .B(n_273), .Y(n_395) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g263 ( .A(n_164), .B(n_191), .Y(n_263) );
AND2x2_ASAP7_75t_L g270 ( .A(n_164), .B(n_179), .Y(n_270) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_164), .Y(n_312) );
OR2x2_ASAP7_75t_L g347 ( .A(n_164), .B(n_190), .Y(n_347) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_177), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_165), .B(n_178), .Y(n_177) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_165), .A2(n_192), .B(n_200), .Y(n_191) );
INVx2_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
INVx2_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_170) );
INVx2_ASAP7_75t_L g173 ( .A(n_171), .Y(n_173) );
INVx4_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_176), .A2(n_193), .B(n_194), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_176), .A2(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
INVx3_ASAP7_75t_L g275 ( .A(n_179), .Y(n_275) );
BUFx2_ASAP7_75t_L g299 ( .A(n_179), .Y(n_299) );
AND2x2_ASAP7_75t_L g332 ( .A(n_179), .B(n_267), .Y(n_332) );
INVx1_ASAP7_75t_L g453 ( .A(n_184), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_188), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_417) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_203), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_190), .B(n_275), .Y(n_279) );
INVx1_ASAP7_75t_L g307 ( .A(n_190), .Y(n_307) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g273 ( .A(n_191), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
INVx2_ASAP7_75t_L g475 ( .A(n_197), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_197), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_197), .A2(n_524), .B(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_199), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_202), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_202), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
NAND2x1_ASAP7_75t_SL g204 ( .A(n_205), .B(n_219), .Y(n_204) );
AND2x2_ASAP7_75t_L g283 ( .A(n_205), .B(n_234), .Y(n_283) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_205), .Y(n_357) );
AND2x2_ASAP7_75t_L g384 ( .A(n_205), .B(n_304), .Y(n_384) );
AND2x2_ASAP7_75t_L g392 ( .A(n_205), .B(n_354), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_205), .B(n_249), .Y(n_419) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g250 ( .A(n_206), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g268 ( .A(n_206), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
INVx1_ASAP7_75t_L g295 ( .A(n_206), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_206), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_206), .B(n_252), .Y(n_328) );
OR2x2_ASAP7_75t_L g366 ( .A(n_206), .B(n_321), .Y(n_366) );
AOI32xp33_ASAP7_75t_L g378 ( .A1(n_206), .A2(n_379), .A3(n_382), .B1(n_383), .B2(n_384), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_206), .B(n_354), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_206), .B(n_314), .Y(n_429) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AOI21xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_209), .B(n_216), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g244 ( .A(n_215), .Y(n_244) );
INVx1_ASAP7_75t_L g259 ( .A(n_216), .Y(n_259) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_216), .A2(n_508), .B(n_517), .Y(n_507) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_216), .A2(n_522), .B(n_529), .Y(n_521) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g340 ( .A(n_220), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
INVx1_ASAP7_75t_L g302 ( .A(n_221), .Y(n_302) );
AND2x2_ASAP7_75t_L g304 ( .A(n_221), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_221), .B(n_251), .Y(n_321) );
AND2x2_ASAP7_75t_L g354 ( .A(n_221), .B(n_330), .Y(n_354) );
AND2x2_ASAP7_75t_L g391 ( .A(n_221), .B(n_252), .Y(n_391) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_222), .B(n_251), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_222), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g329 ( .A(n_222), .B(n_330), .Y(n_329) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_232), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_230), .Y(n_226) );
INVx2_ASAP7_75t_L g305 ( .A(n_234), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_234), .B(n_251), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_234), .B(n_296), .Y(n_377) );
INVx1_ASAP7_75t_L g399 ( .A(n_234), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_234), .Y(n_416) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g269 ( .A(n_235), .B(n_251), .Y(n_269) );
AND2x2_ASAP7_75t_L g291 ( .A(n_235), .B(n_252), .Y(n_291) );
INVx1_ASAP7_75t_L g330 ( .A(n_235), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_241), .B(n_243), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_241), .A2(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g512 ( .A(n_241), .Y(n_512) );
AOI221x1_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_262), .B1(n_268), .B2(n_270), .C(n_271), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_247), .A2(n_335), .B1(n_402), .B2(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
AND2x2_ASAP7_75t_L g293 ( .A(n_248), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g388 ( .A(n_248), .B(n_268), .Y(n_388) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g344 ( .A(n_249), .B(n_269), .Y(n_344) );
INVx1_ASAP7_75t_L g356 ( .A(n_250), .Y(n_356) );
AND2x2_ASAP7_75t_L g367 ( .A(n_250), .B(n_354), .Y(n_367) );
AND2x2_ASAP7_75t_L g434 ( .A(n_250), .B(n_329), .Y(n_434) );
INVx2_ASAP7_75t_L g296 ( .A(n_251), .Y(n_296) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_259), .B(n_260), .Y(n_252) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_263), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_263), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_264), .B(n_347), .Y(n_350) );
INVx3_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_265), .A2(n_386), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_268), .B(n_294), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_269), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g360 ( .A(n_269), .B(n_288), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_269), .B(n_295), .Y(n_437) );
AND2x2_ASAP7_75t_L g306 ( .A(n_270), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g373 ( .A(n_270), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_280), .Y(n_271) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_273), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g322 ( .A(n_273), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g334 ( .A(n_273), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_273), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g358 ( .A(n_274), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_274), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_274), .B(n_277), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_277), .A2(n_316), .B(n_346), .C(n_348), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_277), .A2(n_364), .B1(n_367), .B2(n_368), .C(n_372), .Y(n_363) );
AND2x2_ASAP7_75t_L g359 ( .A(n_278), .B(n_312), .Y(n_359) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g319 ( .A(n_283), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g390 ( .A(n_283), .B(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_292), .C(n_317), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g403 ( .A(n_285), .B(n_404), .C(n_405), .Y(n_403) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
OR2x2_ASAP7_75t_L g376 ( .A(n_287), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_297), .B1(n_300), .B2(n_306), .C(n_308), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_294), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_294), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_299), .A2(n_356), .B1(n_357), .B2(n_358), .Y(n_355) );
OR2x2_ASAP7_75t_L g436 ( .A(n_299), .B(n_347), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVxp67_ASAP7_75t_L g410 ( .A(n_302), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_304), .B(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g311 ( .A(n_305), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_307), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_307), .B(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_307), .B(n_374), .Y(n_413) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_311), .Y(n_337) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g427 ( .A(n_316), .B(n_347), .Y(n_427) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g405 ( .A(n_322), .Y(n_405) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI322xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_331), .A3(n_332), .B1(n_333), .B2(n_336), .C1(n_338), .C2(n_340), .Y(n_325) );
OAI322xp33_ASAP7_75t_L g407 ( .A1(n_326), .A2(n_408), .A3(n_409), .B1(n_410), .B2(n_411), .C1(n_412), .C2(n_414), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx4_ASAP7_75t_L g341 ( .A(n_328), .Y(n_341) );
AND2x2_ASAP7_75t_L g402 ( .A(n_328), .B(n_354), .Y(n_402) );
AND2x2_ASAP7_75t_L g415 ( .A(n_328), .B(n_416), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_331), .Y(n_426) );
INVx1_ASAP7_75t_L g404 ( .A(n_332), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g338 ( .A(n_334), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g421 ( .A(n_334), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_334), .B(n_375), .Y(n_432) );
OR2x2_ASAP7_75t_L g365 ( .A(n_337), .B(n_366), .Y(n_365) );
INVxp33_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g342 ( .A1(n_341), .A2(n_343), .B1(n_345), .B2(n_349), .C(n_351), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_341), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g425 ( .A(n_341), .Y(n_425) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx3_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AOI322xp5_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_373), .A3(n_390), .B1(n_392), .B2(n_393), .C1(n_396), .C2(n_400), .Y(n_389) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_359), .B2(n_360), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_385), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_378), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_366), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp33_ASAP7_75t_SL g383 ( .A(n_369), .B(n_380), .Y(n_383) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI322xp33_ASAP7_75t_L g423 ( .A1(n_371), .A2(n_424), .A3(n_426), .B1(n_427), .B2(n_428), .C1(n_430), .C2(n_433), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_381), .B(n_429), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_387), .B(n_389), .C(n_401), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_417), .C(n_423), .D(n_435), .Y(n_406) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx14_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx6_ASAP7_75t_L g731 ( .A(n_440), .Y(n_731) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_442), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_646), .Y(n_442) );
NAND5xp2_ASAP7_75t_L g443 ( .A(n_444), .B(n_565), .C(n_580), .D(n_606), .E(n_628), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g444 ( .A(n_445), .B(n_545), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_486), .B1(n_518), .B2(n_534), .C(n_535), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_478), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_447), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g722 ( .A(n_447), .Y(n_722) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_459), .Y(n_447) );
INVx1_ASAP7_75t_L g562 ( .A(n_448), .Y(n_562) );
AND2x2_ASAP7_75t_L g564 ( .A(n_448), .B(n_472), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_448), .B(n_471), .Y(n_574) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_448), .Y(n_592) );
INVx1_ASAP7_75t_L g602 ( .A(n_448), .Y(n_602) );
OR2x2_ASAP7_75t_L g640 ( .A(n_448), .B(n_539), .Y(n_640) );
INVx2_ASAP7_75t_L g690 ( .A(n_448), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_448), .B(n_538), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_453), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_461), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_461), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_SL g622 ( .A(n_461), .B(n_562), .Y(n_622) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_462), .Y(n_480) );
INVx2_ASAP7_75t_L g539 ( .A(n_462), .Y(n_539) );
OR2x2_ASAP7_75t_L g601 ( .A(n_462), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g540 ( .A(n_471), .B(n_482), .Y(n_540) );
AND2x2_ASAP7_75t_L g557 ( .A(n_471), .B(n_537), .Y(n_557) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g481 ( .A(n_472), .B(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g560 ( .A(n_472), .Y(n_560) );
AND2x2_ASAP7_75t_L g689 ( .A(n_472), .B(n_690), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_475), .A2(n_503), .B(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_475), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_477), .A2(n_523), .B(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
AND2x2_ASAP7_75t_L g652 ( .A(n_479), .B(n_540), .Y(n_652) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g653 ( .A(n_480), .B(n_564), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_481), .A2(n_621), .B(n_623), .C(n_625), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_481), .B(n_621), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_481), .A2(n_551), .B1(n_694), .B2(n_695), .C(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g537 ( .A(n_482), .Y(n_537) );
INVx1_ASAP7_75t_L g573 ( .A(n_482), .Y(n_573) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_482), .Y(n_582) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
AND2x2_ASAP7_75t_L g599 ( .A(n_488), .B(n_544), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_488), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_489), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g691 ( .A(n_489), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g723 ( .A(n_489), .Y(n_723) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g553 ( .A(n_490), .Y(n_553) );
AND2x2_ASAP7_75t_L g579 ( .A(n_490), .B(n_533), .Y(n_579) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_490), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g595 ( .A(n_490), .B(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_496), .B(n_635), .Y(n_670) );
INVx1_ASAP7_75t_SL g674 ( .A(n_496), .Y(n_674) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
INVx3_ASAP7_75t_L g533 ( .A(n_497), .Y(n_533) );
AND2x2_ASAP7_75t_L g544 ( .A(n_497), .B(n_521), .Y(n_544) );
AND2x2_ASAP7_75t_L g566 ( .A(n_497), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g611 ( .A(n_497), .B(n_605), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_497), .B(n_543), .Y(n_692) );
INVx2_ASAP7_75t_L g514 ( .A(n_505), .Y(n_514) );
AND2x2_ASAP7_75t_L g532 ( .A(n_507), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g543 ( .A(n_507), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_507), .B(n_521), .Y(n_568) );
AND2x2_ASAP7_75t_L g604 ( .A(n_507), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_532), .Y(n_519) );
INVx1_ASAP7_75t_L g584 ( .A(n_520), .Y(n_584) );
AND2x2_ASAP7_75t_L g626 ( .A(n_520), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_520), .B(n_547), .Y(n_632) );
AOI21xp5_ASAP7_75t_SL g706 ( .A1(n_520), .A2(n_538), .B(n_561), .Y(n_706) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
OR2x2_ASAP7_75t_L g549 ( .A(n_521), .B(n_530), .Y(n_549) );
AND2x2_ASAP7_75t_L g596 ( .A(n_521), .B(n_533), .Y(n_596) );
INVx2_ASAP7_75t_L g605 ( .A(n_521), .Y(n_605) );
INVx1_ASAP7_75t_L g711 ( .A(n_521), .Y(n_711) );
AND2x2_ASAP7_75t_L g635 ( .A(n_530), .B(n_605), .Y(n_635) );
INVx1_ASAP7_75t_L g660 ( .A(n_530), .Y(n_660) );
AND2x2_ASAP7_75t_L g569 ( .A(n_532), .B(n_553), .Y(n_569) );
AND2x2_ASAP7_75t_L g581 ( .A(n_532), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g699 ( .A(n_532), .Y(n_699) );
INVx2_ASAP7_75t_L g589 ( .A(n_533), .Y(n_589) );
AND2x2_ASAP7_75t_L g627 ( .A(n_533), .B(n_543), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_533), .B(n_711), .Y(n_710) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_540), .B(n_541), .Y(n_535) );
AND2x2_ASAP7_75t_L g642 ( .A(n_536), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g696 ( .A(n_536), .Y(n_696) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g616 ( .A(n_537), .Y(n_616) );
BUFx2_ASAP7_75t_L g715 ( .A(n_537), .Y(n_715) );
BUFx2_ASAP7_75t_L g586 ( .A(n_538), .Y(n_586) );
AND2x2_ASAP7_75t_L g688 ( .A(n_538), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g671 ( .A(n_539), .Y(n_671) );
AND2x4_ASAP7_75t_L g598 ( .A(n_540), .B(n_561), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_540), .B(n_622), .Y(n_634) );
AOI32xp33_ASAP7_75t_L g558 ( .A1(n_541), .A2(n_559), .A3(n_561), .B1(n_563), .B2(n_564), .Y(n_558) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
INVx3_ASAP7_75t_L g547 ( .A(n_542), .Y(n_547) );
OR2x2_ASAP7_75t_L g683 ( .A(n_542), .B(n_639), .Y(n_683) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g552 ( .A(n_543), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g659 ( .A(n_543), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g551 ( .A(n_544), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g563 ( .A(n_544), .B(n_553), .Y(n_563) );
INVx1_ASAP7_75t_L g684 ( .A(n_544), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_544), .B(n_659), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_550), .B(n_554), .C(n_558), .Y(n_545) );
OAI322xp33_ASAP7_75t_L g654 ( .A1(n_546), .A2(n_591), .A3(n_655), .B1(n_657), .B2(n_661), .C1(n_662), .C2(n_666), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVxp67_ASAP7_75t_L g619 ( .A(n_547), .Y(n_619) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g673 ( .A(n_549), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_549), .B(n_589), .Y(n_720) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g612 ( .A(n_552), .Y(n_612) );
OR2x2_ASAP7_75t_L g698 ( .A(n_553), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_556), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g607 ( .A(n_557), .B(n_586), .Y(n_607) );
AND2x2_ASAP7_75t_L g678 ( .A(n_557), .B(n_591), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_557), .B(n_665), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_559), .A2(n_566), .B1(n_569), .B2(n_570), .C(n_575), .Y(n_565) );
OR2x2_ASAP7_75t_L g576 ( .A(n_559), .B(n_572), .Y(n_576) );
AND2x2_ASAP7_75t_L g664 ( .A(n_559), .B(n_665), .Y(n_664) );
AOI32xp33_ASAP7_75t_L g703 ( .A1(n_559), .A2(n_589), .A3(n_704), .B1(n_705), .B2(n_708), .Y(n_703) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_560), .B(n_596), .C(n_619), .Y(n_637) );
AND2x2_ASAP7_75t_L g663 ( .A(n_560), .B(n_656), .Y(n_663) );
INVxp67_ASAP7_75t_L g643 ( .A(n_561), .Y(n_643) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_564), .B(n_616), .Y(n_672) );
INVx2_ASAP7_75t_L g682 ( .A(n_564), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_564), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g651 ( .A(n_567), .Y(n_651) );
OR2x2_ASAP7_75t_L g577 ( .A(n_568), .B(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_570), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_573), .Y(n_656) );
AND2x2_ASAP7_75t_L g615 ( .A(n_574), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g661 ( .A(n_574), .Y(n_661) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_574), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI21xp33_ASAP7_75t_SL g600 ( .A1(n_576), .A2(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g694 ( .A(n_579), .B(n_604), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .B(n_593), .C(n_600), .Y(n_580) );
AND2x2_ASAP7_75t_L g624 ( .A(n_582), .B(n_592), .Y(n_624) );
INVx2_ASAP7_75t_L g639 ( .A(n_582), .Y(n_639) );
OR2x2_ASAP7_75t_L g677 ( .A(n_582), .B(n_640), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_582), .B(n_720), .Y(n_719) );
AOI211xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_585), .B(n_587), .C(n_590), .Y(n_583) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_586), .B(n_624), .Y(n_623) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_587), .A2(n_682), .B(n_706), .C(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_588), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g645 ( .A(n_589), .B(n_635), .Y(n_645) );
INVx1_ASAP7_75t_L g650 ( .A(n_589), .Y(n_650) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_597), .Y(n_593) );
INVxp33_ASAP7_75t_L g701 ( .A(n_595), .Y(n_701) );
AND2x2_ASAP7_75t_L g680 ( .A(n_596), .B(n_659), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_601), .A2(n_663), .B(n_664), .Y(n_662) );
OAI322xp33_ASAP7_75t_L g681 ( .A1(n_603), .A2(n_682), .A3(n_683), .B1(n_684), .B2(n_685), .C1(n_687), .C2(n_691), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_613), .B2(n_617), .C(n_620), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g658 ( .A(n_611), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g702 ( .A(n_615), .Y(n_702) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_618), .B(n_638), .Y(n_704) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g667 ( .A(n_627), .B(n_635), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_633), .B2(n_635), .C(n_636), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_631), .A2(n_648), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_647) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_635), .B(n_650), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_641), .B2(n_644), .Y(n_636) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx2_ASAP7_75t_SL g665 ( .A(n_640), .Y(n_665) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_647), .B(n_668), .C(n_693), .D(n_703), .E(n_713), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_649), .B(n_651), .Y(n_648) );
NOR4xp25_ASAP7_75t_L g721 ( .A(n_650), .B(n_656), .C(n_722), .D(n_723), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_653), .A2(n_714), .B1(n_716), .B2(n_718), .C(n_721), .Y(n_713) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g712 ( .A(n_659), .Y(n_712) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_663), .A2(n_670), .A3(n_671), .B1(n_672), .B2(n_673), .C1(n_675), .C2(n_679), .Y(n_669) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_681), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g714 ( .A(n_689), .B(n_715), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_697) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g750 ( .A(n_737), .Y(n_750) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g754 ( .A(n_748), .Y(n_754) );
BUFx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule