module fake_netlist_1_3358_n_447 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_447);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_447;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_58;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_SL g58 ( .A(n_51), .Y(n_58) );
INVxp67_ASAP7_75t_SL g59 ( .A(n_36), .Y(n_59) );
BUFx6f_ASAP7_75t_L g60 ( .A(n_4), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_11), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_54), .Y(n_62) );
INVxp67_ASAP7_75t_SL g63 ( .A(n_47), .Y(n_63) );
INVxp33_ASAP7_75t_L g64 ( .A(n_50), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_57), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_23), .Y(n_66) );
INVxp33_ASAP7_75t_L g67 ( .A(n_56), .Y(n_67) );
INVxp33_ASAP7_75t_L g68 ( .A(n_24), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_0), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_30), .Y(n_70) );
CKINVDCx20_ASAP7_75t_R g71 ( .A(n_39), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_41), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_27), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_46), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_11), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_12), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_49), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_42), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_55), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_9), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_9), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_6), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_5), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_14), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_17), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_6), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_3), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_31), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_19), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_5), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_71), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_85), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_85), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_77), .Y(n_99) );
BUFx2_ASAP7_75t_L g100 ( .A(n_85), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_83), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_58), .B(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
INVx4_ASAP7_75t_L g104 ( .A(n_60), .Y(n_104) );
INVx3_ASAP7_75t_L g105 ( .A(n_77), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_62), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_64), .B(n_1), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_95), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_65), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_60), .Y(n_110) );
NOR2xp33_ASAP7_75t_R g111 ( .A(n_74), .B(n_34), .Y(n_111) );
NAND2xp33_ASAP7_75t_R g112 ( .A(n_91), .B(n_2), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_58), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_67), .B(n_2), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_68), .B(n_3), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_61), .B(n_4), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_113), .B(n_78), .Y(n_117) );
OR2x2_ASAP7_75t_SL g118 ( .A(n_113), .B(n_98), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_101), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_105), .Y(n_120) );
AND2x6_ASAP7_75t_L g121 ( .A(n_107), .B(n_65), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_99), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_99), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_100), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_100), .B(n_61), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_99), .Y(n_127) );
OAI221xp5_ASAP7_75t_L g128 ( .A1(n_116), .A2(n_76), .B1(n_87), .B2(n_69), .C(n_75), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_104), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_107), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_101), .B(n_66), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_101), .B(n_66), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_110), .A2(n_76), .B1(n_80), .B2(n_86), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_96), .A2(n_84), .B1(n_94), .B2(n_80), .Y(n_137) );
INVxp67_ASAP7_75t_SL g138 ( .A(n_107), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_98), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_105), .Y(n_140) );
NOR2xp33_ASAP7_75t_R g141 ( .A(n_134), .B(n_112), .Y(n_141) );
O2A1O1Ixp5_ASAP7_75t_L g142 ( .A1(n_133), .A2(n_115), .B(n_102), .C(n_103), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_130), .B(n_100), .Y(n_143) );
OR2x6_ASAP7_75t_L g144 ( .A(n_125), .B(n_116), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
AND2x4_ASAP7_75t_SL g146 ( .A(n_126), .B(n_103), .Y(n_146) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
NOR3xp33_ASAP7_75t_SL g151 ( .A(n_137), .B(n_112), .C(n_115), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_138), .B(n_106), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_130), .B(n_106), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_125), .B(n_109), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_126), .B(n_111), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_126), .B(n_109), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_139), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_121), .A2(n_102), .B1(n_114), .B2(n_87), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_121), .B(n_114), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVxp67_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
AO22x1_ASAP7_75t_L g166 ( .A1(n_121), .A2(n_93), .B1(n_63), .B2(n_59), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_117), .B(n_93), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_126), .B(n_105), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_134), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_157), .A2(n_128), .B1(n_132), .B2(n_137), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx1_ASAP7_75t_SL g174 ( .A(n_146), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
INVx8_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_163), .Y(n_178) );
CKINVDCx8_ASAP7_75t_R g179 ( .A(n_144), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_146), .B(n_135), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_144), .B(n_69), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_157), .B(n_105), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
INVx5_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_157), .A2(n_105), .B1(n_99), .B2(n_97), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_158), .B(n_118), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_152), .A2(n_97), .B(n_88), .C(n_82), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_147), .B(n_129), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_157), .B(n_154), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_162), .A2(n_89), .B(n_70), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_154), .B(n_75), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_154), .B(n_81), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_136), .B(n_131), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_193), .A2(n_148), .B1(n_145), .B2(n_143), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_179), .A2(n_147), .B1(n_145), .B2(n_154), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_179), .A2(n_171), .B1(n_147), .B2(n_152), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_188), .B(n_118), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_193), .B(n_143), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_179), .A2(n_169), .B1(n_162), .B2(n_165), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_186), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_193), .A2(n_143), .B1(n_141), .B2(n_168), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_180), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_177), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_180), .A2(n_156), .B(n_169), .Y(n_213) );
INVx1_ASAP7_75t_SL g214 ( .A(n_174), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_188), .B(n_143), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_180), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_188), .B(n_153), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_173), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_176), .A2(n_170), .B(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_193), .B(n_153), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_193), .B(n_151), .Y(n_223) );
OAI221xp5_ASAP7_75t_L g224 ( .A1(n_172), .A2(n_151), .B1(n_161), .B2(n_142), .C(n_165), .Y(n_224) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_199), .A2(n_160), .B(n_164), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_167), .B1(n_159), .B2(n_170), .Y(n_226) );
BUFx10_ASAP7_75t_L g227 ( .A(n_193), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_186), .A2(n_166), .B1(n_81), .B2(n_82), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_205), .A2(n_177), .B1(n_182), .B2(n_183), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_209), .Y(n_230) );
AOI22xp33_ASAP7_75t_SL g231 ( .A1(n_212), .A2(n_177), .B1(n_189), .B2(n_186), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_211), .A2(n_189), .B1(n_177), .B2(n_186), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_227), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_212), .A2(n_186), .B1(n_177), .B2(n_189), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_215), .B(n_183), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_210), .A2(n_182), .B1(n_177), .B2(n_183), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_216), .B(n_184), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_216), .Y(n_239) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_225), .A2(n_191), .B(n_199), .Y(n_240) );
AOI221xp5_ASAP7_75t_L g241 ( .A1(n_217), .A2(n_172), .B1(n_191), .B2(n_198), .C(n_196), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g242 ( .A1(n_204), .A2(n_177), .B1(n_186), .B2(n_182), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_217), .A2(n_196), .B1(n_198), .B2(n_184), .C(n_88), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_206), .A2(n_183), .B1(n_186), .B2(n_198), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_214), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_176), .B(n_190), .Y(n_247) );
OAI221xp5_ASAP7_75t_L g248 ( .A1(n_203), .A2(n_142), .B1(n_187), .B2(n_196), .C(n_184), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_206), .A2(n_183), .B1(n_186), .B2(n_175), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_209), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g251 ( .A1(n_244), .A2(n_215), .B1(n_224), .B2(n_223), .C(n_222), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_239), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_239), .B(n_219), .Y(n_253) );
OAI211xp5_ASAP7_75t_L g254 ( .A1(n_241), .A2(n_86), .B(n_94), .C(n_187), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_244), .A2(n_183), .B1(n_228), .B2(n_207), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_239), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_233), .A2(n_219), .B(n_220), .Y(n_257) );
OAI211xp5_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_213), .B(n_92), .C(n_79), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_233), .B(n_220), .Y(n_259) );
OAI211xp5_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_90), .B(n_79), .C(n_89), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_233), .B(n_195), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_247), .A2(n_221), .B(n_218), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
OAI33xp33_ASAP7_75t_L g264 ( .A1(n_232), .A2(n_70), .A3(n_72), .B1(n_73), .B2(n_92), .B3(n_90), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_229), .A2(n_208), .B1(n_197), .B2(n_190), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_248), .A2(n_166), .B1(n_60), .B2(n_197), .C(n_195), .Y(n_267) );
AOI33xp33_ASAP7_75t_L g268 ( .A1(n_245), .A2(n_72), .A3(n_73), .B1(n_77), .B2(n_124), .B3(n_127), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_238), .B(n_195), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_247), .Y(n_270) );
NOR2x1_ASAP7_75t_SL g271 ( .A(n_232), .B(n_202), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_266), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_252), .Y(n_274) );
OAI31xp33_ASAP7_75t_L g275 ( .A1(n_260), .A2(n_235), .A3(n_248), .B(n_234), .Y(n_275) );
OAI33xp33_ASAP7_75t_L g276 ( .A1(n_265), .A2(n_236), .A3(n_226), .B1(n_10), .B2(n_12), .B3(n_13), .Y(n_276) );
NAND4xp25_ASAP7_75t_L g277 ( .A(n_254), .B(n_237), .C(n_249), .D(n_242), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_252), .B(n_246), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_256), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_256), .B(n_247), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_270), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_270), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_255), .A2(n_242), .B1(n_231), .B2(n_234), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_253), .B(n_243), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_259), .B(n_238), .Y(n_288) );
OAI31xp33_ASAP7_75t_L g289 ( .A1(n_258), .A2(n_243), .A3(n_236), .B(n_175), .Y(n_289) );
OAI221xp5_ASAP7_75t_L g290 ( .A1(n_251), .A2(n_231), .B1(n_250), .B2(n_218), .C(n_60), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_240), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_266), .B(n_250), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_269), .B(n_240), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_271), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
OAI21xp5_ASAP7_75t_SL g298 ( .A1(n_255), .A2(n_218), .B(n_175), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_265), .B(n_240), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_293), .A2(n_262), .B(n_257), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_291), .B(n_240), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_291), .B(n_240), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_295), .B(n_297), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_290), .A2(n_264), .B(n_267), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_278), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_292), .B(n_262), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_278), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_292), .B(n_60), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_295), .B(n_230), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_299), .B(n_60), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_299), .B(n_230), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_294), .B(n_230), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_294), .B(n_230), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_287), .B(n_230), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_288), .B(n_268), .Y(n_317) );
OAI31xp33_ASAP7_75t_SL g318 ( .A1(n_283), .A2(n_250), .A3(n_8), .B(n_10), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_273), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_287), .B(n_230), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_272), .B(n_7), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_284), .B(n_195), .Y(n_324) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_297), .B(n_175), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_281), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_273), .B(n_52), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_285), .B(n_195), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_282), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_285), .B(n_7), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_286), .B(n_13), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_284), .B(n_14), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_282), .B(n_15), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_273), .B(n_15), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_275), .B(n_298), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_277), .A2(n_276), .B1(n_289), .B2(n_227), .Y(n_339) );
OR2x4_ASAP7_75t_L g340 ( .A(n_295), .B(n_200), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_323), .A2(n_192), .B(n_124), .C(n_127), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_338), .A2(n_227), .B1(n_192), .B2(n_104), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_306), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_309), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_319), .Y(n_346) );
OAI222xp33_ASAP7_75t_L g347 ( .A1(n_338), .A2(n_16), .B1(n_17), .B2(n_18), .C1(n_19), .C2(n_20), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_319), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_304), .Y(n_349) );
OAI31xp33_ASAP7_75t_L g350 ( .A1(n_333), .A2(n_16), .A3(n_18), .B(n_20), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_127), .B(n_131), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_334), .A2(n_104), .B1(n_123), .B2(n_122), .C(n_124), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_311), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_339), .A2(n_104), .B1(n_201), .B2(n_202), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g357 ( .A1(n_332), .A2(n_111), .B(n_136), .C(n_122), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_321), .B(n_104), .Y(n_359) );
AOI21xp33_ASAP7_75t_SL g360 ( .A1(n_332), .A2(n_21), .B(n_22), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_303), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
INVx4_ASAP7_75t_L g365 ( .A(n_320), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_303), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_340), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_317), .B(n_25), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_337), .A2(n_122), .B(n_131), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_326), .A2(n_123), .B1(n_194), .B2(n_202), .C(n_185), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_326), .B(n_123), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_335), .A2(n_123), .B1(n_194), .B2(n_185), .C(n_181), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_314), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_330), .B(n_26), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_337), .A2(n_194), .B1(n_185), .B2(n_181), .Y(n_377) );
OR2x6_ASAP7_75t_SL g378 ( .A(n_330), .B(n_28), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_301), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_379), .B(n_301), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_343), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_374), .B(n_307), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_354), .B(n_312), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g385 ( .A1(n_347), .A2(n_305), .B(n_329), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_349), .B(n_302), .Y(n_386) );
NAND2xp33_ASAP7_75t_R g387 ( .A(n_360), .B(n_329), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_365), .B(n_320), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_329), .B(n_325), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_367), .A2(n_329), .B(n_310), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_353), .B(n_314), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_365), .B(n_310), .Y(n_392) );
XNOR2xp5_ASAP7_75t_L g393 ( .A(n_362), .B(n_315), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_358), .B(n_324), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_345), .B(n_315), .Y(n_395) );
NAND2x1_ASAP7_75t_SL g396 ( .A(n_365), .B(n_310), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_350), .A2(n_300), .B(n_310), .Y(n_397) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_367), .B(n_312), .Y(n_398) );
XOR2xp5_ASAP7_75t_L g399 ( .A(n_375), .B(n_322), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_366), .B(n_316), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_361), .B(n_29), .Y(n_403) );
XNOR2x1_ASAP7_75t_L g404 ( .A(n_356), .B(n_32), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_346), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_181), .B(n_178), .C(n_194), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_400), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_380), .B(n_369), .Y(n_411) );
NAND4xp75_ASAP7_75t_L g412 ( .A(n_385), .B(n_368), .C(n_342), .D(n_376), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g413 ( .A1(n_402), .A2(n_370), .B1(n_377), .B2(n_346), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_386), .B(n_348), .Y(n_414) );
NOR2xp33_ASAP7_75t_SL g415 ( .A(n_402), .B(n_351), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_392), .A2(n_372), .B(n_359), .Y(n_416) );
AOI31xp33_ASAP7_75t_L g417 ( .A1(n_387), .A2(n_373), .A3(n_371), .B(n_352), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_388), .B(n_341), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_396), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_200), .B1(n_37), .B2(n_38), .Y(n_420) );
OAI321xp33_ASAP7_75t_L g421 ( .A1(n_389), .A2(n_200), .A3(n_40), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_391), .B(n_35), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_405), .Y(n_423) );
OAI21xp33_ASAP7_75t_SL g424 ( .A1(n_419), .A2(n_398), .B(n_382), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_413), .A2(n_409), .B(n_383), .C(n_381), .Y(n_425) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_410), .A2(n_384), .A3(n_401), .B1(n_406), .B2(n_407), .C1(n_386), .C2(n_394), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_412), .A2(n_399), .B1(n_393), .B2(n_395), .Y(n_427) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_420), .B(n_404), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_414), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_418), .A2(n_394), .B1(n_408), .B2(n_403), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_423), .A2(n_417), .B1(n_411), .B2(n_414), .C(n_416), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_411), .A2(n_402), .B1(n_378), .B2(n_413), .Y(n_432) );
INVxp33_ASAP7_75t_SL g433 ( .A(n_421), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_413), .A2(n_402), .B1(n_412), .B2(n_415), .Y(n_434) );
OAI311xp33_ASAP7_75t_L g435 ( .A1(n_422), .A2(n_402), .A3(n_385), .B1(n_397), .C1(n_339), .Y(n_435) );
XNOR2xp5_ASAP7_75t_L g436 ( .A(n_432), .B(n_434), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_429), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_431), .B(n_426), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_427), .A2(n_425), .B1(n_433), .B2(n_430), .Y(n_439) );
NOR2xp67_ASAP7_75t_L g440 ( .A(n_436), .B(n_424), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_437), .Y(n_441) );
XOR2xp5_ASAP7_75t_L g442 ( .A(n_439), .B(n_428), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_442), .B(n_438), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_441), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g445 ( .A(n_443), .B(n_440), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_445), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_446), .A2(n_444), .B(n_435), .Y(n_447) );
endmodule