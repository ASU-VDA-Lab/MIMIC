module fake_jpeg_7490_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_28),
.B1(n_20),
.B2(n_33),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_20),
.B1(n_16),
.B2(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_23),
.B(n_25),
.C(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx2_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_23),
.B(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_90),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_76),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_17),
.Y(n_103)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_75),
.B1(n_78),
.B2(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_84),
.B1(n_89),
.B2(n_32),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_21),
.B1(n_28),
.B2(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_18),
.C(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_91),
.Y(n_101)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_16),
.B1(n_17),
.B2(n_31),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_45),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g145 ( 
.A(n_92),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_0),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_116),
.B1(n_88),
.B2(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_60),
.B1(n_47),
.B2(n_58),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_90),
.B1(n_80),
.B2(n_74),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_22),
.B(n_24),
.C(n_54),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_108),
.A3(n_116),
.B1(n_115),
.B2(n_101),
.Y(n_142)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_24),
.B(n_83),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_26),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_31),
.B1(n_26),
.B2(n_19),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_26),
.B1(n_22),
.B2(n_33),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_70),
.B1(n_30),
.B2(n_67),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_77),
.B1(n_65),
.B2(n_9),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_43),
.C(n_63),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_19),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_30),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_83),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_43),
.B1(n_24),
.B2(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_77),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_49),
.C(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_135),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_134),
.B1(n_140),
.B2(n_142),
.Y(n_169)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_133),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_123),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_76),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_88),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_85),
.B1(n_73),
.B2(n_83),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_103),
.B1(n_116),
.B2(n_109),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_99),
.B1(n_111),
.B2(n_116),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_77),
.B1(n_65),
.B2(n_9),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_65),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_159),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_104),
.B(n_102),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_176),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_162),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_94),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_15),
.B(n_11),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_93),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_167),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_112),
.C(n_93),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_4),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_100),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_145),
.C(n_120),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_8),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_95),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_0),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_132),
.B(n_119),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_1),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_1),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_3),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_129),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_181),
.B(n_188),
.Y(n_208)
);

XOR2x2_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_145),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_201),
.C(n_204),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_145),
.B1(n_146),
.B2(n_100),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_145),
.B1(n_130),
.B2(n_133),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_130),
.B(n_2),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_194),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_171),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_192),
.B1(n_196),
.B2(n_175),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_199),
.B1(n_163),
.B2(n_168),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_10),
.B1(n_11),
.B2(n_15),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_173),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_10),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_3),
.B(n_4),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_4),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_165),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_218),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_165),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_156),
.B1(n_155),
.B2(n_168),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_230),
.C(n_180),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_222),
.Y(n_247)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_228),
.B(n_229),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_148),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_176),
.B(n_150),
.C(n_161),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_232),
.A2(n_199),
.B1(n_190),
.B2(n_202),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_208),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_241),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_240),
.C(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_198),
.C(n_189),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_207),
.B(n_198),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_182),
.B(n_158),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_215),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_177),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_231),
.C(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_250),
.C(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_251),
.A2(n_209),
.B1(n_213),
.B2(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_232),
.B1(n_241),
.B2(n_222),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_219),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_258),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_225),
.CI(n_233),
.CON(n_260),
.SN(n_260)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_249),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_267),
.B1(n_268),
.B2(n_243),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_209),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_236),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_211),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_266),
.B1(n_202),
.B2(n_157),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_177),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_272),
.C(n_275),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_247),
.C(n_245),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_236),
.C(n_252),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_265),
.C(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_277),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_282),
.B1(n_255),
.B2(n_220),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_260),
.C(n_226),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_223),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_273),
.B1(n_280),
.B2(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_261),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_149),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_293),
.Y(n_297)
);

OAI211xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_291),
.B(n_260),
.C(n_221),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_153),
.B(n_149),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_167),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_301),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_157),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_285),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_307),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_285),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_309),
.B(n_297),
.Y(n_311)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_304),
.B(n_293),
.C(n_305),
.D(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_312),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_310),
.B(n_305),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_304),
.B(n_296),
.C(n_271),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_174),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_200),
.B(n_6),
.Y(n_318)
);


endmodule