module real_jpeg_24418_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_0),
.A2(n_38),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_0),
.A2(n_47),
.B1(n_65),
.B2(n_66),
.Y(n_170)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_2),
.A2(n_38),
.B1(n_41),
.B2(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_3),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_37),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_50),
.C(n_52),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_3),
.A2(n_38),
.B1(n_41),
.B2(n_161),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_108),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_161),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_3),
.B(n_65),
.C(n_80),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_3),
.A2(n_67),
.B(n_222),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_27),
.B1(n_38),
.B2(n_41),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_27),
.B1(n_65),
.B2(n_66),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_9),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_12),
.A2(n_38),
.B1(n_41),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_12),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_72),
.Y(n_125)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_16),
.Y(n_171)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_143),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_141),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_20),
.B(n_120),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_98),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_25),
.B(n_44),
.C(n_60),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_37),
.B2(n_42),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_28),
.A2(n_35),
.A3(n_41),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_29),
.Y(n_160)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_32),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_32),
.A2(n_138),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_34),
.B(n_38),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_36),
.B(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_38),
.B(n_186),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_42),
.Y(n_135)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_46),
.A2(n_48),
.B1(n_58),
.B2(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_48),
.A2(n_54),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_50),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_50),
.B(n_229),
.Y(n_228)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_55),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_106),
.B1(n_108),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_58),
.A2(n_107),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_76),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_61),
.B(n_76),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_71),
.B2(n_73),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_110)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_68),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_66),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_66),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_71),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_73),
.B(n_88),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_67),
.A2(n_113),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_67),
.B(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_67),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_74),
.B(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_75),
.B(n_161),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_77),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_77),
.A2(n_210),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_94),
.B1(n_95),
.B2(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_78),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_78),
.A2(n_95),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_82),
.A2(n_83),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_82),
.A2(n_154),
.B(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_82),
.B(n_161),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_86),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_95),
.B(n_155),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_98),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_109),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_99),
.B(n_104),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_109),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_115),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_111),
.A2(n_233),
.B1(n_235),
.B2(n_237),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_140),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_139),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B(n_137),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_178),
.B(n_265),
.C(n_270),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_172),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_163),
.C(n_164),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_146),
.A2(n_147),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_152),
.C(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B(n_162),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_163),
.B(n_164),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_171),
.A2(n_234),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_259),
.B(n_264),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_211),
.B(n_258),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_200),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_183),
.B(n_200),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_193),
.C(n_197),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_184),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_187),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B(n_191),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_193),
.A2(n_197),
.B1(n_198),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_263)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_252),
.B(n_257),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_230),
.B(n_251),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_224),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_224),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_228),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_240),
.B(n_250),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_238),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);


endmodule