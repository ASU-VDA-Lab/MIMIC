module fake_jpeg_15066_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_59),
.Y(n_74)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_22),
.B1(n_28),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_79),
.B1(n_37),
.B2(n_39),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_70),
.B(n_76),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_78),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_28),
.B1(n_42),
.B2(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_96),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_42),
.B1(n_61),
.B2(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_105),
.B1(n_41),
.B2(n_27),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_64),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_44),
.CON(n_103),
.SN(n_103)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_123),
.B(n_45),
.Y(n_148)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_27),
.B1(n_41),
.B2(n_46),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_126),
.Y(n_147)
);

BUFx4f_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_116),
.B1(n_124),
.B2(n_43),
.Y(n_128)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_39),
.B1(n_60),
.B2(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_117),
.B1(n_88),
.B2(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_26),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_34),
.B1(n_31),
.B2(n_35),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_21),
.B1(n_29),
.B2(n_34),
.Y(n_117)
);

OA22x2_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_59),
.B1(n_56),
.B2(n_48),
.Y(n_118)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_36),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_32),
.Y(n_151)
);

CKINVDCx11_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_0),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_29),
.B1(n_21),
.B2(n_31),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_26),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_36),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_128),
.Y(n_167)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_73),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_153),
.B(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_149),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_81),
.B1(n_86),
.B2(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_141),
.B1(n_93),
.B2(n_108),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_81),
.B1(n_90),
.B2(n_75),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_144),
.Y(n_172)
);

OAI221xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_45),
.B1(n_32),
.B2(n_43),
.C(n_33),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_33),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_106),
.A2(n_98),
.B1(n_112),
.B2(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_122),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_109),
.C(n_95),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_25),
.C(n_142),
.Y(n_200)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_171),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_180),
.B1(n_148),
.B2(n_147),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_103),
.B(n_118),
.C(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_75),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_174),
.A2(n_113),
.B1(n_158),
.B2(n_31),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_141),
.B1(n_150),
.B2(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_157),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_195),
.C(n_200),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_150),
.B1(n_165),
.B2(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_202),
.B1(n_170),
.B2(n_113),
.Y(n_209)
);

NOR2x1p5_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_118),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_185),
.B(n_192),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_130),
.B(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_191),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_152),
.B1(n_146),
.B2(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_193),
.B1(n_194),
.B2(n_180),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_135),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_146),
.B1(n_151),
.B2(n_133),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_140),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_145),
.B(n_127),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_142),
.B(n_176),
.C(n_179),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_154),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_166),
.B1(n_170),
.B2(n_169),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_59),
.B1(n_107),
.B2(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_129),
.B1(n_131),
.B2(n_137),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_229),
.B1(n_10),
.B2(n_19),
.Y(n_237)
);

OAI22x1_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_168),
.B1(n_161),
.B2(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_228),
.Y(n_240)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_160),
.B1(n_166),
.B2(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_224),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_201),
.B(n_35),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_172),
.B1(n_173),
.B2(n_179),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_181),
.B1(n_188),
.B2(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_199),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_181),
.A2(n_144),
.B1(n_139),
.B2(n_107),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_107),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_0),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_139),
.C(n_25),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_213),
.C(n_229),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_181),
.A2(n_35),
.B1(n_34),
.B2(n_59),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_200),
.B1(n_202),
.B2(n_201),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_232),
.A2(n_217),
.B(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_212),
.C(n_220),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_245),
.B1(n_246),
.B2(n_2),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_25),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_238),
.B(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

NOR4xp25_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_9),
.C(n_16),
.D(n_3),
.Y(n_244)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_1),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_224),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_215),
.B(n_18),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_10),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_16),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_254),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_223),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_213),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_278),
.C(n_231),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_241),
.C(n_240),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_236),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_217),
.B1(n_216),
.B2(n_203),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_10),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_217),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_277),
.B1(n_243),
.B2(n_247),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_217),
.B1(n_7),
.B2(n_8),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_5),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_230),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_231),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_293),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_267),
.B1(n_276),
.B2(n_258),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_289),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_257),
.B(n_235),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_294),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_261),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_239),
.C(n_248),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_241),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_237),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_240),
.Y(n_296)
);

AOI221xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_272),
.B1(n_277),
.B2(n_258),
.C(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_254),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_260),
.C(n_270),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_311),
.C(n_238),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_308),
.B1(n_244),
.B2(n_280),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_275),
.B1(n_276),
.B2(n_267),
.Y(n_303)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_260),
.B(n_266),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_310),
.B(n_279),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_263),
.B1(n_265),
.B2(n_253),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_285),
.B(n_290),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_243),
.C(n_263),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_262),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_311),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_317),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_292),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_319),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_281),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_305),
.B(n_269),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_324),
.B(n_307),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_309),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_246),
.C(n_245),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_5),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_325),
.B(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_304),
.Y(n_330)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_322),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_332),
.A2(n_333),
.B(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_315),
.A2(n_310),
.B(n_7),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_323),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_337),
.B(n_334),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_340),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_5),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_344),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_329),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_342),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_8),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_332),
.C(n_326),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_350),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_11),
.B(n_13),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_342),
.B(n_14),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_349),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);

AOI322xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_353),
.A3(n_348),
.B1(n_345),
.B2(n_354),
.C1(n_346),
.C2(n_338),
.Y(n_357)
);

NOR4xp25_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_15),
.C(n_13),
.D(n_14),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_13),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_15),
.Y(n_360)
);


endmodule