module real_jpeg_32938_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx3_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_0),
.Y(n_110)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_36),
.B1(n_40),
.B2(n_45),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_45),
.B1(n_99),
.B2(n_103),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_2),
.A2(n_62),
.B1(n_256),
.B2(n_261),
.Y(n_255)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_67),
.A3(n_73),
.B1(n_77),
.B2(n_85),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_86),
.B1(n_197),
.B2(n_202),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_3),
.B(n_137),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_3),
.A2(n_95),
.B1(n_289),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_5),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_6),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_7),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_7),
.A2(n_132),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_7),
.A2(n_132),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_9),
.A2(n_147),
.B1(n_150),
.B2(n_153),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_9),
.A2(n_153),
.B1(n_240),
.B2(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_9),
.A2(n_153),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_171),
.B1(n_172),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_217),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_215),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_123),
.B(n_190),
.C(n_191),
.Y(n_16)
);

AOI211xp5_ASAP7_75t_L g216 ( 
.A1(n_17),
.A2(n_123),
.B(n_190),
.C(n_191),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_18),
.B(n_125),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_65),
.B1(n_121),
.B2(n_122),
.Y(n_18)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_19),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_35),
.B1(n_46),
.B2(n_60),
.Y(n_19)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_20),
.A2(n_238),
.B1(n_247),
.B2(n_248),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_20),
.B(n_86),
.Y(n_300)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_21),
.A2(n_61),
.B1(n_206),
.B2(n_214),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_22),
.A2(n_46),
.B1(n_207),
.B2(n_238),
.Y(n_268)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AO21x2_ASAP7_75t_L g46 ( 
.A1(n_24),
.A2(n_47),
.B(n_53),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_24)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_27),
.Y(n_175)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_29),
.Y(n_231)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_39),
.Y(n_244)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_43),
.Y(n_213)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_44),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_46),
.Y(n_214)
);

NAND2xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_53),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_92),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_66),
.A2(n_92),
.B1(n_93),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_66),
.Y(n_193)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_72),
.Y(n_204)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_77),
.A2(n_138),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_86),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_86),
.B(n_233),
.Y(n_232)
);

OA21x2_ASAP7_75t_SL g248 ( 
.A1(n_86),
.A2(n_232),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_86),
.B(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_90),
.Y(n_236)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B1(n_107),
.B2(n_111),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_111),
.B1(n_166),
.B2(n_170),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_94),
.A2(n_274),
.B1(n_281),
.B2(n_282),
.Y(n_273)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_95),
.A2(n_255),
.B1(n_262),
.B2(n_265),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_95),
.A2(n_275),
.B1(n_289),
.B2(n_296),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_98),
.Y(n_265)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_102),
.Y(n_278)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_105),
.Y(n_308)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_110),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_110),
.Y(n_284)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_115),
.Y(n_224)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_119),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_120),
.Y(n_295)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_163),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_136),
.B1(n_146),
.B2(n_154),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_136),
.A2(n_146),
.B1(n_154),
.B2(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_179),
.B2(n_180),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_168),
.Y(n_307)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_178),
.Y(n_291)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_205),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_192),
.B(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_194),
.A2(n_195),
.B1(n_205),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_205),
.Y(n_316)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_214),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21x1_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_312),
.B(n_317),
.Y(n_218)
);

OAI21x1_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_271),
.B(n_311),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_253),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_221),
.B(n_253),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_237),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_222),
.B(n_237),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.B(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_230),
.B(n_232),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx4f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_266),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_254),
.B(n_268),
.C(n_269),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_286),
.B(n_310),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_285),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_285),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_301),
.B(n_309),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_300),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);


endmodule