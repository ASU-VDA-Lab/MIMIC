module real_jpeg_33041_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_653;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_0),
.A2(n_115),
.B1(n_117),
.B2(n_120),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_0),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_0),
.A2(n_120),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_0),
.A2(n_120),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_0),
.A2(n_120),
.B1(n_542),
.B2(n_544),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_1),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_1),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_3),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_3),
.A2(n_237),
.B1(n_413),
.B2(n_416),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_3),
.A2(n_237),
.B1(n_484),
.B2(n_487),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_3),
.A2(n_237),
.B1(n_601),
.B2(n_602),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_4),
.A2(n_129),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_4),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_4),
.A2(n_230),
.B1(n_288),
.B2(n_292),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_4),
.A2(n_230),
.B1(n_441),
.B2(n_446),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_4),
.A2(n_222),
.B1(n_230),
.B2(n_565),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_5),
.A2(n_349),
.B1(n_354),
.B2(n_356),
.Y(n_348)
);

INVx2_ASAP7_75t_R g356 ( 
.A(n_5),
.Y(n_356)
);

AO22x1_ASAP7_75t_L g422 ( 
.A1(n_5),
.A2(n_356),
.B1(n_423),
.B2(n_425),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_5),
.A2(n_356),
.B1(n_495),
.B2(n_498),
.Y(n_494)
);

AO22x1_ASAP7_75t_L g592 ( 
.A1(n_5),
.A2(n_356),
.B1(n_593),
.B2(n_595),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_5),
.A2(n_356),
.B1(n_611),
.B2(n_612),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_6),
.A2(n_332),
.B1(n_334),
.B2(n_337),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_6),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_6),
.A2(n_337),
.B1(n_384),
.B2(n_389),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_6),
.A2(n_337),
.B1(n_470),
.B2(n_472),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_6),
.A2(n_337),
.B1(n_558),
.B2(n_560),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_7),
.A2(n_231),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_7),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_7),
.A2(n_299),
.B1(n_376),
.B2(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_7),
.A2(n_299),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_7),
.A2(n_299),
.B1(n_569),
.B2(n_571),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_35),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_8),
.A2(n_35),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_8),
.A2(n_35),
.B1(n_208),
.B2(n_275),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_11),
.Y(n_353)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_11),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_12),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_12),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_12),
.A2(n_128),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_12),
.A2(n_128),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_12),
.A2(n_128),
.B1(n_506),
.B2(n_508),
.Y(n_505)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_13),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_14),
.A2(n_64),
.B1(n_67),
.B2(n_73),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_14),
.A2(n_73),
.B1(n_103),
.B2(n_108),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_73),
.B1(n_166),
.B2(n_169),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_14),
.A2(n_73),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

CKINVDCx11_ASAP7_75t_R g658 ( 
.A(n_15),
.Y(n_658)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_16),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_17),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_18),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_18),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_19),
.A2(n_197),
.B1(n_278),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_19),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_19),
.B(n_164),
.Y(n_427)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_19),
.A2(n_143),
.A3(n_449),
.B1(n_451),
.B2(n_455),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_19),
.A2(n_340),
.B1(n_465),
.B2(n_467),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_19),
.B(n_238),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_19),
.A2(n_535),
.B(n_554),
.Y(n_553)
);

OAI311xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_178),
.A3(n_184),
.B1(n_655),
.C1(n_657),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_22),
.B(n_178),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_177),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_74),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_25),
.B(n_74),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_61),
.B2(n_63),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_26),
.A2(n_37),
.B1(n_61),
.B2(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_30),
.Y(n_239)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_34),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_34),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_37),
.A2(n_114),
.B1(n_121),
.B2(n_123),
.Y(n_113)
);

OAI22x1_ASAP7_75t_SL g295 ( 
.A1(n_37),
.A2(n_62),
.B1(n_296),
.B2(n_300),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_37),
.A2(n_62),
.B1(n_553),
.B2(n_557),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_37),
.A2(n_62),
.B1(n_296),
.B2(n_610),
.Y(n_609)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_38),
.A2(n_122),
.B1(n_229),
.B2(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_38),
.A2(n_122),
.B1(n_124),
.B2(n_229),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_38),
.A2(n_122),
.B1(n_592),
.B2(n_598),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_51),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_39)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_40),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_40),
.Y(n_612)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_41),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_41),
.Y(n_556)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_42),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_42),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_43),
.Y(n_597)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_46),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_50),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_55),
.Y(n_252)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_57),
.Y(n_533)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_58),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_60),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_60),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_R g509 ( 
.A(n_62),
.B(n_340),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_70),
.Y(n_232)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_72),
.Y(n_236)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_72),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_173),
.C(n_176),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_75),
.A2(n_76),
.B1(n_646),
.B2(n_647),
.Y(n_645)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_113),
.C(n_132),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_77),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_77),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g321 ( 
.A(n_77),
.B(n_133),
.Y(n_321)
);

AO21x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_88),
.B(n_102),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_78),
.A2(n_88),
.B1(n_212),
.B2(n_219),
.Y(n_211)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_78),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_78),
.A2(n_88),
.B1(n_212),
.B2(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_78),
.B(n_340),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_78),
.A2(n_88),
.B1(n_482),
.B2(n_483),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_78),
.A2(n_88),
.B1(n_483),
.B2(n_564),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_78),
.A2(n_88),
.B1(n_266),
.B2(n_564),
.Y(n_582)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AO21x2_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_89),
.B(n_94),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_83),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_83),
.Y(n_277)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_85),
.Y(n_333)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_92),
.Y(n_395)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_92),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_93),
.Y(n_269)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_93),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_94),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_98),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_98),
.Y(n_272)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_102),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_103),
.B(n_340),
.Y(n_455)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_106),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_107),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_111),
.Y(n_218)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_111),
.Y(n_486)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_112),
.Y(n_392)
);

XOR2x1_ASAP7_75t_L g320 ( 
.A(n_113),
.B(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_158),
.B1(n_163),
.B2(n_165),
.Y(n_133)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_134),
.A2(n_158),
.B1(n_163),
.B2(n_309),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_134),
.A2(n_163),
.B1(n_464),
.B2(n_469),
.Y(n_463)
);

OAI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_134),
.A2(n_163),
.B1(n_469),
.B2(n_494),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_134),
.A2(n_163),
.B1(n_494),
.B2(n_568),
.Y(n_567)
);

OA22x2_ASAP7_75t_L g599 ( 
.A1(n_134),
.A2(n_163),
.B1(n_568),
.B2(n_600),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_134),
.A2(n_163),
.B1(n_287),
.B2(n_600),
.Y(n_613)
);

AO21x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_143),
.B(n_149),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_136),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_145),
.Y(n_466)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_145),
.Y(n_572)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_155),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_150),
.Y(n_566)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_164),
.A2(n_174),
.B1(n_243),
.B2(n_250),
.Y(n_242)
);

AOI22x1_ASAP7_75t_L g285 ( 
.A1(n_164),
.A2(n_174),
.B1(n_243),
.B2(n_286),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g454 ( 
.A(n_172),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_173),
.B(n_176),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_178),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_184),
.B(n_656),
.Y(n_655)
);

OAI31xp33_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_322),
.A3(n_644),
.B(n_649),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_314),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_301),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_188),
.B(n_301),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_240),
.C(n_262),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2x1_ASAP7_75t_L g633 ( 
.A(n_190),
.B(n_241),
.Y(n_633)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_226),
.Y(n_190)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_191),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_211),
.Y(n_191)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_192),
.A2(n_228),
.B(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_192),
.A2(n_227),
.B1(n_624),
.B2(n_625),
.Y(n_623)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_204),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_195),
.Y(n_342)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_197),
.A2(n_274),
.B1(n_278),
.B2(n_283),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_197),
.A2(n_331),
.B1(n_348),
.B2(n_357),
.Y(n_347)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_197),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_197),
.A2(n_399),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_197),
.A2(n_274),
.B1(n_541),
.B2(n_584),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_200),
.Y(n_439)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_200),
.Y(n_539)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g345 ( 
.A(n_202),
.Y(n_345)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_202),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_203),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_211),
.Y(n_625)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

BUFx4f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_233),
.Y(n_300)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_256),
.B(n_261),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_256),
.Y(n_261)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_249),
.Y(n_474)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_258),
.A2(n_259),
.B1(n_383),
.B2(n_393),
.Y(n_382)
);

NAND2x1_ASAP7_75t_SL g421 ( 
.A(n_258),
.B(n_422),
.Y(n_421)
);

AOI22x1_ASAP7_75t_L g458 ( 
.A1(n_258),
.A2(n_259),
.B1(n_422),
.B2(n_459),
.Y(n_458)
);

NAND2x1_ASAP7_75t_L g420 ( 
.A(n_259),
.B(n_383),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_262),
.B(n_633),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_284),
.C(n_294),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_263),
.A2(n_264),
.B1(n_627),
.B2(n_628),
.Y(n_626)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_265),
.B(n_273),
.Y(n_616)
);

BUFx6f_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_269),
.Y(n_424)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_272),
.Y(n_426)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_277),
.Y(n_543)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_277),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_282),
.Y(n_410)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_282),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g627 ( 
.A(n_285),
.B(n_295),
.Y(n_627)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_291),
.Y(n_471)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_291),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_293),
.Y(n_497)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_293),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_310),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_311),
.C(n_313),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_304),
.B(n_318),
.C(n_320),
.Y(n_648)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_315),
.A2(n_652),
.B(n_653),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g653 ( 
.A(n_316),
.B(n_317),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_575),
.B(n_639),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_513),
.B(n_574),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_476),
.B(n_512),
.Y(n_324)
);

AOI21x1_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_429),
.B(n_475),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_406),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_361),
.B(n_403),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_346),
.B(n_360),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_338),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_336),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_373),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_SL g393 ( 
.A1(n_340),
.A2(n_372),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_398),
.B1(n_401),
.B2(n_402),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_359),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_347),
.B(n_359),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_352),
.Y(n_507)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_397),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_381),
.B1(n_382),
.B2(n_396),
.Y(n_362)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g404 ( 
.A(n_363),
.B(n_381),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_371),
.B1(n_375),
.B2(n_380),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_381),
.B(n_396),
.Y(n_407)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_396),
.Y(n_405)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_397),
.A2(n_404),
.B(n_405),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AO22x1_ASAP7_75t_L g436 ( 
.A1(n_401),
.A2(n_412),
.B1(n_437),
.B2(n_440),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_401),
.A2(n_440),
.B1(n_503),
.B2(n_505),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_401),
.A2(n_505),
.B1(n_537),
.B2(n_540),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_407),
.A2(n_430),
.B(n_431),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_408),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_419),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g432 ( 
.A(n_409),
.B(n_427),
.C(n_433),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B(n_427),
.C(n_428),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_421),
.C(n_427),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_R g433 ( 
.A(n_420),
.B(n_421),
.Y(n_433)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

NOR2x1_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_432),
.B(n_434),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_456),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_435),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_448),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_448),
.Y(n_480)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_SL g468 ( 
.A(n_453),
.Y(n_468)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_454),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_462),
.B2(n_463),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_462),
.C(n_511),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_460),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_470),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_510),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_510),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_491),
.B2(n_492),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_480),
.A2(n_481),
.B1(n_489),
.B2(n_490),
.Y(n_479)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_480),
.Y(n_490)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_481),
.B(n_490),
.C(n_491),
.Y(n_573)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_501),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_493),
.B(n_509),
.C(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_500),
.Y(n_570)
);

XNOR2x1_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_509),
.Y(n_501)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_502),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_573),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_514),
.B(n_573),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_550),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_548),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_548),
.C(n_550),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_536),
.B1(n_546),
.B2(n_547),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_517),
.B(n_547),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_517),
.B(n_547),
.Y(n_615)
);

OAI32xp33_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_520),
.A3(n_523),
.B1(n_527),
.B2(n_534),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx3_ASAP7_75t_SL g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_536),
.Y(n_547)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx2_ASAP7_75t_SL g544 ( 
.A(n_545),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_551),
.B(n_562),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_SL g580 ( 
.A(n_552),
.B(n_563),
.C(n_567),
.Y(n_580)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx3_ASAP7_75t_SL g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_557),
.Y(n_598)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_567),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

NAND4xp25_ASAP7_75t_SL g575 ( 
.A(n_576),
.B(n_603),
.C(n_629),
.D(n_634),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_577),
.B(n_578),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_577),
.B(n_578),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_588),
.Y(n_578)
);

XNOR2x1_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_581),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_580),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_581),
.B(n_588),
.C(n_636),
.Y(n_635)
);

XOR2x2_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_583),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_582),
.B(n_583),
.Y(n_607)
);

INVx3_ASAP7_75t_SL g584 ( 
.A(n_585),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

XNOR2x1_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_590),
.Y(n_588)
);

XNOR2x1_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_599),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_591),
.B(n_599),
.C(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_597),
.Y(n_596)
);

A2O1A1O1Ixp25_ASAP7_75t_L g639 ( 
.A1(n_603),
.A2(n_629),
.B(n_640),
.C(n_642),
.D(n_643),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_604),
.B(n_617),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_604),
.B(n_617),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_614),
.C(n_616),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_606),
.B(n_616),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_608),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_619),
.C(n_621),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_609),
.B(n_613),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_609),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_613),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_614),
.B(n_638),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_622),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_623),
.C(n_631),
.Y(n_630)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_626),
.Y(n_622)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_626),
.Y(n_631)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_627),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_632),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_630),
.B(n_632),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_635),
.B(n_637),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_635),
.B(n_637),
.C(n_641),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_644),
.A2(n_651),
.B(n_654),
.Y(n_650)
);

NOR2x1_ASAP7_75t_R g644 ( 
.A(n_645),
.B(n_648),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_645),
.B(n_648),
.Y(n_654)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_658),
.B(n_659),
.Y(n_657)
);


endmodule