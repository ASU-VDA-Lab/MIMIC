module fake_netlist_5_988_n_108 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_108);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_108;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVxp33_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx2_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_7),
.Y(n_48)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_29),
.B1(n_5),
.B2(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI221xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_29),
.B1(n_34),
.B2(n_22),
.C(n_24),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_4),
.B1(n_5),
.B2(n_20),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_26),
.B1(n_31),
.B2(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_48),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_52),
.B(n_57),
.C(n_44),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_59),
.Y(n_71)
);

OR2x6_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_65),
.B(n_68),
.C(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_78),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AO21x2_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_68),
.B(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_78),
.B1(n_49),
.B2(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_72),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_88),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_86),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_38),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_38),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_48),
.B(n_37),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_40),
.B(n_45),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_98),
.B1(n_100),
.B2(n_48),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_103),
.B1(n_40),
.B2(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_13),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_40),
.B1(n_45),
.B2(n_18),
.C(n_19),
.Y(n_108)
);


endmodule