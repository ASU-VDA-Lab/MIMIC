module real_jpeg_25534_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_0),
.B(n_69),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_54),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_59),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_0),
.B(n_28),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_0),
.B(n_45),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_69),
.Y(n_96)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_59),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_3),
.B(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_28),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_42),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_4),
.B(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_4),
.B(n_59),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_17),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_4),
.B(n_28),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_8),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_9),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_9),
.B(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_9),
.B(n_54),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_59),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_9),
.B(n_69),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_9),
.B(n_28),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_45),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_13),
.B(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_13),
.B(n_59),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_13),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_14),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_14),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_42),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_16),
.B(n_54),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_16),
.B(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_16),
.B(n_69),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_16),
.B(n_28),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_16),
.B(n_50),
.Y(n_238)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_155),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_132),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_63),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_22),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_48),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_23),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_30),
.C(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_40),
.A2(n_41),
.B(n_44),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_40),
.B(n_48),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_42),
.Y(n_222)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_43),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_55),
.Y(n_48)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_49),
.B(n_53),
.CI(n_55),
.CON(n_136),
.SN(n_136)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_56),
.B(n_63),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_61),
.C(n_62),
.Y(n_121)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_59),
.Y(n_217)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.C(n_73),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_64),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.C(n_68),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_65),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_66),
.B(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_67),
.B(n_68),
.Y(n_259)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_98),
.B2(n_131),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_88),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_86),
.B1(n_90),
.B2(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_90),
.C(n_91),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_92),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_94),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.CI(n_97),
.CON(n_94),
.SN(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_120),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.C(n_116),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_105),
.C(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_106),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_116),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.C(n_114),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_130),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_151),
.C(n_153),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_133),
.A2(n_134),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_147),
.C(n_149),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_135),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.C(n_143),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_136),
.B(n_252),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_136),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_143),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_144),
.B(n_145),
.CI(n_146),
.CON(n_233),
.SN(n_233)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_147),
.B(n_149),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_151),
.B(n_153),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_272),
.C(n_273),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_262),
.C(n_263),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_245),
.C(n_246),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_227),
.C(n_228),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_187),
.C(n_199),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_174),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_169),
.C(n_174),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_164),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_175),
.B(n_181),
.C(n_182),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_186),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_198),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_192),
.B1(n_198),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_223),
.C(n_224),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.C(n_214),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_206),
.C(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.C(n_218),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_235),
.C(n_244),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_232),
.C(n_233),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_233),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_244),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_238),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_250),
.C(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_258),
.C(n_260),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_257),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_258),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_268),
.C(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);


endmodule