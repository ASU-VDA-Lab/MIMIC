module real_aes_4038_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_1135, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_1134, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_1136, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_1133, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_1135;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_1134;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_1136;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_1133;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_1034;
wire n_923;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_884;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_976;
wire n_559;
wire n_636;
wire n_872;
wire n_1053;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_1081;
wire n_960;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_1031;
wire n_1037;
wire n_880;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1105;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_1033;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_968;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_717;
wire n_456;
wire n_1090;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1114;
wire n_465;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_1045;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_1104;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_0), .A2(n_273), .B1(n_414), .B2(n_430), .Y(n_742) );
INVx1_ASAP7_75t_L g712 ( .A(n_1), .Y(n_712) );
INVx1_ASAP7_75t_L g686 ( .A(n_2), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_3), .A2(n_226), .B1(n_358), .B2(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g802 ( .A(n_4), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_5), .A2(n_208), .B1(n_400), .B2(n_430), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_6), .A2(n_240), .B1(n_471), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g567 ( .A(n_7), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_8), .A2(n_256), .B1(n_514), .B2(n_515), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_9), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_10), .A2(n_244), .B1(n_390), .B2(n_396), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_11), .A2(n_125), .B1(n_566), .B2(n_569), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_12), .A2(n_179), .B1(n_358), .B2(n_828), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_13), .A2(n_235), .B1(n_445), .B2(n_676), .C(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_14), .A2(n_195), .B1(n_401), .B2(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g715 ( .A(n_15), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_16), .A2(n_17), .B1(n_519), .B2(n_756), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_18), .B(n_340), .Y(n_350) );
AOI21xp33_ASAP7_75t_L g790 ( .A1(n_19), .A2(n_595), .B(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_20), .A2(n_86), .B1(n_471), .B2(n_472), .Y(n_1091) );
INVx1_ASAP7_75t_L g710 ( .A(n_21), .Y(n_710) );
AOI221x1_ASAP7_75t_L g363 ( .A1(n_22), .A2(n_76), .B1(n_364), .B2(n_371), .C(n_374), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_23), .A2(n_239), .B1(n_471), .B2(n_583), .Y(n_644) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_24), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_25), .A2(n_26), .B1(n_517), .B2(n_519), .Y(n_516) );
INVx1_ASAP7_75t_L g532 ( .A(n_27), .Y(n_532) );
AOI21xp33_ASAP7_75t_L g837 ( .A1(n_28), .A2(n_541), .B(n_838), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_29), .A2(n_148), .B1(n_476), .B2(n_613), .Y(n_1090) );
INVx1_ASAP7_75t_L g747 ( .A(n_30), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_31), .A2(n_108), .B1(n_560), .B2(n_638), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_32), .A2(n_203), .B1(n_637), .B2(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_33), .A2(n_248), .B1(n_594), .B2(n_596), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_34), .A2(n_98), .B1(n_548), .B2(n_549), .Y(n_657) );
INVx1_ASAP7_75t_L g685 ( .A(n_35), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_36), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_37), .A2(n_257), .B1(n_515), .B2(n_759), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_38), .A2(n_138), .B1(n_883), .B2(n_891), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_39), .A2(n_251), .B1(n_464), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_40), .A2(n_189), .B1(n_358), .B2(n_487), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_41), .A2(n_48), .B1(n_517), .B2(n_757), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_42), .A2(n_118), .B1(n_548), .B2(n_549), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_43), .A2(n_120), .B1(n_486), .B2(n_487), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_44), .A2(n_281), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_45), .A2(n_201), .B1(n_515), .B2(n_759), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_46), .A2(n_191), .B1(n_756), .B2(n_757), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_47), .A2(n_294), .B1(n_536), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_49), .A2(n_282), .B1(n_423), .B2(n_536), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_50), .A2(n_93), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_51), .A2(n_598), .B(n_600), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g1116 ( .A1(n_52), .A2(n_306), .B1(n_472), .B2(n_521), .Y(n_1116) );
OA22x2_ASAP7_75t_L g345 ( .A1(n_53), .A2(n_137), .B1(n_340), .B2(n_344), .Y(n_345) );
INVx1_ASAP7_75t_L g386 ( .A(n_53), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_54), .A2(n_162), .B1(n_505), .B2(n_651), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_55), .A2(n_66), .B1(n_501), .B2(n_1094), .C(n_1095), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_56), .A2(n_269), .B1(n_401), .B2(n_409), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_57), .A2(n_97), .B1(n_505), .B2(n_789), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_58), .Y(n_412) );
INVx1_ASAP7_75t_L g870 ( .A(n_59), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_60), .A2(n_129), .B1(n_858), .B2(n_861), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_61), .A2(n_298), .B1(n_336), .B2(n_358), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_62), .A2(n_186), .B1(n_514), .B2(n_515), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_63), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g872 ( .A(n_64), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_65), .B(n_155), .Y(n_322) );
INVx1_ASAP7_75t_L g343 ( .A(n_65), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g403 ( .A1(n_65), .A2(n_137), .B(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_67), .A2(n_95), .B1(n_881), .B2(n_889), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_68), .A2(n_209), .B1(n_512), .B2(n_609), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_69), .A2(n_217), .B1(n_472), .B2(n_521), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_70), .A2(n_197), .B1(n_464), .B2(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g571 ( .A(n_71), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g1123 ( .A1(n_72), .A2(n_445), .B(n_1124), .Y(n_1123) );
XOR2x2_ASAP7_75t_L g550 ( .A(n_73), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g853 ( .A(n_74), .Y(n_853) );
AND2x4_ASAP7_75t_L g856 ( .A(n_74), .B(n_225), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_75), .A2(n_271), .B1(n_855), .B2(n_881), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_77), .A2(n_241), .B1(n_472), .B2(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g443 ( .A(n_78), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_79), .A2(n_132), .B1(n_464), .B2(n_708), .Y(n_761) );
INVx1_ASAP7_75t_L g575 ( .A(n_80), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_81), .A2(n_293), .B1(n_471), .B2(n_472), .Y(n_470) );
AO22x1_ASAP7_75t_L g1113 ( .A1(n_82), .A2(n_266), .B1(n_512), .B2(n_1114), .Y(n_1113) );
AO22x2_ASAP7_75t_L g880 ( .A1(n_83), .A2(n_247), .B1(n_855), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_84), .A2(n_106), .B1(n_390), .B2(n_396), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_85), .A2(n_127), .B1(n_708), .B2(n_834), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_87), .A2(n_188), .B1(n_505), .B2(n_708), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_88), .A2(n_101), .B1(n_499), .B2(n_560), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_89), .A2(n_124), .B1(n_517), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_90), .A2(n_115), .B1(n_861), .B2(n_901), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_91), .A2(n_249), .B1(n_474), .B2(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g749 ( .A(n_92), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_92), .A2(n_117), .B1(n_883), .B2(n_891), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_94), .A2(n_110), .B1(n_643), .B2(n_759), .Y(n_758) );
AND2x4_ASAP7_75t_L g854 ( .A(n_96), .B(n_318), .Y(n_854) );
INVx1_ASAP7_75t_L g860 ( .A(n_96), .Y(n_860) );
INVx1_ASAP7_75t_SL g884 ( .A(n_96), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_99), .A2(n_291), .B1(n_641), .B2(n_643), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g1126 ( .A(n_100), .B(n_599), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_102), .A2(n_107), .B1(n_514), .B2(n_643), .Y(n_1089) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_103), .A2(n_105), .B1(n_481), .B2(n_483), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_104), .B(n_539), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_109), .A2(n_122), .B1(n_855), .B2(n_881), .Y(n_896) );
INVx1_ASAP7_75t_L g776 ( .A(n_111), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_111), .A2(n_310), .B1(n_858), .B2(n_881), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_112), .A2(n_274), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_113), .A2(n_220), .B1(n_400), .B2(n_408), .Y(n_739) );
AO22x1_ASAP7_75t_L g806 ( .A1(n_114), .A2(n_270), .B1(n_474), .B2(n_486), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_116), .A2(n_199), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_119), .A2(n_213), .B1(n_364), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_121), .A2(n_216), .B1(n_408), .B2(n_544), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_123), .A2(n_194), .B1(n_573), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_126), .A2(n_128), .B1(n_486), .B2(n_487), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_130), .B(n_599), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_131), .A2(n_255), .B1(n_472), .B2(n_521), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_133), .A2(n_147), .B1(n_487), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_134), .A2(n_279), .B1(n_507), .B2(n_508), .Y(n_506) );
CKINVDCx6p67_ASAP7_75t_R g439 ( .A(n_135), .Y(n_439) );
INVx1_ASAP7_75t_L g357 ( .A(n_136), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_136), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_136), .B(n_183), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_137), .B(n_234), .Y(n_321) );
XNOR2x1_ASAP7_75t_L g734 ( .A(n_138), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g824 ( .A(n_139), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_140), .A2(n_145), .B1(n_486), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_141), .A2(n_146), .B1(n_449), .B2(n_1099), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_142), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_143), .A2(n_158), .B1(n_336), .B2(n_409), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_144), .A2(n_212), .B1(n_474), .B2(n_486), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_149), .A2(n_231), .B1(n_519), .B2(n_756), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_150), .Y(n_670) );
INVx1_ASAP7_75t_L g564 ( .A(n_151), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_152), .A2(n_308), .B1(n_445), .B2(n_569), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_153), .A2(n_164), .B1(n_560), .B2(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g680 ( .A(n_154), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_155), .B(n_349), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_156), .A2(n_174), .B1(n_483), .B2(n_487), .Y(n_584) );
INVx1_ASAP7_75t_L g683 ( .A(n_157), .Y(n_683) );
XNOR2x1_ASAP7_75t_L g626 ( .A(n_159), .B(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_160), .A2(n_307), .B1(n_617), .B2(n_618), .Y(n_616) );
INVxp33_ASAP7_75t_SL g876 ( .A(n_161), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_163), .A2(n_254), .B1(n_474), .B2(n_476), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_165), .Y(n_425) );
INVx1_ASAP7_75t_L g839 ( .A(n_166), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_167), .A2(n_193), .B1(n_472), .B2(n_521), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_168), .B(n_566), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_169), .A2(n_297), .B1(n_336), .B2(n_544), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_170), .A2(n_311), .B1(n_708), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_171), .A2(n_295), .B1(n_849), .B2(n_855), .Y(n_848) );
INVx1_ASAP7_75t_L g704 ( .A(n_172), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_173), .A2(n_301), .B1(n_541), .B2(n_562), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_175), .A2(n_267), .B1(n_481), .B2(n_723), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_176), .A2(n_205), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_177), .A2(n_232), .B1(n_408), .B2(n_409), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_178), .A2(n_250), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_180), .A2(n_230), .B1(n_336), .B2(n_427), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_181), .B(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_182), .A2(n_292), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g341 ( .A(n_183), .Y(n_341) );
INVx1_ASAP7_75t_L g798 ( .A(n_184), .Y(n_798) );
OAI222xp33_ASAP7_75t_L g807 ( .A1(n_184), .A2(n_808), .B1(n_811), .B2(n_812), .C1(n_1135), .C2(n_1136), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_184), .B(n_812), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_185), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_187), .A2(n_290), .B1(n_400), .B2(n_408), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_190), .A2(n_206), .B1(n_474), .B2(n_623), .Y(n_645) );
XNOR2x1_ASAP7_75t_L g587 ( .A(n_192), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_196), .B(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_198), .A2(n_210), .B1(n_371), .B2(n_445), .C(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g1096 ( .A(n_200), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_202), .A2(n_296), .B1(n_423), .B2(n_541), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_204), .A2(n_289), .B1(n_858), .B2(n_885), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_207), .A2(n_268), .B1(n_481), .B2(n_483), .Y(n_691) );
INVx1_ASAP7_75t_L g457 ( .A(n_211), .Y(n_457) );
INVx1_ASAP7_75t_L g792 ( .A(n_214), .Y(n_792) );
INVx1_ASAP7_75t_L g601 ( .A(n_215), .Y(n_601) );
INVx1_ASAP7_75t_L g674 ( .A(n_218), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_219), .A2(n_246), .B1(n_514), .B2(n_515), .Y(n_721) );
INVx1_ASAP7_75t_L g554 ( .A(n_221), .Y(n_554) );
INVx1_ASAP7_75t_L g765 ( .A(n_222), .Y(n_765) );
AO22x1_ASAP7_75t_L g882 ( .A1(n_223), .A2(n_229), .B1(n_883), .B2(n_885), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_224), .A2(n_262), .B1(n_481), .B2(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_225), .Y(n_323) );
AND2x4_ASAP7_75t_L g852 ( .A(n_225), .B(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_227), .A2(n_233), .B1(n_401), .B2(n_409), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_228), .Y(n_421) );
INVx1_ASAP7_75t_L g355 ( .A(n_234), .Y(n_355) );
INVxp67_ASAP7_75t_L g420 ( .A(n_234), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_236), .A2(n_300), .B1(n_612), .B2(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g1125 ( .A(n_237), .Y(n_1125) );
INVx1_ASAP7_75t_L g447 ( .A(n_238), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_242), .A2(n_277), .B1(n_471), .B2(n_583), .Y(n_811) );
INVx2_ASAP7_75t_L g318 ( .A(n_243), .Y(n_318) );
INVxp33_ASAP7_75t_SL g979 ( .A(n_245), .Y(n_979) );
INVx1_ASAP7_75t_SL g362 ( .A(n_252), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_252), .B(n_436), .C(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g706 ( .A(n_253), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_258), .A2(n_261), .B1(n_423), .B2(n_430), .Y(n_537) );
AO221x2_ASAP7_75t_L g975 ( .A1(n_259), .A2(n_260), .B1(n_849), .B2(n_976), .C(n_977), .Y(n_975) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_263), .A2(n_427), .B(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_264), .A2(n_278), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_265), .A2(n_275), .B1(n_427), .B2(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g1085 ( .A(n_271), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_271), .A2(n_1107), .B1(n_1127), .B2(n_1129), .Y(n_1106) );
INVx1_ASAP7_75t_L g453 ( .A(n_272), .Y(n_453) );
XOR2xp5_ASAP7_75t_L g647 ( .A(n_276), .B(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_280), .A2(n_284), .B1(n_505), .B2(n_651), .Y(n_1120) );
INVx1_ASAP7_75t_L g522 ( .A(n_283), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_285), .A2(n_305), .B1(n_466), .B2(n_539), .Y(n_538) );
AO22x2_ASAP7_75t_L g698 ( .A1(n_286), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_286), .Y(n_699) );
AND2x2_ASAP7_75t_L g374 ( .A(n_287), .B(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_288), .A2(n_303), .B1(n_476), .B2(n_579), .Y(n_578) );
XNOR2xp5_ASAP7_75t_L g1107 ( .A(n_299), .B(n_1108), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_302), .A2(n_309), .B1(n_637), .B2(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g461 ( .A(n_304), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_324), .B(n_841), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_316), .B(n_1104), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_316), .B(n_1105), .Y(n_1128) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OA21x2_ASAP7_75t_L g1130 ( .A1(n_317), .A2(n_884), .B(n_1131), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g859 ( .A(n_318), .B(n_860), .Y(n_859) );
AND3x4_ASAP7_75t_L g883 ( .A(n_318), .B(n_852), .C(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_319), .B(n_1105), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g378 ( .A1(n_320), .A2(n_379), .B(n_381), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g1105 ( .A(n_323), .Y(n_1105) );
XNOR2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_664), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_585), .B1(n_662), .B2(n_663), .Y(n_325) );
INVx1_ASAP7_75t_L g662 ( .A(n_326), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_527), .B2(n_528), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AO22x2_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_490), .B1(n_523), .B2(n_524), .Y(n_328) );
INVx2_ASAP7_75t_L g523 ( .A(n_329), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_331), .B1(n_438), .B2(n_489), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2x1_ASAP7_75t_L g332 ( .A(n_333), .B(n_431), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_387), .C(n_406), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_362), .B1(n_363), .B2(n_1133), .Y(n_334) );
INVx1_ASAP7_75t_L g436 ( .A(n_335), .Y(n_436) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_346), .Y(n_336) );
AND2x4_ASAP7_75t_L g359 ( .A(n_337), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g373 ( .A(n_337), .B(n_368), .Y(n_373) );
AND2x4_ASAP7_75t_L g430 ( .A(n_337), .B(n_395), .Y(n_430) );
AND2x2_ASAP7_75t_L g451 ( .A(n_337), .B(n_395), .Y(n_451) );
AND2x2_ASAP7_75t_L g475 ( .A(n_337), .B(n_346), .Y(n_475) );
AND2x2_ASAP7_75t_L g518 ( .A(n_337), .B(n_346), .Y(n_518) );
AND2x2_ASAP7_75t_L g541 ( .A(n_337), .B(n_368), .Y(n_541) );
AND2x4_ASAP7_75t_L g544 ( .A(n_337), .B(n_405), .Y(n_544) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_345), .Y(n_337) );
INVx1_ASAP7_75t_L g367 ( .A(n_338), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
NAND2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx2_ASAP7_75t_L g344 ( .A(n_340), .Y(n_344) );
INVx3_ASAP7_75t_L g349 ( .A(n_340), .Y(n_349) );
NAND2xp33_ASAP7_75t_L g356 ( .A(n_340), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_340), .Y(n_380) );
INVx1_ASAP7_75t_L g404 ( .A(n_340), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_341), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_343), .A2(n_404), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g366 ( .A(n_345), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
AND2x2_ASAP7_75t_L g418 ( .A(n_345), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g408 ( .A(n_346), .B(n_393), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_346), .B(n_402), .Y(n_409) );
AND2x4_ASAP7_75t_L g478 ( .A(n_346), .B(n_402), .Y(n_478) );
AND2x4_ASAP7_75t_L g482 ( .A(n_346), .B(n_393), .Y(n_482) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_351), .Y(n_346) );
OR2x2_ASAP7_75t_L g361 ( .A(n_347), .B(n_352), .Y(n_361) );
INVx2_ASAP7_75t_L g369 ( .A(n_347), .Y(n_369) );
AND2x4_ASAP7_75t_L g395 ( .A(n_347), .B(n_370), .Y(n_395) );
AND2x2_ASAP7_75t_L g415 ( .A(n_347), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_349), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g381 ( .A(n_350), .B(n_382), .C(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g370 ( .A(n_353), .Y(n_370) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_359), .Y(n_486) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_359), .Y(n_512) );
BUFx12f_ASAP7_75t_L g615 ( .A(n_359), .Y(n_615) );
AND2x4_ASAP7_75t_L g400 ( .A(n_360), .B(n_393), .Y(n_400) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g405 ( .A(n_361), .Y(n_405) );
NOR2xp67_ASAP7_75t_L g387 ( .A(n_362), .B(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_362), .A2(n_407), .B1(n_410), .B2(n_1134), .Y(n_406) );
INVx1_ASAP7_75t_L g433 ( .A(n_363), .Y(n_433) );
BUFx8_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g456 ( .A(n_365), .Y(n_456) );
INVx2_ASAP7_75t_L g502 ( .A(n_365), .Y(n_502) );
BUFx3_ASAP7_75t_L g566 ( .A(n_365), .Y(n_566) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_365), .Y(n_595) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_365), .Y(n_651) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
AND2x4_ASAP7_75t_L g427 ( .A(n_366), .B(n_395), .Y(n_427) );
AND2x4_ASAP7_75t_L g446 ( .A(n_366), .B(n_395), .Y(n_446) );
AND2x2_ASAP7_75t_L g539 ( .A(n_366), .B(n_368), .Y(n_539) );
AND2x4_ASAP7_75t_L g393 ( .A(n_367), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_393), .Y(n_398) );
AND2x4_ASAP7_75t_L g423 ( .A(n_368), .B(n_402), .Y(n_423) );
AND2x4_ASAP7_75t_L g459 ( .A(n_368), .B(n_402), .Y(n_459) );
AND2x4_ASAP7_75t_L g549 ( .A(n_368), .B(n_393), .Y(n_549) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g462 ( .A(n_371), .Y(n_462) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g599 ( .A(n_372), .Y(n_599) );
INVx3_ASAP7_75t_SL g1094 ( .A(n_372), .Y(n_1094) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g507 ( .A(n_373), .Y(n_507) );
INVx2_ASAP7_75t_L g558 ( .A(n_373), .Y(n_558) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx4_ASAP7_75t_L g604 ( .A(n_377), .Y(n_604) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_378), .Y(n_467) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_380), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_383), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g402 ( .A(n_384), .B(n_403), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_388), .B(n_432), .C(n_435), .Y(n_431) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_399), .Y(n_388) );
BUFx4f_ASAP7_75t_L g582 ( .A(n_390), .Y(n_582) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_392), .Y(n_471) );
BUFx12f_ASAP7_75t_L g521 ( .A(n_392), .Y(n_521) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AND2x4_ASAP7_75t_L g484 ( .A(n_393), .B(n_405), .Y(n_484) );
AND2x4_ASAP7_75t_L g548 ( .A(n_393), .B(n_395), .Y(n_548) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_396), .Y(n_693) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_398), .Y(n_472) );
BUFx5_ASAP7_75t_L g583 ( .A(n_398), .Y(n_583) );
BUFx3_ASAP7_75t_L g619 ( .A(n_398), .Y(n_619) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
AND2x4_ASAP7_75t_L g488 ( .A(n_402), .B(n_405), .Y(n_488) );
INVx1_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
INVx1_ASAP7_75t_L g434 ( .A(n_410), .Y(n_434) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_424), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_421), .B2(n_422), .Y(n_411) );
INVx4_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
AND2x4_ASAP7_75t_L g465 ( .A(n_415), .B(n_418), .Y(n_465) );
AND2x2_ASAP7_75t_L g536 ( .A(n_415), .B(n_418), .Y(n_536) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_428), .B2(n_429), .Y(n_424) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_438), .Y(n_489) );
XNOR2x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_468), .Y(n_440) );
NOR3xp33_ASAP7_75t_SL g441 ( .A(n_442), .B(n_452), .C(n_460), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_444), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g504 ( .A(n_446), .Y(n_504) );
INVx1_ASAP7_75t_L g574 ( .A(n_446), .Y(n_574) );
BUFx3_ASAP7_75t_L g789 ( .A(n_446), .Y(n_789) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_450), .Y(n_633) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_451), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_457), .B2(n_458), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g596 ( .A(n_458), .Y(n_596) );
INVx3_ASAP7_75t_L g635 ( .A(n_458), .Y(n_635) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_459), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_463), .Y(n_460) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx5_ASAP7_75t_L g561 ( .A(n_465), .Y(n_561) );
BUFx4f_ASAP7_75t_L g834 ( .A(n_465), .Y(n_834) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
INVx2_ASAP7_75t_SL g562 ( .A(n_467), .Y(n_562) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_467), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_467), .B(n_747), .Y(n_746) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
BUFx8_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_475), .Y(n_613) );
INVx4_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
INVx1_ASAP7_75t_L g623 ( .A(n_477), .Y(n_623) );
INVx1_ASAP7_75t_L g695 ( .A(n_477), .Y(n_695) );
INVx4_ASAP7_75t_L g723 ( .A(n_477), .Y(n_723) );
INVx2_ASAP7_75t_SL g757 ( .A(n_477), .Y(n_757) );
INVx8_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_485), .Y(n_479) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx12f_ASAP7_75t_L g514 ( .A(n_482), .Y(n_514) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_482), .Y(n_759) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_483), .Y(n_607) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_484), .Y(n_515) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_484), .Y(n_643) );
BUFx12f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx6_ASAP7_75t_L g610 ( .A(n_488), .Y(n_610) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g526 ( .A(n_493), .Y(n_526) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
XOR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_522), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_497), .B(n_510), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .C(n_503), .D(n_506), .Y(n_497) );
INVx2_ASAP7_75t_L g576 ( .A(n_499), .Y(n_576) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g591 ( .A(n_504), .Y(n_591) );
INVx1_ASAP7_75t_L g705 ( .A(n_504), .Y(n_705) );
INVx3_ASAP7_75t_L g713 ( .A(n_505), .Y(n_713) );
INVx2_ASAP7_75t_L g677 ( .A(n_507), .Y(n_677) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_509), .B(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g1124 ( .A(n_509), .B(n_1125), .Y(n_1124) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .C(n_516), .D(n_520), .Y(n_510) );
BUFx12f_ASAP7_75t_L g579 ( .A(n_514), .Y(n_579) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_514), .Y(n_621) );
BUFx4f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_518), .Y(n_756) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
XNOR2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_550), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
XNOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_542), .Y(n_533) );
NAND4xp25_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .C(n_538), .D(n_540), .Y(n_534) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .C(n_546), .D(n_547), .Y(n_542) );
NAND2x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_577), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_563), .C(n_570), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_559), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g630 ( .A(n_557), .Y(n_630) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_561), .A2(n_601), .B(n_602), .Y(n_600) );
INVx4_ASAP7_75t_L g637 ( .A(n_561), .Y(n_637) );
INVx2_ASAP7_75t_L g1099 ( .A(n_561), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_567), .B2(n_568), .Y(n_563) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_568), .A2(n_680), .B1(n_681), .B2(n_683), .Y(n_679) );
INVx4_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_575), .B2(n_576), .Y(n_570) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g592 ( .A(n_576), .Y(n_592) );
AND4x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .C(n_581), .D(n_584), .Y(n_577) );
INVx1_ASAP7_75t_L g663 ( .A(n_585), .Y(n_663) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_624), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_605), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .C(n_597), .Y(n_589) );
BUFx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx4_ASAP7_75t_L g638 ( .A(n_604), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_604), .B(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_604), .B(n_802), .Y(n_801) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_606), .B(n_611), .C(n_616), .D(n_620), .Y(n_605) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g641 ( .A(n_610), .Y(n_641) );
INVx3_ASAP7_75t_L g727 ( .A(n_610), .Y(n_727) );
INVx2_ASAP7_75t_L g828 ( .A(n_610), .Y(n_828) );
INVx5_ASAP7_75t_L g1114 ( .A(n_610), .Y(n_1114) );
BUFx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AO22x2_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_646), .B1(n_660), .B2(n_661), .Y(n_625) );
INVx2_ASAP7_75t_L g660 ( .A(n_626), .Y(n_660) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_639), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .C(n_634), .D(n_636), .Y(n_628) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g688 ( .A(n_633), .Y(n_688) );
INVx2_ASAP7_75t_L g1097 ( .A(n_638), .Y(n_1097) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .C(n_644), .D(n_645), .Y(n_639) );
INVx1_ASAP7_75t_L g661 ( .A(n_646), .Y(n_661) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_655), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .C(n_653), .D(n_654), .Y(n_649) );
BUFx3_ASAP7_75t_L g682 ( .A(n_651), .Y(n_682) );
INVx2_ASAP7_75t_L g711 ( .A(n_651), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .C(n_658), .D(n_659), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_770), .B2(n_771), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_731), .B1(n_767), .B2(n_769), .Y(n_666) );
INVx1_ASAP7_75t_L g769 ( .A(n_667), .Y(n_769) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_696), .B1(n_728), .B2(n_729), .Y(n_667) );
INVx4_ASAP7_75t_R g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g728 ( .A(n_669), .Y(n_728) );
XNOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_670), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
AND2x4_ASAP7_75t_L g671 ( .A(n_672), .B(n_689), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_679), .C(n_684), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_678), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_677), .A2(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND4x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .C(n_692), .D(n_694), .Y(n_689) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g730 ( .A(n_698), .Y(n_730) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_719), .Y(n_701) );
NOR3xp33_ASAP7_75t_SL g702 ( .A(n_703), .B(n_709), .C(n_714), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_703) );
INVx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_718), .B(n_765), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_L g768 ( .A(n_732), .Y(n_768) );
AO22x2_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B1(n_748), .B2(n_766), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_741), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .C(n_739), .D(n_740), .Y(n_736) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .C(n_744), .D(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g766 ( .A(n_748), .Y(n_766) );
XNOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND4xp75_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .C(n_760), .D(n_763), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .Y(n_754) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_793), .B2(n_794), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
NOR4xp75_ASAP7_75t_L g777 ( .A(n_778), .B(n_781), .C(n_784), .D(n_787), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_788), .B(n_790), .Y(n_787) );
INVx2_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
OA22x2_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .B1(n_820), .B2(n_840), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x4_ASAP7_75t_L g796 ( .A(n_797), .B(n_813), .Y(n_796) );
AOI21x1_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B(n_807), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_803), .Y(n_799) );
BUFx2_ASAP7_75t_L g814 ( .A(n_800), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g818 ( .A(n_805), .B(n_811), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_806), .Y(n_819) );
INVx1_ASAP7_75t_L g817 ( .A(n_808), .Y(n_817) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
NAND4xp75_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .C(n_818), .D(n_819), .Y(n_813) );
NOR2x1_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx1_ASAP7_75t_L g840 ( .A(n_820), .Y(n_840) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
XNOR2x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
NOR2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_832), .Y(n_825) );
NAND4xp25_ASAP7_75t_L g826 ( .A(n_827), .B(n_829), .C(n_830), .D(n_831), .Y(n_826) );
NAND4xp25_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .C(n_836), .D(n_837), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_1081), .B1(n_1082), .B2(n_1101), .C(n_1106), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_987), .B(n_1035), .Y(n_842) );
OAI211xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_862), .B(n_920), .C(n_954), .Y(n_843) );
CKINVDCx14_ASAP7_75t_R g998 ( .A(n_844), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_844), .A2(n_951), .B1(n_1022), .B2(n_1024), .C(n_1031), .Y(n_1021) );
O2A1O1Ixp33_ASAP7_75t_L g1036 ( .A1(n_844), .A2(n_1037), .B(n_1040), .C(n_1044), .Y(n_1036) );
OAI222xp33_ASAP7_75t_L g1053 ( .A1(n_844), .A2(n_971), .B1(n_1006), .B2(n_1054), .C1(n_1056), .C2(n_1059), .Y(n_1053) );
INVx5_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_845), .B(n_933), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_845), .B(n_970), .Y(n_969) );
INVx3_ASAP7_75t_L g1063 ( .A(n_845), .Y(n_1063) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AND2x2_ASAP7_75t_L g921 ( .A(n_846), .B(n_922), .Y(n_921) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_846), .B(n_886), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_846), .B(n_937), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_846), .B(n_878), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_846), .B(n_879), .Y(n_1080) );
INVx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g947 ( .A(n_847), .B(n_937), .Y(n_947) );
OR2x2_ASAP7_75t_L g952 ( .A(n_847), .B(n_953), .Y(n_952) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_847), .B(n_986), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_857), .Y(n_847) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_852), .B(n_854), .Y(n_851) );
AND2x4_ASAP7_75t_L g858 ( .A(n_852), .B(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_852), .B(n_854), .Y(n_875) );
AND2x4_ASAP7_75t_L g881 ( .A(n_852), .B(n_854), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_852), .Y(n_1131) );
AND2x4_ASAP7_75t_L g855 ( .A(n_854), .B(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g889 ( .A(n_854), .B(n_856), .Y(n_889) );
AND2x2_ASAP7_75t_L g901 ( .A(n_854), .B(n_856), .Y(n_901) );
INVx2_ASAP7_75t_L g871 ( .A(n_855), .Y(n_871) );
AND2x4_ASAP7_75t_L g861 ( .A(n_856), .B(n_859), .Y(n_861) );
AND2x2_ASAP7_75t_L g885 ( .A(n_856), .B(n_859), .Y(n_885) );
AND2x2_ASAP7_75t_L g891 ( .A(n_856), .B(n_859), .Y(n_891) );
INVx3_ASAP7_75t_L g874 ( .A(n_858), .Y(n_874) );
INVx3_ASAP7_75t_L g869 ( .A(n_861), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_878), .B1(n_892), .B2(n_903), .C(n_910), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_877), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_865), .B(n_905), .Y(n_904) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_865), .B(n_929), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_865), .B(n_934), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_865), .B(n_942), .Y(n_1038) );
INVx1_ASAP7_75t_SL g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g928 ( .A(n_866), .B(n_929), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_866), .B(n_887), .Y(n_941) );
AND2x2_ASAP7_75t_L g984 ( .A(n_866), .B(n_985), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_866), .B(n_899), .Y(n_1073) );
INVx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g916 ( .A(n_867), .Y(n_916) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_867), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_867), .B(n_909), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_867), .B(n_887), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_867), .B(n_970), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_867), .B(n_879), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_867), .B(n_913), .Y(n_1065) );
OR2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_873), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_869), .A2(n_871), .B1(n_978), .B2(n_979), .Y(n_977) );
INVx1_ASAP7_75t_L g976 ( .A(n_874), .Y(n_976) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_875), .Y(n_1081) );
INVx1_ASAP7_75t_L g1029 ( .A(n_877), .Y(n_1029) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_886), .Y(n_877) );
OAI211xp5_ASAP7_75t_SL g926 ( .A1(n_878), .A2(n_927), .B(n_930), .C(n_944), .Y(n_926) );
INVx1_ASAP7_75t_L g1015 ( .A(n_878), .Y(n_1015) );
CKINVDCx6p67_ASAP7_75t_R g878 ( .A(n_879), .Y(n_878) );
AND2x2_ASAP7_75t_L g933 ( .A(n_879), .B(n_887), .Y(n_933) );
INVx1_ASAP7_75t_L g938 ( .A(n_879), .Y(n_938) );
AND2x2_ASAP7_75t_L g970 ( .A(n_879), .B(n_913), .Y(n_970) );
OR2x2_ASAP7_75t_L g986 ( .A(n_879), .B(n_887), .Y(n_986) );
OAI322xp33_ASAP7_75t_L g989 ( .A1(n_879), .A2(n_963), .A3(n_973), .B1(n_990), .B2(n_991), .C1(n_992), .C2(n_994), .Y(n_989) );
OR2x6_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .Y(n_879) );
BUFx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_887), .Y(n_913) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_887), .Y(n_1041) );
AND2x4_ASAP7_75t_L g887 ( .A(n_888), .B(n_890), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_892), .B(n_961), .Y(n_960) );
CKINVDCx16_ASAP7_75t_R g991 ( .A(n_892), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_892), .B(n_1019), .Y(n_1018) );
AND2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_897), .Y(n_892) );
AND2x2_ASAP7_75t_L g929 ( .A(n_893), .B(n_906), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_893), .B(n_909), .Y(n_935) );
OR2x2_ASAP7_75t_L g943 ( .A(n_893), .B(n_909), .Y(n_943) );
OR2x2_ASAP7_75t_L g964 ( .A(n_893), .B(n_906), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_893), .B(n_897), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_894), .Y(n_893) );
OR2x2_ASAP7_75t_L g919 ( .A(n_894), .B(n_906), .Y(n_919) );
AND2x2_ASAP7_75t_L g946 ( .A(n_894), .B(n_906), .Y(n_946) );
AND2x2_ASAP7_75t_L g894 ( .A(n_895), .B(n_896), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_897), .B(n_928), .Y(n_927) );
AND2x2_ASAP7_75t_L g945 ( .A(n_897), .B(n_946), .Y(n_945) );
AND2x2_ASAP7_75t_L g950 ( .A(n_897), .B(n_929), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_897), .B(n_967), .Y(n_1001) );
O2A1O1Ixp33_ASAP7_75t_SL g1044 ( .A1(n_897), .A2(n_1045), .B(n_1048), .C(n_1050), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_897), .B(n_1016), .Y(n_1049) );
AND3x1_ASAP7_75t_L g1055 ( .A(n_897), .B(n_922), .C(n_928), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_897), .B(n_906), .Y(n_1058) );
INVx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx3_ASAP7_75t_L g909 ( .A(n_899), .Y(n_909) );
OR2x2_ASAP7_75t_L g996 ( .A(n_899), .B(n_906), .Y(n_996) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AOI31xp33_ASAP7_75t_L g1037 ( .A1(n_904), .A2(n_1029), .A3(n_1038), .B(n_1039), .Y(n_1037) );
INVxp67_ASAP7_75t_SL g1030 ( .A(n_905), .Y(n_1030) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_909), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
OR2x2_ASAP7_75t_L g918 ( .A(n_909), .B(n_919), .Y(n_918) );
AND2x2_ASAP7_75t_L g924 ( .A(n_909), .B(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_909), .B(n_963), .Y(n_962) );
AND2x2_ASAP7_75t_L g972 ( .A(n_909), .B(n_946), .Y(n_972) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_909), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_909), .B(n_964), .Y(n_1011) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_914), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_911), .B(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g922 ( .A(n_912), .Y(n_922) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_917), .Y(n_914) );
AND2x2_ASAP7_75t_L g923 ( .A(n_915), .B(n_924), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g944 ( .A(n_915), .B(n_945), .C(n_947), .Y(n_944) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_916), .B(n_964), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_916), .B(n_996), .Y(n_995) );
O2A1O1Ixp33_ASAP7_75t_L g1031 ( .A1(n_916), .A2(n_991), .B(n_1032), .C(n_1034), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_916), .B(n_946), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_916), .B(n_972), .Y(n_1076) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g925 ( .A(n_919), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_919), .B(n_1047), .Y(n_1046) );
AOI211xp5_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_923), .B(n_926), .C(n_948), .Y(n_920) );
INVx1_ASAP7_75t_L g1034 ( .A(n_921), .Y(n_1034) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_922), .A2(n_1013), .B1(n_1014), .B2(n_1016), .C(n_1017), .Y(n_1012) );
INVx1_ASAP7_75t_L g1007 ( .A(n_924), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_927), .Y(n_997) );
AND2x2_ASAP7_75t_L g982 ( .A(n_929), .B(n_983), .Y(n_982) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_929), .B(n_1043), .Y(n_1042) );
AOI21xp33_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_934), .B(n_936), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g953 ( .A(n_933), .Y(n_953) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_935), .B(n_941), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_937), .B(n_939), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_937), .B(n_993), .Y(n_1006) );
AOI211xp5_ASAP7_75t_L g1051 ( .A1(n_937), .A2(n_1052), .B(n_1053), .C(n_1060), .Y(n_1051) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
AOI21xp33_ASAP7_75t_SL g1079 ( .A1(n_939), .A2(n_1010), .B(n_1080), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .Y(n_939) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_940), .B(n_950), .Y(n_1052) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g1068 ( .A(n_945), .Y(n_1068) );
INVx1_ASAP7_75t_L g1047 ( .A(n_946), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_947), .B(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g1059 ( .A(n_947), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_950), .B(n_985), .Y(n_1004) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
AOI211xp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_959), .B(n_965), .C(n_980), .Y(n_954) );
INVxp67_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVxp67_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
OAI21xp5_ASAP7_75t_L g981 ( .A1(n_963), .A2(n_982), .B(n_984), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_963), .B(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_968), .B1(n_971), .B2(n_973), .C(n_974), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVxp67_ASAP7_75t_SL g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g973 ( .A(n_970), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_971), .B(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
NOR3xp33_ASAP7_75t_L g1002 ( .A(n_974), .B(n_1003), .C(n_1005), .Y(n_1002) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g1039 ( .A(n_982), .Y(n_1039) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND5xp2_ASAP7_75t_SL g987 ( .A(n_988), .B(n_999), .C(n_1002), .D(n_1012), .E(n_1021), .Y(n_987) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_997), .B(n_998), .Y(n_988) );
INVx1_ASAP7_75t_L g1043 ( .A(n_990), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_1000), .Y(n_999) );
INVxp67_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1007), .B1(n_1008), .B2(n_1010), .Y(n_1005) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
CKINVDCx14_ASAP7_75t_R g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_1020), .A2(n_1061), .B(n_1066), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1027), .B1(n_1029), .B2(n_1030), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVxp67_ASAP7_75t_SL g1032 ( .A(n_1033), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1051), .C(n_1069), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1039), .B(n_1068), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_1041), .B(n_1058), .Y(n_1057) );
NOR2xp33_ASAP7_75t_L g1070 ( .A(n_1041), .B(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g1056 ( .A(n_1057), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1064), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1074), .B1(n_1075), .B2(n_1077), .C(n_1079), .Y(n_1069) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
XNOR2x1_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
NOR2x1_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1092), .Y(n_1086) );
NAND4xp25_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .C(n_1090), .D(n_1091), .Y(n_1087) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1098), .C(n_1100), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1118), .Y(n_1109) );
NOR3xp33_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1113), .C(n_1115), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1122), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1126), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
endmodule