module fake_ariane_3200_n_1432 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1432);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1432;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_186),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_2),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_142),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_40),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_137),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_255),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_14),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_244),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_104),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_56),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_133),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_65),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_39),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_113),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_16),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_125),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_230),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_126),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_159),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_210),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_236),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_83),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_175),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_7),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_4),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_228),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_114),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_88),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_18),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_238),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_43),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_20),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_270),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_202),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_220),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_178),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_91),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_239),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_257),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_48),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_89),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_140),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_0),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_34),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_165),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_13),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_112),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_20),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_102),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_106),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_10),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_90),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_19),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_43),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_222),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_163),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_219),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_17),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_96),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_82),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_119),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_232),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_116),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_152),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_240),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_78),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_190),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_91),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_109),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_100),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_87),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_283),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_33),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_121),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_169),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_243),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_208),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_273),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_188),
.Y(n_397)
);

BUFx5_ASAP7_75t_L g398 ( 
.A(n_15),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_166),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_150),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_135),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_192),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_143),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_268),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_131),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_33),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_227),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_73),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_307),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_129),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_292),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_304),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_47),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_115),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_145),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_10),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_158),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_39),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_70),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_34),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_308),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_50),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_171),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_38),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_84),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_2),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_261),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_302),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_63),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_267),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_128),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_48),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_136),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_139),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_313),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_144),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_312),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_231),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_256),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_277),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_29),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_249),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_61),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_97),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_284),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_17),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_300),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_84),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_262),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_141),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_79),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_306),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_213),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_111),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_303),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_1),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_120),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_81),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_223),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_275),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_68),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_24),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_309),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_13),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_148),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_310),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_274),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_263),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_173),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_161),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_88),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_168),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_55),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_234),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_26),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_258),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_248),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_288),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_46),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_315),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_4),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_28),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_207),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_92),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_187),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_56),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_52),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_172),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_107),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_297),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_21),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_200),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_174),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_281),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_211),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_59),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_197),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_149),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_28),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_250),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_242),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_98),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_167),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_259),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_138),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_69),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_25),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_193),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_181),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_286),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_195),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_179),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_59),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_85),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_8),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_21),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_75),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_92),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_108),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_241),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_285),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_206),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_209),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_82),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_185),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_254),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_81),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_251),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_147),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_99),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_118),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_290),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_226),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_29),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_235),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_105),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_225),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_1),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_224),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_287),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_26),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_212),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_473),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_473),
.B(n_0),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_316),
.Y(n_545)
);

BUFx8_ASAP7_75t_SL g546 ( 
.A(n_329),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_316),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_473),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_398),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_316),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_316),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_413),
.B(n_3),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_498),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_398),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_398),
.B(n_3),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_367),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_398),
.B(n_435),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_406),
.B(n_446),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_413),
.B(n_5),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_398),
.B(n_5),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_398),
.B(n_6),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_498),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_498),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_462),
.B(n_6),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_462),
.B(n_7),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_538),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_498),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_538),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_538),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_344),
.B(n_8),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_322),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_344),
.B(n_9),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_332),
.B(n_93),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_361),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_361),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_340),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_514),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_363),
.Y(n_580)
);

BUFx8_ASAP7_75t_SL g581 ( 
.A(n_329),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_322),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_337),
.B(n_9),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_432),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_363),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_341),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_535),
.B(n_11),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_324),
.B(n_11),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_322),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_407),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_357),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_416),
.B(n_12),
.Y(n_592)
);

NOR2x1_ASAP7_75t_L g593 ( 
.A(n_476),
.B(n_94),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_327),
.B(n_12),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_330),
.B(n_14),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_369),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_416),
.B(n_15),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_542),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_323),
.B(n_16),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_425),
.B(n_18),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_334),
.B(n_19),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_358),
.B(n_22),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_420),
.B(n_22),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_407),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_346),
.B(n_23),
.Y(n_608)
);

BUFx8_ASAP7_75t_SL g609 ( 
.A(n_432),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_355),
.B(n_23),
.Y(n_610)
);

BUFx12f_ASAP7_75t_L g611 ( 
.A(n_455),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_386),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_317),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_441),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_373),
.B(n_27),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_332),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_441),
.B(n_27),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_426),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_455),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_448),
.B(n_30),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_374),
.B(n_30),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_443),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_448),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_456),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_497),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_471),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_484),
.B(n_31),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_507),
.B(n_31),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_497),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_497),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_482),
.B(n_391),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_377),
.B(n_32),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_392),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_382),
.B(n_32),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_391),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_383),
.B(n_35),
.Y(n_638)
);

NOR2x1_ASAP7_75t_L g639 ( 
.A(n_397),
.B(n_95),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_392),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_404),
.B(n_35),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_391),
.B(n_36),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_409),
.B(n_36),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_516),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_423),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_423),
.B(n_101),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_328),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_524),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_517),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_333),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_518),
.B(n_405),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_524),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_505),
.B(n_379),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_405),
.B(n_434),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_524),
.B(n_37),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_379),
.B(n_37),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_399),
.B(n_38),
.Y(n_657)
);

BUFx12f_ASAP7_75t_L g658 ( 
.A(n_328),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_411),
.B(n_40),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_333),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_434),
.B(n_41),
.Y(n_661)
);

BUFx12f_ASAP7_75t_L g662 ( 
.A(n_331),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_521),
.B(n_41),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_430),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_521),
.B(n_42),
.Y(n_665)
);

BUFx8_ASAP7_75t_L g666 ( 
.A(n_430),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_414),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_417),
.B(n_42),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_494),
.B(n_44),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_428),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_431),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_335),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_494),
.B(n_44),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_527),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_520),
.B(n_45),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_436),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_527),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_534),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_534),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_445),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_520),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_532),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_447),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_449),
.B(n_46),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_319),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_450),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_459),
.B(n_463),
.Y(n_688)
);

BUFx8_ASAP7_75t_SL g689 ( 
.A(n_506),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_326),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_478),
.B(n_47),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_336),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_490),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_500),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_502),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_653),
.A2(n_509),
.B1(n_442),
.B2(n_506),
.Y(n_696)
);

AO22x2_ASAP7_75t_L g697 ( 
.A1(n_632),
.A2(n_429),
.B1(n_347),
.B2(n_385),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_653),
.A2(n_509),
.B1(n_442),
.B2(n_338),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_571),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_660),
.B(n_439),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_637),
.B(n_508),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_571),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_657),
.A2(n_348),
.B1(n_353),
.B2(n_345),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_656),
.A2(n_359),
.B1(n_360),
.B2(n_356),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_605),
.A2(n_364),
.B1(n_368),
.B2(n_362),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_605),
.A2(n_541),
.B1(n_376),
.B2(n_378),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_590),
.B(n_597),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_582),
.B(n_370),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_656),
.A2(n_389),
.B1(n_408),
.B2(n_384),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_589),
.B(n_418),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_556),
.B(n_419),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_601),
.A2(n_424),
.B1(n_451),
.B2(n_422),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_606),
.A2(n_558),
.B1(n_587),
.B2(n_583),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_583),
.A2(n_461),
.B1(n_464),
.B2(n_458),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_569),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_661),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_587),
.A2(n_479),
.B1(n_481),
.B2(n_475),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_557),
.A2(n_487),
.B1(n_491),
.B2(n_486),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_647),
.A2(n_499),
.B1(n_513),
.B2(n_496),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_661),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_677),
.A2(n_342),
.B1(n_394),
.B2(n_336),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_642),
.A2(n_530),
.B1(n_537),
.B2(n_528),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_522),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_654),
.A2(n_529),
.B1(n_531),
.B2(n_525),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_654),
.A2(n_536),
.B1(n_533),
.B2(n_51),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_637),
.B(n_528),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_655),
.A2(n_537),
.B1(n_530),
.B2(n_320),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_556),
.A2(n_321),
.B1(n_325),
.B2(n_318),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_674),
.A2(n_343),
.B1(n_349),
.B2(n_339),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_663),
.A2(n_351),
.B1(n_352),
.B2(n_350),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_570),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

AO22x2_ASAP7_75t_L g734 ( 
.A1(n_552),
.A2(n_560),
.B1(n_566),
.B2(n_565),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_548),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_545),
.Y(n_736)
);

OAI22xp33_ASAP7_75t_L g737 ( 
.A1(n_674),
.A2(n_365),
.B1(n_366),
.B2(n_354),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_545),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_573),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_611),
.B(n_49),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_577),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_663),
.A2(n_372),
.B1(n_375),
.B2(n_371),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_648),
.A2(n_381),
.B1(n_387),
.B2(n_380),
.Y(n_743)
);

OA22x2_ASAP7_75t_L g744 ( 
.A1(n_652),
.A2(n_390),
.B1(n_393),
.B2(n_388),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_690),
.A2(n_396),
.B1(n_400),
.B2(n_395),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_614),
.A2(n_402),
.B1(n_403),
.B2(n_401),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_665),
.A2(n_412),
.B1(n_415),
.B2(n_410),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_651),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_590),
.B(n_421),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_SL g750 ( 
.A(n_631),
.B(n_427),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_545),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_665),
.A2(n_437),
.B1(n_438),
.B2(n_433),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_658),
.B(n_49),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_590),
.B(n_440),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_690),
.A2(n_452),
.B1(n_453),
.B2(n_444),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_678),
.A2(n_540),
.B1(n_539),
.B2(n_526),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_669),
.A2(n_675),
.B1(n_673),
.B2(n_552),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_669),
.A2(n_523),
.B1(n_519),
.B2(n_512),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_560),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_543),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_549),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_546),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_673),
.A2(n_511),
.B1(n_510),
.B2(n_504),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_559),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_578),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_675),
.A2(n_503),
.B1(n_501),
.B2(n_495),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_586),
.Y(n_767)
);

INVx5_ASAP7_75t_L g768 ( 
.A(n_590),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_597),
.Y(n_769)
);

OA22x2_ASAP7_75t_L g770 ( 
.A1(n_613),
.A2(n_493),
.B1(n_492),
.B2(n_489),
.Y(n_770)
);

AO22x2_ASAP7_75t_L g771 ( 
.A1(n_565),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_597),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_566),
.A2(n_488),
.B1(n_485),
.B2(n_483),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_557),
.A2(n_688),
.B1(n_595),
.B2(n_610),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_SL g775 ( 
.A1(n_662),
.A2(n_480),
.B1(n_477),
.B2(n_474),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_597),
.A2(n_472),
.B1(n_470),
.B2(n_469),
.Y(n_776)
);

CKINVDCx6p67_ASAP7_75t_R g777 ( 
.A(n_607),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_619),
.B(n_54),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_591),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_454),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_651),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_679),
.A2(n_468),
.B1(n_467),
.B2(n_466),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_679),
.A2(n_465),
.B1(n_460),
.B2(n_457),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_607),
.B(n_57),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_547),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_547),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_607),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_SL g788 ( 
.A1(n_581),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_584),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_596),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_612),
.B(n_62),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_550),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_550),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_688),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_612),
.B(n_64),
.Y(n_795)
);

BUFx6f_ASAP7_75t_SL g796 ( 
.A(n_577),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_741),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_735),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_698),
.B(n_572),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_757),
.B(n_612),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_765),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_767),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_739),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_779),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_774),
.B(n_672),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_790),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_760),
.Y(n_807)
);

INVxp33_ASAP7_75t_L g808 ( 
.A(n_712),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_733),
.Y(n_809)
);

INVxp33_ASAP7_75t_L g810 ( 
.A(n_708),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_761),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_764),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_699),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_702),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_710),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_716),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_732),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_717),
.Y(n_818)
);

XNOR2x2_ASAP7_75t_L g819 ( 
.A(n_696),
.B(n_726),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_717),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_721),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_721),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_701),
.Y(n_823)
);

BUFx5_ASAP7_75t_L g824 ( 
.A(n_784),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_736),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_704),
.B(n_572),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_701),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_762),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_739),
.B(n_574),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_734),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_781),
.Y(n_832)
);

XNOR2x2_ASAP7_75t_L g833 ( 
.A(n_726),
.B(n_609),
.Y(n_833)
);

AND2x6_ASAP7_75t_L g834 ( 
.A(n_791),
.B(n_574),
.Y(n_834)
);

AND2x6_ASAP7_75t_L g835 ( 
.A(n_795),
.B(n_592),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_738),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_751),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_711),
.B(n_612),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_727),
.B(n_692),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_714),
.B(n_620),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_785),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_786),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_792),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_793),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_720),
.B(n_686),
.Y(n_845)
);

XNOR2x2_ASAP7_75t_L g846 ( 
.A(n_697),
.B(n_689),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_796),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_731),
.B(n_742),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_778),
.B(n_620),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_724),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_778),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_SL g852 ( 
.A(n_775),
.B(n_588),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_737),
.B(n_555),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_770),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_749),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_754),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_728),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_722),
.B(n_620),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_780),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_725),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_725),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_744),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_789),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_777),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_769),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_772),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_707),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_758),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_768),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_763),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_768),
.B(n_592),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_766),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_723),
.B(n_620),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_750),
.B(n_626),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_709),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_759),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_768),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_759),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_771),
.Y(n_879)
);

XNOR2xp5_ASAP7_75t_L g880 ( 
.A(n_697),
.B(n_598),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_747),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_771),
.B(n_588),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_782),
.Y(n_883)
);

INVxp33_ASAP7_75t_L g884 ( 
.A(n_715),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_805),
.A2(n_752),
.B(n_773),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_834),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_809),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_829),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_811),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_830),
.B(n_626),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_805),
.A2(n_783),
.B(n_703),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_863),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_840),
.B(n_626),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_826),
.B(n_745),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_850),
.B(n_630),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_800),
.B(n_630),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_812),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_857),
.B(n_630),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_800),
.B(n_628),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_884),
.B(n_713),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_860),
.B(n_628),
.Y(n_901)
);

OR2x2_ASAP7_75t_SL g902 ( 
.A(n_875),
.B(n_788),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_829),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_857),
.B(n_746),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_825),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_849),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_798),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_801),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_815),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_829),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_802),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_826),
.B(n_629),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_849),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_799),
.B(n_629),
.Y(n_914)
);

AND2x6_ASAP7_75t_L g915 ( 
.A(n_861),
.B(n_874),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_834),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_828),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_834),
.B(n_730),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_873),
.B(n_598),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_834),
.B(n_756),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_835),
.B(n_755),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_803),
.B(n_579),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_816),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_873),
.B(n_603),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_835),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_853),
.A2(n_544),
.B(n_595),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_817),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_848),
.A2(n_853),
.B1(n_882),
.B2(n_835),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_804),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_823),
.B(n_603),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_813),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_827),
.B(n_618),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_881),
.B(n_776),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_807),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_SL g935 ( 
.A(n_818),
.B(n_544),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_810),
.B(n_808),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_810),
.B(n_883),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_855),
.A2(n_561),
.B(n_555),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_858),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_835),
.B(n_743),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_876),
.B(n_753),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_856),
.B(n_666),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_867),
.B(n_681),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_878),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_879),
.B(n_753),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_868),
.B(n_621),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_859),
.B(n_666),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_864),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_870),
.B(n_621),
.Y(n_949)
);

AND2x2_ASAP7_75t_SL g950 ( 
.A(n_848),
.B(n_561),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_872),
.B(n_671),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_814),
.B(n_729),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_839),
.B(n_683),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_847),
.B(n_579),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_839),
.B(n_695),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_836),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_838),
.B(n_576),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_814),
.B(n_610),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_806),
.B(n_580),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_854),
.B(n_585),
.Y(n_960)
);

INVxp33_ASAP7_75t_L g961 ( 
.A(n_880),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_SL g962 ( 
.A(n_831),
.B(n_705),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_862),
.B(n_740),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_869),
.B(n_639),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_837),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_871),
.B(n_599),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_824),
.B(n_616),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_824),
.B(n_622),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_820),
.B(n_740),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_845),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_841),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_842),
.Y(n_972)
);

BUFx12f_ASAP7_75t_SL g973 ( 
.A(n_819),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_821),
.B(n_627),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_936),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_950),
.B(n_824),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_931),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_944),
.B(n_822),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_950),
.B(n_824),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_886),
.B(n_794),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_886),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_948),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_904),
.B(n_900),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_892),
.B(n_970),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_936),
.B(n_832),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_950),
.B(n_824),
.Y(n_986)
);

AND2x6_ASAP7_75t_L g987 ( 
.A(n_912),
.B(n_851),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_917),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_928),
.B(n_843),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_916),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_937),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_916),
.B(n_877),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_916),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_925),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_925),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_912),
.B(n_914),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_925),
.B(n_797),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_948),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_958),
.B(n_844),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_913),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_944),
.B(n_865),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_906),
.B(n_866),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_897),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_931),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_906),
.B(n_623),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_927),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_919),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_967),
.B(n_852),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_914),
.B(n_625),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_953),
.B(n_833),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_894),
.B(n_706),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_968),
.B(n_719),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_926),
.B(n_667),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_919),
.B(n_593),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_887),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_898),
.B(n_670),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_953),
.B(n_955),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_960),
.Y(n_1018)
);

BUFx8_ASAP7_75t_L g1019 ( 
.A(n_969),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_915),
.Y(n_1020)
);

NAND2x1p5_ASAP7_75t_L g1021 ( 
.A(n_907),
.B(n_617),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_915),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_907),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_908),
.B(n_617),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_915),
.B(n_676),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_960),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_966),
.B(n_644),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_915),
.B(n_680),
.Y(n_1028)
);

CKINVDCx16_ASAP7_75t_R g1029 ( 
.A(n_922),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_908),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_927),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_915),
.B(n_694),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_911),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_911),
.B(n_617),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_929),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_966),
.B(n_901),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_887),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_SL g1038 ( 
.A(n_891),
.B(n_885),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_927),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_909),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_909),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_974),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_955),
.B(n_615),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_901),
.B(n_899),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_927),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_SL g1046 ( 
.A(n_918),
.B(n_562),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_901),
.B(n_649),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_971),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_902),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_915),
.B(n_718),
.Y(n_1050)
);

BUFx2_ASAP7_75t_SL g1051 ( 
.A(n_988),
.Y(n_1051)
);

INVx8_ASAP7_75t_L g1052 ( 
.A(n_1022),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_1019),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_1019),
.Y(n_1054)
);

AND2x6_ASAP7_75t_L g1055 ( 
.A(n_981),
.B(n_924),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_984),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_1045),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_983),
.B(n_946),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_1036),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_1022),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1003),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_1036),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_981),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_1022),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_982),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1023),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_983),
.B(n_946),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_981),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_1042),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1030),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1033),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1035),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_1022),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_994),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_1038),
.A2(n_846),
.B1(n_973),
.B2(n_924),
.Y(n_1075)
);

NAND2x1p5_ASAP7_75t_L g1076 ( 
.A(n_1020),
.B(n_889),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_1029),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_1000),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_1020),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_SL g1080 ( 
.A(n_998),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_991),
.B(n_949),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_975),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_994),
.Y(n_1083)
);

BUFx2_ASAP7_75t_SL g1084 ( 
.A(n_998),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_978),
.Y(n_1085)
);

BUFx2_ASAP7_75t_SL g1086 ( 
.A(n_978),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_994),
.Y(n_1087)
);

CKINVDCx16_ASAP7_75t_R g1088 ( 
.A(n_1049),
.Y(n_1088)
);

BUFx24_ASAP7_75t_L g1089 ( 
.A(n_1044),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_995),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_985),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_995),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_977),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1044),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1038),
.B(n_920),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_991),
.B(n_949),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1009),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_987),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1004),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_995),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_1001),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_1027),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_L g1103 ( 
.A(n_987),
.Y(n_1103)
);

BUFx2_ASAP7_75t_SL g1104 ( 
.A(n_1001),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1017),
.B(n_951),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1015),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1043),
.B(n_899),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1045),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_SL g1109 ( 
.A(n_1047),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1007),
.B(n_951),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_1045),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1047),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_1077),
.Y(n_1113)
);

OAI21xp33_ASAP7_75t_L g1114 ( 
.A1(n_1058),
.A2(n_1008),
.B(n_604),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_1053),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1051),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1110),
.A2(n_1007),
.B1(n_1008),
.B2(n_1012),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1054),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1061),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1091),
.A2(n_996),
.B1(n_980),
.B2(n_1011),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1075),
.A2(n_902),
.B1(n_1011),
.B2(n_1010),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1067),
.A2(n_1012),
.B1(n_979),
.B2(n_986),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_1080),
.Y(n_1123)
);

INVx8_ASAP7_75t_L g1124 ( 
.A(n_1055),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1066),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1080),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_1082),
.Y(n_1127)
);

BUFx8_ASAP7_75t_SL g1128 ( 
.A(n_1065),
.Y(n_1128)
);

BUFx8_ASAP7_75t_L g1129 ( 
.A(n_1054),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1075),
.A2(n_973),
.B1(n_996),
.B2(n_961),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1052),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1091),
.A2(n_996),
.B1(n_1097),
.B2(n_939),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1070),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1059),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1071),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1072),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1078),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_1065),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1093),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1108),
.Y(n_1140)
);

BUFx2_ASAP7_75t_R g1141 ( 
.A(n_1104),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1099),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1105),
.A2(n_1037),
.B1(n_1041),
.B2(n_1040),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1106),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1056),
.Y(n_1145)
);

INVx6_ASAP7_75t_L g1146 ( 
.A(n_1101),
.Y(n_1146)
);

CKINVDCx8_ASAP7_75t_R g1147 ( 
.A(n_1086),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1081),
.A2(n_980),
.B1(n_1050),
.B2(n_1016),
.Y(n_1148)
);

INVx6_ASAP7_75t_L g1149 ( 
.A(n_1101),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1093),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1095),
.B(n_976),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1107),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1096),
.A2(n_1050),
.B1(n_934),
.B2(n_987),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1103),
.A2(n_979),
.B1(n_986),
.B2(n_976),
.Y(n_1154)
);

CKINVDCx11_ASAP7_75t_R g1155 ( 
.A(n_1101),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1078),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1085),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1095),
.A2(n_787),
.B(n_604),
.Y(n_1158)
);

BUFx8_ASAP7_75t_L g1159 ( 
.A(n_1069),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1103),
.A2(n_929),
.B1(n_1013),
.B2(n_1016),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1084),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1098),
.A2(n_934),
.B1(n_987),
.B2(n_1014),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1062),
.Y(n_1163)
);

CKINVDCx8_ASAP7_75t_R g1164 ( 
.A(n_1088),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1098),
.A2(n_1014),
.B1(n_923),
.B2(n_933),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1094),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1109),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1102),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1094),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1089),
.A2(n_1013),
.B1(n_938),
.B2(n_999),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1069),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1112),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1109),
.Y(n_1173)
);

BUFx4f_ASAP7_75t_SL g1174 ( 
.A(n_1108),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1055),
.A2(n_1018),
.B1(n_1026),
.B2(n_1014),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1057),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1055),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1052),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1120),
.A2(n_1158),
.B1(n_1121),
.B2(n_1153),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1170),
.A2(n_962),
.B1(n_921),
.B2(n_940),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1130),
.A2(n_1014),
.B1(n_947),
.B2(n_942),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1170),
.A2(n_954),
.B1(n_1089),
.B2(n_1046),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1119),
.B(n_1057),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1151),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1148),
.A2(n_923),
.B1(n_893),
.B2(n_956),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1139),
.Y(n_1186)
);

OAI222xp33_ASAP7_75t_L g1187 ( 
.A1(n_1165),
.A2(n_1032),
.B1(n_1028),
.B2(n_1025),
.C1(n_952),
.C2(n_972),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1156),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_SL g1189 ( 
.A(n_1118),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1117),
.B(n_1079),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1153),
.A2(n_1117),
.B1(n_1161),
.B2(n_1152),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1132),
.A2(n_1005),
.B1(n_974),
.B2(n_957),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1113),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1160),
.A2(n_1032),
.B1(n_895),
.B2(n_999),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1125),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1146),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1133),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1135),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1122),
.A2(n_965),
.B1(n_972),
.B2(n_971),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1159),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1124),
.A2(n_945),
.B1(n_941),
.B2(n_963),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1114),
.A2(n_608),
.B(n_594),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1128),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1136),
.Y(n_1204)
);

BUFx4f_ASAP7_75t_SL g1205 ( 
.A(n_1129),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1162),
.A2(n_965),
.B1(n_971),
.B2(n_1055),
.Y(n_1206)
);

AND2x2_ASAP7_75t_SL g1207 ( 
.A(n_1162),
.B(n_1060),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1172),
.A2(n_971),
.B1(n_1055),
.B2(n_959),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1164),
.A2(n_969),
.B1(n_945),
.B2(n_941),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1142),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1157),
.B(n_888),
.Y(n_1211)
);

OAI222xp33_ASAP7_75t_L g1212 ( 
.A1(n_1145),
.A2(n_989),
.B1(n_643),
.B2(n_684),
.C1(n_668),
.C2(n_636),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1145),
.A2(n_905),
.B1(n_945),
.B2(n_941),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1144),
.Y(n_1214)
);

AOI222xp33_ASAP7_75t_L g1215 ( 
.A1(n_1175),
.A2(n_641),
.B1(n_691),
.B2(n_659),
.C1(n_638),
.C2(n_963),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1124),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1154),
.A2(n_905),
.B1(n_896),
.B2(n_963),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1143),
.A2(n_905),
.B1(n_896),
.B2(n_943),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1151),
.A2(n_935),
.B(n_641),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1150),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1137),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1166),
.A2(n_602),
.B1(n_1002),
.B2(n_659),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1176),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1127),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1169),
.B(n_1111),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1141),
.B(n_903),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1155),
.A2(n_910),
.B1(n_1002),
.B2(n_691),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1168),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1171),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1116),
.A2(n_638),
.B1(n_932),
.B2(n_930),
.Y(n_1230)
);

OAI222xp33_ASAP7_75t_L g1231 ( 
.A1(n_1147),
.A2(n_684),
.B1(n_668),
.B2(n_643),
.C1(n_636),
.C2(n_633),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1177),
.A2(n_600),
.B1(n_932),
.B2(n_930),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1138),
.Y(n_1233)
);

OAI222xp33_ASAP7_75t_L g1234 ( 
.A1(n_1179),
.A2(n_964),
.B1(n_1034),
.B2(n_1024),
.C1(n_1021),
.C2(n_562),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1181),
.A2(n_693),
.B1(n_687),
.B2(n_615),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1207),
.A2(n_1146),
.B1(n_1149),
.B2(n_1134),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1184),
.B(n_1134),
.Y(n_1237)
);

OAI221xp5_ASAP7_75t_L g1238 ( 
.A1(n_1202),
.A2(n_634),
.B1(n_964),
.B2(n_1167),
.C(n_1173),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1207),
.A2(n_1146),
.B1(n_1149),
.B2(n_1134),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1182),
.A2(n_1126),
.B1(n_1174),
.B2(n_1149),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1215),
.A2(n_693),
.B1(n_687),
.B2(n_624),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1183),
.B(n_1163),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1180),
.A2(n_1163),
.B1(n_1115),
.B2(n_1159),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1191),
.A2(n_1163),
.B1(n_693),
.B2(n_687),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1196),
.B(n_1174),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1211),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1230),
.A2(n_1131),
.B1(n_1006),
.B2(n_1076),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1192),
.A2(n_640),
.B1(n_645),
.B2(n_664),
.Y(n_1248)
);

AOI222xp33_ASAP7_75t_L g1249 ( 
.A1(n_1212),
.A2(n_575),
.B1(n_646),
.B2(n_635),
.C1(n_682),
.C2(n_890),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1195),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1194),
.A2(n_1123),
.B1(n_1060),
.B2(n_1064),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1183),
.B(n_1140),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1185),
.A2(n_682),
.B1(n_1039),
.B2(n_1031),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1209),
.A2(n_997),
.B1(n_1073),
.B2(n_1039),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1217),
.A2(n_997),
.B1(n_1178),
.B2(n_1079),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1226),
.A2(n_1064),
.B1(n_1060),
.B2(n_1048),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1227),
.A2(n_1199),
.B1(n_1206),
.B2(n_1232),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1229),
.A2(n_1073),
.B1(n_575),
.B2(n_646),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1197),
.B(n_1108),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1224),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1196),
.B(n_1140),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1201),
.A2(n_1063),
.B1(n_1100),
.B2(n_1068),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1190),
.A2(n_1074),
.B1(n_1083),
.B2(n_1064),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1218),
.A2(n_646),
.B1(n_575),
.B2(n_1074),
.Y(n_1264)
);

NAND4xp25_ASAP7_75t_L g1265 ( 
.A(n_1219),
.B(n_66),
.C(n_67),
.D(n_68),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1220),
.A2(n_685),
.B1(n_681),
.B2(n_890),
.Y(n_1266)
);

OAI211xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1188),
.A2(n_67),
.B(n_69),
.C(n_70),
.Y(n_1267)
);

AOI222xp33_ASAP7_75t_L g1268 ( 
.A1(n_1231),
.A2(n_681),
.B1(n_685),
.B2(n_73),
.C1(n_74),
.C2(n_76),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1213),
.A2(n_685),
.B1(n_1092),
.B2(n_1090),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1208),
.A2(n_1083),
.B1(n_1111),
.B2(n_1090),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1225),
.B(n_71),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1210),
.A2(n_1092),
.B1(n_1090),
.B2(n_1087),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1222),
.B(n_1090),
.C(n_1087),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1187),
.A2(n_71),
.B(n_72),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1221),
.A2(n_1092),
.B1(n_1087),
.B2(n_993),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1214),
.A2(n_1092),
.B1(n_1087),
.B2(n_993),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1228),
.A2(n_990),
.B1(n_992),
.B2(n_564),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1220),
.A2(n_551),
.B(n_550),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1198),
.A2(n_1204),
.B1(n_1233),
.B2(n_1200),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1200),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1233),
.A2(n_551),
.B1(n_563),
.B2(n_564),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1242),
.B(n_1246),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1252),
.B(n_1223),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1251),
.B(n_1236),
.Y(n_1284)
);

NAND4xp25_ASAP7_75t_L g1285 ( 
.A(n_1265),
.B(n_1268),
.C(n_1267),
.D(n_1274),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1250),
.B(n_1186),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1260),
.B(n_79),
.Y(n_1287)
);

NAND4xp25_ASAP7_75t_L g1288 ( 
.A(n_1280),
.B(n_1279),
.C(n_1241),
.D(n_1238),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1239),
.B(n_1216),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1260),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1257),
.A2(n_1193),
.B1(n_1205),
.B2(n_1189),
.Y(n_1291)
);

AND2x2_ASAP7_75t_SL g1292 ( 
.A(n_1244),
.B(n_1203),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1271),
.B(n_80),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1237),
.B(n_85),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1259),
.B(n_1272),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1272),
.B(n_86),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1276),
.B(n_90),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1243),
.B(n_103),
.Y(n_1298)
);

NAND2x1_ASAP7_75t_L g1299 ( 
.A(n_1263),
.B(n_551),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1240),
.A2(n_564),
.B(n_563),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1261),
.B(n_1247),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1278),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1234),
.A2(n_553),
.B(n_568),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1245),
.B(n_110),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_568),
.C(n_553),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1275),
.B(n_117),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1277),
.A2(n_122),
.B(n_123),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1254),
.B(n_124),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1270),
.A2(n_568),
.B1(n_553),
.B2(n_132),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1255),
.B(n_314),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1256),
.B(n_127),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1290),
.B(n_1278),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1291),
.B(n_1292),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1285),
.A2(n_1235),
.B1(n_1248),
.B2(n_1249),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1302),
.A2(n_1278),
.B(n_1262),
.Y(n_1315)
);

NOR2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1288),
.B(n_1281),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1286),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1290),
.B(n_1277),
.Y(n_1318)
);

NAND4xp75_ASAP7_75t_L g1319 ( 
.A(n_1284),
.B(n_1292),
.C(n_1289),
.D(n_1297),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1283),
.B(n_1281),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1282),
.B(n_1253),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1295),
.B(n_1269),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1301),
.B(n_1266),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1308),
.A2(n_1264),
.B1(n_1258),
.B2(n_134),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1287),
.B(n_130),
.Y(n_1325)
);

AO21x2_ASAP7_75t_L g1326 ( 
.A1(n_1296),
.A2(n_146),
.B(n_151),
.Y(n_1326)
);

NAND4xp75_ASAP7_75t_L g1327 ( 
.A(n_1289),
.B(n_153),
.C(n_154),
.D(n_155),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1310),
.A2(n_156),
.B(n_157),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1293),
.A2(n_160),
.B1(n_162),
.B2(n_164),
.C(n_170),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1308),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1294),
.B(n_182),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1317),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1317),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1313),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1318),
.B(n_1308),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1312),
.Y(n_1336)
);

AO22x2_ASAP7_75t_L g1337 ( 
.A1(n_1319),
.A2(n_1300),
.B1(n_1303),
.B2(n_1298),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_SL g1338 ( 
.A(n_1316),
.B(n_1306),
.Y(n_1338)
);

XNOR2x2_ASAP7_75t_SL g1339 ( 
.A(n_1319),
.B(n_1305),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1312),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1326),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1322),
.B(n_1299),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1322),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1320),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1315),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1315),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1321),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1343),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1347),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1338),
.A2(n_1328),
.B1(n_1323),
.B2(n_1326),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1343),
.Y(n_1351)
);

AO22x2_ASAP7_75t_L g1352 ( 
.A1(n_1344),
.A2(n_1323),
.B1(n_1331),
.B2(n_1327),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1334),
.B(n_1325),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1342),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1334),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1336),
.Y(n_1356)
);

OA22x2_ASAP7_75t_L g1357 ( 
.A1(n_1335),
.A2(n_1330),
.B1(n_1311),
.B2(n_1304),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1345),
.Y(n_1358)
);

AOI22x1_ASAP7_75t_L g1359 ( 
.A1(n_1352),
.A2(n_1337),
.B1(n_1340),
.B2(n_1341),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1349),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1354),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1351),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1350),
.A2(n_1336),
.B1(n_1314),
.B2(n_1339),
.Y(n_1363)
);

AO22x2_ASAP7_75t_L g1364 ( 
.A1(n_1355),
.A2(n_1346),
.B1(n_1333),
.B2(n_1332),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1356),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1358),
.Y(n_1366)
);

AO22x1_ASAP7_75t_L g1367 ( 
.A1(n_1353),
.A2(n_1336),
.B1(n_1346),
.B2(n_1326),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1357),
.A2(n_1324),
.B1(n_1329),
.B2(n_1307),
.Y(n_1368)
);

AO22x1_ASAP7_75t_L g1369 ( 
.A1(n_1348),
.A2(n_1328),
.B1(n_1315),
.B2(n_1309),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1360),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1359),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1362),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1366),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1361),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1373),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1370),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1371),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1371),
.B(n_1365),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1370),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1376),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1377),
.A2(n_1363),
.B(n_1368),
.C(n_1372),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1379),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1375),
.Y(n_1383)
);

NAND4xp25_ASAP7_75t_SL g1384 ( 
.A(n_1378),
.B(n_1374),
.C(n_1369),
.D(n_1367),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1384),
.A2(n_1364),
.B1(n_184),
.B2(n_189),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1383),
.B(n_183),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1380),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1381),
.A2(n_191),
.B1(n_194),
.B2(n_196),
.Y(n_1388)
);

AO22x1_ASAP7_75t_L g1389 ( 
.A1(n_1382),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_1389)
);

OAI22x1_ASAP7_75t_L g1390 ( 
.A1(n_1385),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1387),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1386),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1388),
.Y(n_1393)
);

AND4x1_ASAP7_75t_L g1394 ( 
.A(n_1391),
.B(n_1389),
.C(n_215),
.D(n_216),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1392),
.B(n_214),
.Y(n_1395)
);

AO22x2_ASAP7_75t_L g1396 ( 
.A1(n_1393),
.A2(n_217),
.B1(n_218),
.B2(n_221),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1390),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1391),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1395),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1398),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1397),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1396),
.B(n_233),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1396),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1394),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1397),
.A2(n_237),
.B1(n_245),
.B2(n_246),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1395),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1399),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1401),
.Y(n_1408)
);

OA22x2_ASAP7_75t_L g1409 ( 
.A1(n_1404),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1406),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1400),
.A2(n_266),
.B1(n_269),
.B2(n_271),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1403),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1402),
.Y(n_1413)
);

OAI22x1_ASAP7_75t_L g1414 ( 
.A1(n_1405),
.A2(n_272),
.B1(n_276),
.B2(n_278),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1408),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1410),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1409),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1413),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1414),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1412),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1411),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1407),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1418),
.A2(n_1420),
.B1(n_1416),
.B2(n_1417),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1419),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1423),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1424),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1425),
.A2(n_1415),
.B1(n_1421),
.B2(n_1422),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1426),
.A2(n_289),
.B1(n_293),
.B2(n_294),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1427),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1428),
.Y(n_1430)
);

AOI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1429),
.A2(n_295),
.B1(n_296),
.B2(n_298),
.C(n_299),
.Y(n_1431)
);

AOI211xp5_ASAP7_75t_L g1432 ( 
.A1(n_1431),
.A2(n_1430),
.B(n_305),
.C(n_311),
.Y(n_1432)
);


endmodule