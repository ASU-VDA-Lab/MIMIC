module fake_jpeg_2998_n_593 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_593);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_593;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_58),
.B(n_62),
.Y(n_135)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g208 ( 
.A(n_61),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_65),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_68),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_67),
.B(n_71),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_14),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_25),
.B(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_77),
.B(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_81),
.Y(n_161)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_103),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_33),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

CKINVDCx6p67_ASAP7_75t_R g168 ( 
.A(n_105),
.Y(n_168)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_114),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_55),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_40),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_42),
.Y(n_155)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_125),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_26),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_121),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_0),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_42),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_58),
.B(n_66),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_138),
.B(n_184),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_20),
.B(n_52),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_140),
.B(n_173),
.Y(n_288)
);

BUFx2_ASAP7_75t_SL g148 ( 
.A(n_105),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_148),
.Y(n_220)
);

HAxp5_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_55),
.CON(n_152),
.SN(n_152)
);

NAND2x1_ASAP7_75t_SL g247 ( 
.A(n_152),
.B(n_218),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_159),
.B(n_202),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_165),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_60),
.A2(n_108),
.B1(n_79),
.B2(n_90),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_169),
.A2(n_181),
.B1(n_134),
.B2(n_206),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_52),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_54),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_54),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_187),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_69),
.A2(n_22),
.B1(n_36),
.B2(n_39),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_61),
.A2(n_22),
.B1(n_36),
.B2(n_39),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g272 ( 
.A1(n_182),
.A2(n_195),
.B1(n_209),
.B2(n_157),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_65),
.A2(n_43),
.B(n_23),
.C(n_30),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_124),
.B(n_43),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_61),
.B(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_189),
.B(n_192),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_100),
.B(n_23),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_100),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_194),
.B(n_200),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_98),
.A2(n_39),
.B1(n_36),
.B2(n_22),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_87),
.B(n_1),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_91),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_89),
.B(n_1),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_80),
.C(n_112),
.Y(n_225)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_109),
.A2(n_34),
.B1(n_29),
.B2(n_41),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_75),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_12),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_93),
.B(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_217),
.B(n_208),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_73),
.B(n_41),
.Y(n_218)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_223),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_225),
.A2(n_278),
.B(n_279),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_144),
.A2(n_106),
.B1(n_97),
.B2(n_34),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_226),
.A2(n_230),
.B1(n_231),
.B2(n_282),
.Y(n_318)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_163),
.Y(n_227)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_143),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_234),
.A2(n_240),
.B1(n_243),
.B2(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_235),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_133),
.B(n_5),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_236),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_237),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_238),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_167),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_181),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_249),
.B1(n_252),
.B2(n_292),
.Y(n_303)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_152),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_204),
.B(n_151),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_246),
.B(n_260),
.C(n_295),
.Y(n_324)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_135),
.A2(n_218),
.B1(n_154),
.B2(n_130),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_147),
.A2(n_190),
.B1(n_182),
.B2(n_156),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_161),
.Y(n_251)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_211),
.A2(n_214),
.B1(n_195),
.B2(n_186),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_161),
.Y(n_253)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_146),
.Y(n_254)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx4_ASAP7_75t_SL g255 ( 
.A(n_168),
.Y(n_255)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_175),
.Y(n_257)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_170),
.Y(n_258)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_153),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_259),
.B(n_268),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_129),
.B(n_162),
.C(n_160),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_134),
.Y(n_261)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_136),
.Y(n_262)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_131),
.B(n_168),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_265),
.B(n_270),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_128),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_267),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_168),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_142),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_272),
.A2(n_280),
.B1(n_281),
.B2(n_255),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_188),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_276),
.Y(n_297)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_274),
.Y(n_350)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_275),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_164),
.B(n_201),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_191),
.A2(n_214),
.B1(n_211),
.B2(n_215),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_137),
.A2(n_145),
.B1(n_199),
.B2(n_185),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_193),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_188),
.B(n_132),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_287),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_137),
.Y(n_285)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_193),
.Y(n_286)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_198),
.B(n_145),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_247),
.Y(n_326)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_206),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_291),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_158),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_290),
.Y(n_321)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_166),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_166),
.A2(n_158),
.B1(n_199),
.B2(n_185),
.Y(n_292)
);

CKINVDCx12_ASAP7_75t_R g293 ( 
.A(n_174),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_293),
.Y(n_332)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_294),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_173),
.B(n_157),
.C(n_179),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_228),
.B(n_141),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_299),
.B(n_300),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_141),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_179),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_312),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_247),
.A2(n_174),
.B(n_179),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_310),
.A2(n_349),
.B(n_264),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_219),
.B(n_174),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_231),
.A2(n_205),
.B1(n_175),
.B2(n_170),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_319),
.A2(n_325),
.B1(n_333),
.B2(n_346),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_277),
.A2(n_234),
.B1(n_269),
.B2(n_281),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_326),
.B(n_318),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_233),
.A2(n_250),
.B1(n_243),
.B2(n_252),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_266),
.B(n_236),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_221),
.C(n_276),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_339),
.A2(n_351),
.B1(n_271),
.B2(n_239),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_229),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_264),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_272),
.A2(n_241),
.B1(n_292),
.B2(n_262),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_272),
.A2(n_274),
.B(n_220),
.C(n_271),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_224),
.A2(n_240),
.B1(n_290),
.B2(n_237),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_SL g397 ( 
.A1(n_352),
.A2(n_371),
.B(n_390),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_224),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_354),
.B(n_355),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_220),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_223),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_367),
.Y(n_395)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_303),
.A2(n_285),
.B1(n_232),
.B2(n_238),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_359),
.A2(n_360),
.B1(n_377),
.B2(n_383),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_303),
.A2(n_222),
.B1(n_227),
.B2(n_248),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_299),
.B(n_222),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_368),
.Y(n_409)
);

INVx13_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_362),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_363),
.Y(n_422)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_326),
.A2(n_221),
.B(n_276),
.C(n_258),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_221),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_375),
.Y(n_402)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_386),
.Y(n_412)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_389),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_300),
.A2(n_257),
.B1(n_275),
.B2(n_346),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_379),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_310),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_317),
.B(n_305),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_382),
.Y(n_418)
);

INVx2_ASAP7_75t_R g381 ( 
.A(n_296),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_394),
.B(n_322),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_337),
.B(n_335),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_307),
.A2(n_306),
.B1(n_312),
.B2(n_325),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_302),
.B(n_332),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_384),
.B(n_385),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_336),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_324),
.B(n_336),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_324),
.B(n_347),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_392),
.Y(n_414)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_388),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_343),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_391),
.Y(n_416)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

NOR2x1p5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_343),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_309),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_319),
.A2(n_321),
.B1(n_330),
.B2(n_301),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_331),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_399),
.B(n_404),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_393),
.B(n_368),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_405),
.B(n_379),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_331),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_393),
.A2(n_322),
.B(n_338),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_345),
.C(n_311),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_407),
.B(n_411),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_311),
.C(n_313),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_366),
.A2(n_341),
.B1(n_327),
.B2(n_329),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_413),
.A2(n_373),
.B1(n_372),
.B2(n_364),
.Y(n_452)
);

AO21x2_ASAP7_75t_SL g415 ( 
.A1(n_377),
.A2(n_330),
.B(n_338),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_313),
.C(n_323),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_417),
.B(n_404),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_419),
.A2(n_381),
.B(n_374),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_426),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_366),
.A2(n_341),
.B1(n_329),
.B2(n_327),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_424),
.A2(n_378),
.B1(n_391),
.B2(n_375),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_298),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_418),
.B(n_395),
.Y(n_430)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_430),
.B(n_434),
.C(n_443),
.Y(n_472)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_427),
.Y(n_433)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_423),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_427),
.Y(n_435)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_435),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_436),
.B(n_414),
.Y(n_474)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_429),
.Y(n_437)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_437),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_420),
.A2(n_353),
.B1(n_383),
.B2(n_365),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_441),
.A2(n_455),
.B1(n_413),
.B2(n_416),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_450),
.B(n_461),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_402),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_414),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_445),
.B(n_459),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_400),
.B(n_357),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_446),
.B(n_449),
.Y(n_473)
);

CKINVDCx12_ASAP7_75t_R g447 ( 
.A(n_415),
.Y(n_447)
);

BUFx5_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

AO22x1_ASAP7_75t_SL g448 ( 
.A1(n_415),
.A2(n_359),
.B1(n_360),
.B2(n_358),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_451),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_400),
.B(n_367),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_454),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_420),
.A2(n_381),
.B1(n_382),
.B2(n_392),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_403),
.B1(n_409),
.B2(n_405),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g454 ( 
.A(n_410),
.B(n_362),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_425),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_457),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_426),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_309),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_458),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_408),
.B(n_323),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_445),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_409),
.A2(n_370),
.B(n_362),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_412),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_463),
.B(n_467),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_398),
.C(n_439),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_468),
.C(n_477),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_398),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_475),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_412),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_399),
.C(n_407),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_453),
.Y(n_471)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_471),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_411),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_476),
.A2(n_457),
.B1(n_440),
.B2(n_431),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_417),
.C(n_406),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_421),
.B1(n_415),
.B2(n_424),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_478),
.A2(n_488),
.B1(n_433),
.B2(n_451),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_396),
.Y(n_480)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_397),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_490),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_492),
.A2(n_503),
.B1(n_506),
.B2(n_511),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_431),
.Y(n_493)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_493),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_471),
.A2(n_469),
.B1(n_470),
.B2(n_489),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_469),
.A2(n_440),
.B1(n_447),
.B2(n_452),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_490),
.Y(n_499)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_499),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_SL g501 ( 
.A(n_473),
.B(n_454),
.C(n_435),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_501),
.B(n_505),
.Y(n_531)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_481),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_502),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_481),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_473),
.A2(n_419),
.B1(n_455),
.B2(n_444),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_482),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_509),
.Y(n_533)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_484),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_510),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_476),
.A2(n_478),
.B1(n_464),
.B2(n_485),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_460),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_512),
.Y(n_530)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_514),
.Y(n_523)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_485),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_475),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_516),
.B(n_520),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_465),
.C(n_477),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_519),
.B(n_521),
.C(n_529),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_468),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_466),
.C(n_474),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_507),
.A2(n_470),
.B(n_486),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_528),
.C(n_502),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_497),
.B(n_487),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_461),
.C(n_486),
.Y(n_529)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_534),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_532),
.B(n_500),
.Y(n_535)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

XOR2x2_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_496),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_538),
.Y(n_559)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_537),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_532),
.B(n_493),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_539),
.B(n_540),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_531),
.A2(n_492),
.B1(n_488),
.B2(n_504),
.Y(n_540)
);

AOI322xp5_ASAP7_75t_SL g542 ( 
.A1(n_533),
.A2(n_472),
.A3(n_501),
.B1(n_396),
.B2(n_512),
.C1(n_483),
.C2(n_416),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_542),
.B(n_513),
.Y(n_550)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_543),
.A2(n_544),
.B1(n_510),
.B2(n_479),
.Y(n_557)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_524),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_524),
.A2(n_494),
.B(n_499),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_546),
.A2(n_530),
.B(n_518),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_525),
.B(n_494),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_548),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_498),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_550),
.A2(n_556),
.B(n_554),
.Y(n_562)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_551),
.Y(n_565)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_545),
.Y(n_552)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_552),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_543),
.A2(n_530),
.B1(n_517),
.B2(n_514),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_553),
.A2(n_558),
.B1(n_538),
.B2(n_548),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_539),
.A2(n_547),
.B(n_546),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_535),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_544),
.A2(n_462),
.B1(n_529),
.B2(n_448),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_562),
.B(n_564),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_566),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_536),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_537),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_569),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_545),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_556),
.A2(n_551),
.B(n_559),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_570),
.A2(n_561),
.B1(n_559),
.B2(n_558),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_555),
.B(n_541),
.C(n_516),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_552),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_541),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_572),
.B(n_575),
.C(n_578),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_573),
.A2(n_549),
.B(n_520),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_570),
.B(n_519),
.Y(n_578)
);

AOI322xp5_ASAP7_75t_L g579 ( 
.A1(n_574),
.A2(n_565),
.A3(n_567),
.B1(n_563),
.B2(n_564),
.C1(n_549),
.C2(n_557),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_579),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_580),
.A2(n_581),
.B(n_583),
.Y(n_585)
);

AOI221xp5_ASAP7_75t_L g581 ( 
.A1(n_575),
.A2(n_462),
.B1(n_456),
.B2(n_450),
.C(n_429),
.Y(n_581)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_577),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_582),
.A2(n_576),
.B(n_437),
.Y(n_586)
);

AOI31xp33_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_579),
.A3(n_401),
.B(n_422),
.Y(n_587)
);

BUFx24_ASAP7_75t_SL g589 ( 
.A(n_587),
.Y(n_589)
);

A2O1A1Ixp33_ASAP7_75t_SL g588 ( 
.A1(n_585),
.A2(n_448),
.B(n_401),
.C(n_422),
.Y(n_588)
);

AOI31xp33_ASAP7_75t_L g590 ( 
.A1(n_589),
.A2(n_584),
.A3(n_588),
.B(n_298),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_590),
.B(n_363),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_363),
.C(n_388),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_592),
.B(n_388),
.Y(n_593)
);


endmodule