module fake_netlist_6_4471_n_1934 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1934);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1934;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_166;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_55),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_76),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_30),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_51),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_20),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_2),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_45),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_29),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_21),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_37),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_41),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_37),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_137),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_90),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_12),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_24),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_66),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_74),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_58),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_12),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_10),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_44),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_10),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_48),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_89),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_14),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_46),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_6),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_102),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_39),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_81),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_97),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_36),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_117),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_144),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_108),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_59),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_73),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_19),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_92),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_42),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_22),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_114),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_25),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_101),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_57),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_31),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_27),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_62),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_70),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_28),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_26),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_125),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_78),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_155),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_110),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_23),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_32),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_69),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_42),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_146),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_79),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_4),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_94),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_95),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_133),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_29),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_126),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_145),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_104),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_71),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_17),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_6),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_103),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_50),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_138),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_75),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_25),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_129),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_40),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_82),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_47),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_24),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_154),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_109),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_139),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_113),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_49),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_54),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_53),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_41),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_118),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_26),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_136),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_61),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_93),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_16),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_112),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_17),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_123),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_63),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_14),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_152),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_8),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_96),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_167),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_167),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_176),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_181),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_162),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_167),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_167),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_167),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_167),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_166),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_159),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_169),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_195),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_218),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_218),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_200),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_218),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_180),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_203),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_220),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_218),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_189),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_311),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_190),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_218),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_222),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_159),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_222),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_241),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_163),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_173),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_178),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_224),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_198),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_179),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_179),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_250),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_210),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_232),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_234),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_237),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_303),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_206),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_260),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_193),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_193),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_242),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_263),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_206),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_213),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_267),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_206),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_206),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_286),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_206),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_196),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_201),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_201),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_216),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_228),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_217),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_228),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_279),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_279),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_319),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_254),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_315),
.A2(n_255),
.B(n_225),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_326),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_328),
.B(n_225),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_292),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_254),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_338),
.Y(n_403)
);

BUFx8_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_320),
.A2(n_280),
.B(n_255),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_321),
.B(n_170),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_324),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_346),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_329),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_371),
.A2(n_280),
.B(n_160),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_332),
.B(n_158),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_305),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

AND3x2_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_168),
.C(n_161),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_316),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_381),
.Y(n_435)
);

NAND2x1p5_ASAP7_75t_L g436 ( 
.A(n_339),
.B(n_233),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_339),
.B(n_171),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_343),
.B(n_172),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_365),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_365),
.B(n_174),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_381),
.B(n_196),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_376),
.B(n_175),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_177),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_327),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_185),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_345),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_353),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_344),
.A2(n_188),
.B(n_187),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_436),
.B(n_328),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_356),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_396),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_399),
.B(n_336),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_399),
.B(n_340),
.Y(n_471)
);

OAI21xp33_ASAP7_75t_SL g472 ( 
.A1(n_399),
.A2(n_359),
.B(n_337),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_342),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_436),
.B(n_361),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_401),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_R g480 ( 
.A(n_418),
.B(n_358),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_426),
.B(n_220),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_420),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_394),
.B(n_361),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_408),
.B(n_369),
.Y(n_487)
);

NOR2x1p5_ASAP7_75t_L g488 ( 
.A(n_391),
.B(n_331),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_448),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_454),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_426),
.B(n_364),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_401),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_426),
.B(n_364),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_426),
.B(n_220),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_433),
.B(n_355),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_418),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_457),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_390),
.B(n_357),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_437),
.B(n_220),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_437),
.B(n_360),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_457),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_446),
.A2(n_305),
.B1(n_341),
.B2(n_183),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_457),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_390),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_416),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_406),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_429),
.B(n_394),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_409),
.B(n_372),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_410),
.B(n_419),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_419),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_402),
.B(n_349),
.Y(n_526)
);

BUFx6f_ASAP7_75t_SL g527 ( 
.A(n_437),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_425),
.A2(n_197),
.B(n_192),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_452),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_415),
.B(n_385),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_450),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_429),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_402),
.B(n_387),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_431),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_421),
.B(n_424),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_424),
.B(n_318),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_417),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_435),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_423),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_435),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_437),
.B(n_205),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_432),
.B(n_223),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_432),
.A2(n_434),
.B(n_443),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_434),
.B(n_438),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_423),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_438),
.B(n_226),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_442),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_438),
.B(n_215),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_438),
.B(n_231),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_439),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_443),
.B(n_229),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_443),
.B(n_230),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_403),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_422),
.Y(n_567)
);

OA22x2_ASAP7_75t_L g568 ( 
.A1(n_444),
.A2(n_389),
.B1(n_388),
.B2(n_386),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_443),
.B(n_447),
.Y(n_570)
);

BUFx6f_ASAP7_75t_SL g571 ( 
.A(n_447),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_456),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_422),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_411),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_411),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_422),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_404),
.B(n_350),
.C(n_325),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_456),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_444),
.B(n_354),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_440),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_447),
.B(n_239),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_456),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_411),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_411),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_447),
.B(n_244),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_404),
.B(n_350),
.C(n_186),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_404),
.A2(n_214),
.B1(n_163),
.B2(n_164),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_404),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_422),
.Y(n_591)
);

INVx11_ASAP7_75t_L g592 ( 
.A(n_453),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_449),
.B(n_240),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_453),
.A2(n_182),
.B1(n_261),
.B2(n_211),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_440),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_455),
.B(n_344),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_440),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_445),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_445),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_455),
.B(n_351),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_445),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_445),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_445),
.Y(n_604)
);

AOI21x1_ASAP7_75t_L g605 ( 
.A1(n_449),
.A2(n_248),
.B(n_243),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_411),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_449),
.A2(n_164),
.B1(n_214),
.B2(n_282),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_449),
.A2(n_282),
.B1(n_306),
.B2(n_270),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_572),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_580),
.B(n_382),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_596),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_530),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_596),
.Y(n_613)
);

AO22x2_ASAP7_75t_L g614 ( 
.A1(n_462),
.A2(n_266),
.B1(n_256),
.B2(n_304),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_514),
.B(n_395),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_477),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_477),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_485),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_469),
.A2(n_306),
.B1(n_451),
.B2(n_313),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_514),
.B(n_170),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_462),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_471),
.B(n_236),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_482),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_479),
.B(n_362),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_479),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_575),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_493),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_487),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_493),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_575),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_468),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_519),
.B(n_534),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_534),
.B(n_557),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_461),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_590),
.B(n_425),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_487),
.B(n_236),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_530),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_465),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_519),
.B(n_264),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_607),
.A2(n_312),
.B1(n_242),
.B2(n_301),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_475),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_484),
.B(n_395),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_486),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_489),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_590),
.B(n_382),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_579),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_497),
.B(n_395),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_503),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_592),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_601),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_505),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_515),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_500),
.B(n_383),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_518),
.B(n_362),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_592),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_526),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_521),
.B(n_363),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_SL g664 ( 
.A1(n_526),
.A2(n_276),
.B1(n_275),
.B2(n_273),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_524),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_525),
.B(n_363),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_468),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_507),
.B(n_300),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_537),
.B(n_543),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_474),
.B(n_269),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_544),
.B(n_366),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_472),
.A2(n_451),
.B1(n_294),
.B2(n_245),
.Y(n_673)
);

INVxp67_ASAP7_75t_SL g674 ( 
.A(n_523),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_547),
.B(n_395),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_549),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_583),
.Y(n_677)
);

NAND2x1p5_ASAP7_75t_L g678 ( 
.A(n_593),
.B(n_407),
.Y(n_678)
);

BUFx4f_ASAP7_75t_L g679 ( 
.A(n_526),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_468),
.Y(n_680)
);

NAND3x1_ASAP7_75t_L g681 ( 
.A(n_589),
.B(n_389),
.C(n_388),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_539),
.B(n_407),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_526),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_483),
.B(n_300),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_532),
.B(n_312),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_538),
.B(n_366),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_535),
.A2(n_451),
.B1(n_285),
.B2(n_268),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_554),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_533),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_595),
.B(n_271),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_583),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_570),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_460),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_516),
.B(n_407),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_463),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_542),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_538),
.B(n_492),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_545),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_571),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_460),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_466),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_512),
.A2(n_407),
.B1(n_528),
.B2(n_458),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_466),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_470),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_512),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_516),
.B(n_517),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_463),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_470),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_473),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_473),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_480),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_512),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_492),
.B(n_370),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_517),
.B(n_428),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_608),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_478),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_496),
.B(n_370),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_464),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_478),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_490),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_490),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_568),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_522),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_468),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_491),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_522),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_531),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_508),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_540),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_496),
.B(n_373),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_459),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_499),
.B(n_302),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_595),
.B(n_451),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_L g736 ( 
.A(n_550),
.B(n_458),
.C(n_428),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_373),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_488),
.B(n_383),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_491),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_531),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_494),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_571),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_536),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_459),
.A2(n_386),
.B1(n_374),
.B2(n_377),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_536),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_541),
.B(n_428),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_458),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_510),
.B(n_374),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_520),
.B(n_302),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_476),
.A2(n_301),
.B1(n_207),
.B2(n_272),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_510),
.B(n_308),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_494),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_587),
.B(n_377),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_476),
.B(n_378),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_541),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_546),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_546),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_551),
.B(n_308),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_463),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_556),
.B(n_238),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_571),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_561),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_550),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_508),
.Y(n_764)
);

BUFx10_ASAP7_75t_L g765 ( 
.A(n_527),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_562),
.B(n_238),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_552),
.B(n_555),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_552),
.B(n_428),
.Y(n_768)
);

AND2x2_ASAP7_75t_SL g769 ( 
.A(n_582),
.B(n_378),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_504),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_559),
.B(n_458),
.C(n_428),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_586),
.B(n_309),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_504),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_559),
.A2(n_380),
.B1(n_347),
.B2(n_3),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_594),
.B(n_309),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_506),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_527),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_555),
.B(n_428),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_527),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_506),
.Y(n_780)
);

AO22x2_ASAP7_75t_L g781 ( 
.A1(n_498),
.A2(n_509),
.B1(n_380),
.B2(n_560),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_696),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_655),
.B(n_553),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_777),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_609),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_777),
.B(n_498),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_655),
.B(n_567),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_637),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_688),
.A2(n_558),
.B1(n_509),
.B2(n_528),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_636),
.B(n_257),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_641),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_674),
.B(n_563),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_674),
.A2(n_558),
.B1(n_573),
.B2(n_569),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_692),
.B(n_563),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_751),
.A2(n_598),
.B(n_604),
.C(n_603),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_636),
.B(n_635),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_654),
.B(n_597),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_689),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_777),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_630),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_635),
.B(n_564),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_619),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_654),
.B(n_597),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_630),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_645),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_620),
.B(n_495),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_644),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_731),
.B(n_685),
.Y(n_809)
);

AND2x6_ASAP7_75t_L g810 ( 
.A(n_723),
.B(n_598),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_615),
.Y(n_811)
);

NAND2x1p5_ASAP7_75t_L g812 ( 
.A(n_620),
.B(n_495),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_749),
.B(n_599),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_668),
.B(n_599),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_668),
.B(n_600),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_731),
.B(n_577),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_646),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_633),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_642),
.A2(n_558),
.B1(n_591),
.B2(n_603),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_685),
.B(n_495),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_658),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_651),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_662),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_612),
.B(n_640),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_616),
.B(n_564),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_679),
.B(n_258),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_648),
.Y(n_827)
);

INVx6_ASAP7_75t_L g828 ( 
.A(n_765),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_724),
.A2(n_558),
.B1(n_528),
.B2(n_481),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_623),
.B(n_501),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_616),
.B(n_511),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_660),
.B(n_600),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_698),
.B(n_511),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_670),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_677),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_700),
.B(n_513),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_661),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_R g838 ( 
.A(n_779),
.B(n_719),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_611),
.B(n_613),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_649),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_623),
.B(n_347),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_769),
.B(n_513),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_SL g843 ( 
.A(n_660),
.B(n_196),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_653),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_639),
.A2(n_604),
.B(n_602),
.C(n_502),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_642),
.A2(n_558),
.B1(n_602),
.B2(n_481),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_763),
.B(n_558),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_661),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_686),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_679),
.B(n_262),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_699),
.B(n_742),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_691),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_693),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_758),
.B(n_502),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_695),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_702),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_699),
.B(n_742),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_656),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_683),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_763),
.B(n_502),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_762),
.B(n_566),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_657),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_626),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_665),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_676),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_682),
.B(n_566),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_761),
.B(n_628),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_761),
.B(n_501),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_627),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_631),
.B(n_501),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_631),
.B(n_184),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_682),
.B(n_566),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_694),
.A2(n_588),
.B(n_581),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_704),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_669),
.B(n_697),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_748),
.B(n_265),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_642),
.A2(n_748),
.B1(n_718),
.B2(n_732),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_639),
.B(n_191),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_627),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_632),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_738),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_686),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_706),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_712),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_705),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_617),
.B(n_581),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_712),
.Y(n_887)
);

NOR2x2_ASAP7_75t_L g888 ( 
.A(n_650),
.B(n_212),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_SL g889 ( 
.A(n_634),
.B(n_508),
.Y(n_889)
);

INVxp33_ASAP7_75t_L g890 ( 
.A(n_684),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_758),
.B(n_274),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_618),
.Y(n_892)
);

O2A1O1Ixp5_ASAP7_75t_L g893 ( 
.A1(n_624),
.A2(n_605),
.B(n_581),
.C(n_588),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_610),
.B(n_647),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_625),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_733),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_714),
.B(n_718),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_709),
.Y(n_898)
);

BUFx6f_ASAP7_75t_SL g899 ( 
.A(n_765),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_669),
.B(n_576),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_710),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_684),
.B(n_194),
.Y(n_902)
);

AO22x2_ASAP7_75t_L g903 ( 
.A1(n_750),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_725),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_728),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_714),
.A2(n_606),
.B(n_584),
.C(n_576),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_729),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_740),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_733),
.B(n_588),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_642),
.A2(n_481),
.B1(n_606),
.B2(n_584),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_732),
.A2(n_481),
.B1(n_206),
.B2(n_576),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_664),
.A2(n_716),
.B(n_643),
.C(n_683),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_743),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_671),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_634),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_671),
.A2(n_481),
.B1(n_606),
.B2(n_584),
.Y(n_916)
);

OAI22xp33_ASAP7_75t_L g917 ( 
.A1(n_621),
.A2(n_209),
.B1(n_202),
.B2(n_204),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_647),
.B(n_508),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_652),
.B(n_529),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_697),
.B(n_281),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_754),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_694),
.A2(n_481),
.B(n_400),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_745),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_687),
.B(n_283),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_755),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_756),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_722),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_737),
.Y(n_928)
);

BUFx5_ASAP7_75t_L g929 ( 
.A(n_735),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_716),
.A2(n_206),
.B1(n_212),
.B2(n_227),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_757),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_671),
.B(n_529),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_659),
.B(n_287),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_659),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_734),
.B(n_208),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_760),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_663),
.B(n_288),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_766),
.B(n_219),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_727),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_673),
.A2(n_290),
.B(n_291),
.C(n_296),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_739),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_741),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_643),
.B(n_212),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_737),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_634),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_663),
.B(n_585),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_666),
.B(n_298),
.Y(n_947)
);

AND2x6_ASAP7_75t_L g948 ( 
.A(n_753),
.B(n_585),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_753),
.Y(n_949)
);

OR2x6_ASAP7_75t_L g950 ( 
.A(n_650),
.B(n_585),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_671),
.B(n_574),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_666),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_SL g953 ( 
.A1(n_703),
.A2(n_413),
.B(n_400),
.C(n_414),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_672),
.B(n_585),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_667),
.B(n_565),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_672),
.B(n_650),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_744),
.A2(n_227),
.B1(n_297),
.B2(n_529),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_752),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_622),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_744),
.A2(n_227),
.B1(n_574),
.B2(n_529),
.Y(n_960)
);

NOR2x1p5_ASAP7_75t_L g961 ( 
.A(n_652),
.B(n_259),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_770),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_701),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_773),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_SL g965 ( 
.A1(n_713),
.A2(n_253),
.B1(n_235),
.B2(n_246),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_711),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_775),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_695),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_SL g969 ( 
.A1(n_750),
.A2(n_221),
.B1(n_247),
.B2(n_249),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_744),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_675),
.B(n_574),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_667),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_708),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_717),
.B(n_574),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_894),
.B(n_675),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_903),
.A2(n_774),
.B1(n_614),
.B2(n_664),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_868),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_897),
.A2(n_772),
.B1(n_681),
.B2(n_735),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_921),
.B(n_614),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_782),
.Y(n_980)
);

CKINVDCx6p67_ASAP7_75t_R g981 ( 
.A(n_799),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_869),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_879),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_808),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_853),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_868),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_788),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_935),
.A2(n_736),
.B(n_771),
.C(n_703),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_896),
.Y(n_989)
);

BUFx6f_ASAP7_75t_SL g990 ( 
.A(n_784),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_894),
.B(n_707),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_890),
.B(n_720),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_856),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_875),
.B(n_708),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_784),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_821),
.B(n_759),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_811),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_801),
.B(n_707),
.Y(n_998)
);

AND3x1_ASAP7_75t_L g999 ( 
.A(n_943),
.B(n_614),
.C(n_774),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_921),
.B(n_747),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_801),
.B(n_767),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_783),
.B(n_897),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_884),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_834),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_887),
.B(n_721),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_897),
.B(n_767),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_784),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_863),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_809),
.B(n_759),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_896),
.B(n_747),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_903),
.A2(n_774),
.B1(n_781),
.B2(n_736),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_791),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_799),
.B(n_667),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_897),
.B(n_781),
.Y(n_1014)
);

AOI22x1_ASAP7_75t_L g1015 ( 
.A1(n_961),
.A2(n_781),
.B1(n_638),
.B2(n_678),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_806),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_800),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_SL g1018 ( 
.A1(n_820),
.A2(n_780),
.B(n_776),
.C(n_778),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_915),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_838),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_817),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_827),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_877),
.B(n_764),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_SL g1024 ( 
.A1(n_798),
.A2(n_251),
.B1(n_295),
.B2(n_252),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_837),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_792),
.B(n_778),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_792),
.B(n_768),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_848),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_833),
.B(n_768),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_912),
.A2(n_771),
.B(n_715),
.C(n_746),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_828),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_878),
.B(n_638),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_859),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_874),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_943),
.A2(n_690),
.B1(n_735),
.B2(n_678),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_824),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_915),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_950),
.B(n_764),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_800),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_833),
.B(n_715),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_836),
.B(n_794),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_875),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_915),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_836),
.B(n_746),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_885),
.Y(n_1045)
);

BUFx4f_ASAP7_75t_L g1046 ( 
.A(n_828),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_796),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_902),
.A2(n_843),
.B1(n_969),
.B2(n_970),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_804),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_967),
.B(n_278),
.C(n_284),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_794),
.B(n_787),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_839),
.B(n_735),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_839),
.B(n_764),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_SL g1055 ( 
.A(n_799),
.B(n_289),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_860),
.B(n_730),
.Y(n_1056)
);

OR2x6_ASAP7_75t_SL g1057 ( 
.A(n_914),
.B(n_293),
.Y(n_1057)
);

AND2x4_ASAP7_75t_SL g1058 ( 
.A(n_851),
.B(n_730),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_944),
.A2(n_730),
.B(n_726),
.C(n_680),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_957),
.A2(n_690),
.B1(n_726),
.B2(n_680),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_956),
.B(n_726),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_898),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_936),
.A2(n_680),
.B(n_413),
.C(n_400),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_840),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_901),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_927),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_816),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_860),
.B(n_690),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_841),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_829),
.A2(n_565),
.B1(n_413),
.B2(n_414),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_844),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_881),
.B(n_7),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_956),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_945),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_950),
.B(n_412),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_959),
.B(n_7),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_804),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_899),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_814),
.B(n_690),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_815),
.B(n_565),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_866),
.B(n_565),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_851),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_883),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_871),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_945),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_866),
.B(n_872),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_849),
.B(n_8),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_939),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_938),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_882),
.B(n_9),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_858),
.Y(n_1091)
);

AOI22x1_ASAP7_75t_L g1092 ( 
.A1(n_855),
.A2(n_414),
.B1(n_411),
.B2(n_565),
.Y(n_1092)
);

AND2x4_ASAP7_75t_SL g1093 ( 
.A(n_857),
.B(n_414),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_862),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_941),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_857),
.B(n_56),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_872),
.B(n_412),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_949),
.B(n_11),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_864),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_928),
.B(n_11),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_945),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_865),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_883),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_946),
.B(n_954),
.Y(n_1104)
);

AND2x6_ASAP7_75t_L g1105 ( 
.A(n_847),
.B(n_67),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_867),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_950),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_972),
.B(n_889),
.Y(n_1108)
);

CKINVDCx6p67_ASAP7_75t_R g1109 ( 
.A(n_899),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_934),
.B(n_15),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_965),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_942),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_786),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_867),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_972),
.B(n_72),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_825),
.B(n_412),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_L g1117 ( 
.A(n_892),
.B(n_43),
.Y(n_1117)
);

AO22x1_ASAP7_75t_L g1118 ( 
.A1(n_948),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_904),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_847),
.A2(n_842),
.B(n_880),
.C(n_940),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_946),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_790),
.B(n_18),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_954),
.B(n_85),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_825),
.B(n_412),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_786),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_958),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_920),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_895),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_980),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_991),
.A2(n_854),
.B(n_813),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1052),
.B(n_842),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_991),
.A2(n_919),
.B(n_971),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1038),
.Y(n_1133)
);

INVx5_ASAP7_75t_L g1134 ( 
.A(n_1038),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1067),
.B(n_917),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1069),
.B(n_876),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_987),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1012),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1016),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1021),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1086),
.A2(n_918),
.B(n_971),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1052),
.B(n_831),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1048),
.A2(n_891),
.B1(n_930),
.B2(n_843),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1038),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1022),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1064),
.Y(n_1146)
);

BUFx4_ASAP7_75t_SL g1147 ( 
.A(n_1031),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1082),
.B(n_797),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1041),
.B(n_831),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_1002),
.A2(n_932),
.B(n_951),
.Y(n_1150)
);

BUFx10_ASAP7_75t_L g1151 ( 
.A(n_990),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1041),
.B(n_830),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_977),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1071),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_989),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_989),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1019),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1073),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1019),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1028),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1004),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_990),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1086),
.A2(n_918),
.B(n_919),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1111),
.A2(n_826),
.B1(n_850),
.B2(n_924),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1091),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1094),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1048),
.A2(n_870),
.B(n_909),
.C(n_793),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1019),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1020),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1084),
.B(n_933),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1089),
.B(n_937),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1099),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1102),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_1096),
.B(n_1107),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1119),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_985),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1078),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_1037),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_1083),
.Y(n_1179)
);

INVxp67_ASAP7_75t_SL g1180 ( 
.A(n_975),
.Y(n_1180)
);

CKINVDCx11_ASAP7_75t_R g1181 ( 
.A(n_1057),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1109),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_977),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1037),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1046),
.B(n_948),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1028),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_993),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_1037),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1121),
.B(n_797),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1034),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1043),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1045),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_997),
.Y(n_1193)
);

NOR2x1_ASAP7_75t_SL g1194 ( 
.A(n_1075),
.B(n_786),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1033),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1008),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1043),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1062),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1046),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1003),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1065),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1049),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_995),
.Y(n_1203)
);

BUFx5_ASAP7_75t_L g1204 ( 
.A(n_1105),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1010),
.Y(n_1205)
);

AOI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1079),
.A2(n_873),
.B(n_974),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1066),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_995),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_976),
.A2(n_907),
.B1(n_966),
.B2(n_905),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1088),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_998),
.A2(n_922),
.B(n_789),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1043),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_998),
.A2(n_922),
.B(n_953),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1095),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1112),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1067),
.B(n_947),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1001),
.B(n_861),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_986),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1001),
.B(n_861),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1126),
.Y(n_1220)
);

CKINVDCx14_ASAP7_75t_R g1221 ( 
.A(n_1103),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_984),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_981),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1042),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1025),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1074),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_986),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1074),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_976),
.A2(n_908),
.B1(n_913),
.B2(n_923),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1036),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_982),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_983),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1054),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1113),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1011),
.A2(n_925),
.B1(n_926),
.B2(n_963),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1007),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1128),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1121),
.B(n_973),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1074),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1054),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1127),
.A2(n_948),
.B1(n_900),
.B2(n_832),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_979),
.B(n_852),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_975),
.B(n_810),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_994),
.B(n_832),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_994),
.B(n_803),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1000),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1047),
.B(n_931),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1007),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1047),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1017),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1107),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1025),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1107),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_992),
.B(n_805),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1017),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1005),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1005),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1125),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1011),
.A2(n_960),
.B1(n_948),
.B2(n_835),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_999),
.A2(n_911),
.B1(n_906),
.B2(n_973),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1122),
.A2(n_785),
.B1(n_822),
.B2(n_818),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1056),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1056),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1039),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1039),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1104),
.B(n_803),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1035),
.A2(n_968),
.B1(n_855),
.B2(n_807),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1101),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1101),
.Y(n_1269)
);

OAI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1076),
.A2(n_992),
.B1(n_1100),
.B2(n_1051),
.C(n_1072),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1029),
.B(n_810),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1058),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1050),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1050),
.Y(n_1274)
);

INVx8_ASAP7_75t_L g1275 ( 
.A(n_1101),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1098),
.A2(n_802),
.B1(n_823),
.B2(n_962),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1096),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1035),
.A2(n_988),
.B1(n_1060),
.B2(n_1026),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1026),
.A2(n_845),
.B(n_795),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1077),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1060),
.A2(n_968),
.B1(n_807),
.B2(n_812),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1032),
.A2(n_964),
.B1(n_810),
.B2(n_929),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1013),
.Y(n_1283)
);

OAI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1270),
.A2(n_1055),
.B1(n_978),
.B2(n_1002),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_SL g1285 ( 
.A(n_1185),
.B(n_1134),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1137),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1242),
.B(n_1090),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1279),
.A2(n_1030),
.B(n_1079),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1167),
.A2(n_1120),
.B(n_1068),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1138),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1130),
.A2(n_1068),
.B(n_1053),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1275),
.Y(n_1292)
);

INVx8_ASAP7_75t_L g1293 ( 
.A(n_1275),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1279),
.A2(n_1015),
.B(n_1080),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1206),
.A2(n_1097),
.B(n_1124),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1200),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1139),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1213),
.A2(n_1018),
.B(n_1080),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1161),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1135),
.A2(n_1009),
.B(n_1117),
.C(n_996),
.Y(n_1300)
);

AO21x2_ASAP7_75t_L g1301 ( 
.A1(n_1213),
.A2(n_1059),
.B(n_1014),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1141),
.A2(n_1097),
.B(n_1116),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1135),
.A2(n_1024),
.B1(n_1105),
.B2(n_1118),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1134),
.B(n_1106),
.Y(n_1304)
);

AOI22x1_ASAP7_75t_L g1305 ( 
.A1(n_1180),
.A2(n_1108),
.B1(n_1013),
.B2(n_1115),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1140),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1130),
.A2(n_1081),
.B(n_1014),
.Y(n_1307)
);

BUFx12f_ASAP7_75t_L g1308 ( 
.A(n_1151),
.Y(n_1308)
);

AOI21xp33_ASAP7_75t_L g1309 ( 
.A1(n_1278),
.A2(n_1053),
.B(n_1027),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1180),
.A2(n_1027),
.B1(n_1087),
.B2(n_1029),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1205),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1211),
.A2(n_1040),
.B(n_1044),
.Y(n_1312)
);

INVx8_ASAP7_75t_L g1313 ( 
.A(n_1275),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1278),
.A2(n_1006),
.B(n_1124),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1174),
.B(n_1114),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1143),
.A2(n_1270),
.B1(n_1216),
.B2(n_1170),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1216),
.A2(n_1105),
.B1(n_1110),
.B2(n_1115),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1141),
.A2(n_1116),
.B(n_1081),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1150),
.A2(n_1063),
.B(n_1040),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1129),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1211),
.A2(n_1023),
.B(n_1006),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1146),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1174),
.B(n_1108),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1165),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1147),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1283),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1143),
.B(n_1123),
.C(n_1061),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1283),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1131),
.B(n_1044),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1164),
.A2(n_1077),
.B1(n_819),
.B2(n_846),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1283),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1175),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1174),
.B(n_1075),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1202),
.Y(n_1334)
);

NAND2x1_ASAP7_75t_L g1335 ( 
.A(n_1153),
.B(n_1105),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1194),
.A2(n_1092),
.B(n_1085),
.Y(n_1336)
);

AND2x6_ASAP7_75t_SL g1337 ( 
.A(n_1171),
.B(n_1075),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1178),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1133),
.B(n_886),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1163),
.A2(n_893),
.B(n_1070),
.Y(n_1340)
);

NOR2xp67_ASAP7_75t_L g1341 ( 
.A(n_1169),
.B(n_1085),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1189),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1131),
.B(n_1105),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1145),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1205),
.B(n_1254),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1163),
.A2(n_1070),
.B(n_929),
.Y(n_1346)
);

AOI222xp33_ASAP7_75t_L g1347 ( 
.A1(n_1256),
.A2(n_888),
.B1(n_810),
.B2(n_23),
.C1(n_30),
.C2(n_31),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1154),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1277),
.B(n_1093),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1132),
.A2(n_886),
.B(n_812),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1142),
.B(n_929),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1166),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1232),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1247),
.B(n_916),
.C(n_910),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1132),
.A2(n_955),
.B(n_929),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1152),
.A2(n_955),
.B(n_929),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1152),
.A2(n_412),
.B(n_98),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1267),
.A2(n_86),
.B(n_148),
.Y(n_1358)
);

BUFx8_ASAP7_75t_L g1359 ( 
.A(n_1196),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1142),
.B(n_21),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1267),
.A2(n_100),
.B(n_127),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1149),
.A2(n_77),
.B(n_121),
.Y(n_1362)
);

OR2x6_ASAP7_75t_L g1363 ( 
.A(n_1133),
.B(n_153),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1246),
.B(n_22),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1136),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_SL g1366 ( 
.A1(n_1259),
.A2(n_33),
.B(n_34),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1172),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1277),
.A2(n_35),
.B(n_38),
.C(n_107),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1244),
.B(n_111),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1178),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1266),
.A2(n_35),
.B1(n_38),
.B2(n_115),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1281),
.A2(n_1271),
.B(n_1219),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1259),
.A2(n_1257),
.B1(n_1149),
.B2(n_1134),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1187),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_SL g1375 ( 
.A1(n_1271),
.A2(n_1217),
.B(n_1219),
.C(n_1243),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1155),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1281),
.A2(n_1217),
.B(n_1276),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1151),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1173),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1243),
.A2(n_1282),
.B(n_1262),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1260),
.A2(n_1282),
.B(n_1263),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1260),
.A2(n_1233),
.B(n_1240),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1231),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1185),
.A2(n_1134),
.B1(n_1204),
.B2(n_1249),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1156),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1195),
.B(n_1158),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1238),
.A2(n_1280),
.B(n_1274),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1176),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1160),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1247),
.A2(n_1241),
.B(n_1276),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1264),
.A2(n_1273),
.A3(n_1265),
.B(n_1255),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1209),
.A2(n_1229),
.B1(n_1235),
.B2(n_1144),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1195),
.B(n_1186),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1144),
.B(n_1162),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1190),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1261),
.A2(n_1209),
.B(n_1229),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1266),
.A2(n_1224),
.B1(n_1244),
.B2(n_1245),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1193),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1238),
.A2(n_1218),
.B(n_1153),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1225),
.B(n_1252),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1183),
.A2(n_1218),
.B(n_1227),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1210),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1268),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1183),
.A2(n_1227),
.B(n_1235),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1192),
.B(n_1201),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1261),
.B(n_1215),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1198),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1237),
.B(n_1148),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1207),
.Y(n_1409)
);

INVx6_ASAP7_75t_L g1410 ( 
.A(n_1178),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1214),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1222),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1250),
.A2(n_1220),
.B(n_1204),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1178),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1272),
.A2(n_1204),
.B(n_1188),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1245),
.A2(n_1258),
.B1(n_1148),
.B2(n_1199),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1230),
.B(n_1177),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1204),
.A2(n_1179),
.B1(n_1189),
.B2(n_1181),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1204),
.B(n_1253),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1272),
.B(n_1251),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1204),
.A2(n_1188),
.B(n_1184),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1184),
.A2(n_1188),
.B(n_1203),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1236),
.A2(n_1248),
.B(n_1188),
.C(n_1184),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1184),
.B(n_1162),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1203),
.B(n_1212),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1157),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1157),
.B(n_1269),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1157),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1159),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1159),
.B(n_1269),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1159),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1286),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1345),
.B(n_1269),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1306),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1347),
.A2(n_1221),
.B1(n_1234),
.B2(n_1208),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1287),
.B(n_1212),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1316),
.A2(n_1223),
.B1(n_1182),
.B2(n_1168),
.C(n_1191),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1338),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1393),
.B(n_1212),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1296),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1332),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1370),
.Y(n_1442)
);

OAI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1347),
.A2(n_1168),
.B1(n_1191),
.B2(n_1197),
.C(n_1226),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1370),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1373),
.B(n_1390),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1405),
.B(n_1168),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1295),
.A2(n_1191),
.B(n_1197),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1285),
.A2(n_1197),
.B1(n_1226),
.B2(n_1228),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1318),
.A2(n_1226),
.B(n_1228),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1311),
.B(n_1228),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1303),
.A2(n_1147),
.B1(n_1239),
.B2(n_1365),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1303),
.A2(n_1239),
.B1(n_1284),
.B2(n_1390),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_1308),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1320),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1302),
.A2(n_1239),
.B(n_1350),
.Y(n_1455)
);

BUFx8_ASAP7_75t_SL g1456 ( 
.A(n_1325),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1333),
.B(n_1315),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1344),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1353),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1368),
.A2(n_1423),
.B(n_1300),
.C(n_1362),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1311),
.B(n_1360),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1299),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1374),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1370),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1348),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1352),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1382),
.B(n_1305),
.Y(n_1467)
);

NAND2xp33_ASAP7_75t_R g1468 ( 
.A(n_1380),
.B(n_1323),
.Y(n_1468)
);

OAI222xp33_ASAP7_75t_L g1469 ( 
.A1(n_1392),
.A2(n_1373),
.B1(n_1371),
.B2(n_1317),
.C1(n_1384),
.C2(n_1329),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1376),
.B(n_1385),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1376),
.Y(n_1471)
);

AOI21xp33_ASAP7_75t_L g1472 ( 
.A1(n_1327),
.A2(n_1289),
.B(n_1330),
.Y(n_1472)
);

CKINVDCx16_ASAP7_75t_R g1473 ( 
.A(n_1417),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1346),
.A2(n_1340),
.B(n_1355),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1355),
.A2(n_1291),
.B(n_1312),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1359),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1385),
.B(n_1389),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1396),
.A2(n_1392),
.B1(n_1289),
.B2(n_1362),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1396),
.A2(n_1366),
.B1(n_1360),
.B2(n_1317),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1397),
.A2(n_1416),
.B1(n_1418),
.B2(n_1384),
.Y(n_1480)
);

AOI21xp33_ASAP7_75t_L g1481 ( 
.A1(n_1310),
.A2(n_1354),
.B(n_1291),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1338),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1337),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_SL g1484 ( 
.A1(n_1329),
.A2(n_1422),
.B(n_1414),
.C(n_1408),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1285),
.A2(n_1363),
.B1(n_1364),
.B2(n_1400),
.Y(n_1485)
);

BUFx10_ASAP7_75t_L g1486 ( 
.A(n_1386),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1367),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1312),
.A2(n_1314),
.B(n_1381),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1389),
.B(n_1290),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1407),
.B(n_1409),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1309),
.A2(n_1314),
.B1(n_1310),
.B2(n_1377),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1333),
.B(n_1315),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1359),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1379),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1297),
.B(n_1322),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1334),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1426),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1398),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_L g1499 ( 
.A1(n_1406),
.A2(n_1343),
.B(n_1321),
.Y(n_1499)
);

OAI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1309),
.A2(n_1363),
.B1(n_1412),
.B2(n_1394),
.C(n_1343),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1341),
.A2(n_1323),
.B1(n_1394),
.B2(n_1419),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1358),
.A2(n_1361),
.B(n_1335),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1323),
.A2(n_1394),
.B1(n_1419),
.B2(n_1406),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1372),
.A2(n_1356),
.B(n_1387),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1426),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1383),
.Y(n_1506)
);

CKINVDCx9p33_ASAP7_75t_R g1507 ( 
.A(n_1403),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1338),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1342),
.A2(n_1363),
.B1(n_1424),
.B2(n_1304),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1378),
.Y(n_1510)
);

BUFx12f_ASAP7_75t_L g1511 ( 
.A(n_1292),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1324),
.B(n_1411),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1388),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1427),
.B(n_1342),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1395),
.B(n_1402),
.Y(n_1515)
);

INVx6_ASAP7_75t_L g1516 ( 
.A(n_1293),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1377),
.A2(n_1369),
.B1(n_1321),
.B2(n_1288),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1391),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1307),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1420),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1307),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1375),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1422),
.B(n_1415),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1369),
.A2(n_1288),
.B1(n_1351),
.B2(n_1380),
.Y(n_1524)
);

BUFx4f_ASAP7_75t_L g1525 ( 
.A(n_1292),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1414),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_SL g1527 ( 
.A(n_1356),
.B(n_1304),
.C(n_1424),
.Y(n_1527)
);

OAI22x1_ASAP7_75t_L g1528 ( 
.A1(n_1428),
.A2(n_1357),
.B1(n_1420),
.B2(n_1319),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1351),
.B(n_1331),
.Y(n_1529)
);

AOI21xp33_ASAP7_75t_L g1530 ( 
.A1(n_1301),
.A2(n_1298),
.B(n_1294),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_R g1531 ( 
.A(n_1339),
.B(n_1357),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1431),
.B(n_1429),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1326),
.B(n_1331),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1326),
.B(n_1328),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1301),
.A2(n_1319),
.B1(n_1349),
.B2(n_1339),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1349),
.A2(n_1339),
.B1(n_1298),
.B2(n_1404),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1410),
.A2(n_1294),
.B1(n_1421),
.B2(n_1313),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1328),
.B(n_1429),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1293),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1410),
.A2(n_1292),
.B1(n_1425),
.B2(n_1313),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1410),
.B(n_1425),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1413),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1430),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1413),
.A2(n_1336),
.B1(n_1313),
.B2(n_1293),
.Y(n_1544)
);

AOI21xp33_ASAP7_75t_L g1545 ( 
.A1(n_1401),
.A2(n_1399),
.B(n_1430),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1345),
.B(n_1316),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1400),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1296),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1285),
.A2(n_943),
.B1(n_685),
.B2(n_1270),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1400),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1316),
.A2(n_1048),
.B1(n_1111),
.B2(n_1143),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1312),
.A2(n_1180),
.B(n_1130),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1461),
.B(n_1478),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_R g1554 ( 
.A(n_1440),
.B(n_1548),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1456),
.Y(n_1555)
);

AND2x2_ASAP7_75t_SL g1556 ( 
.A(n_1478),
.B(n_1452),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1450),
.B(n_1514),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1458),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1481),
.B(n_1471),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1470),
.B(n_1477),
.Y(n_1560)
);

NAND2xp33_ASAP7_75t_R g1561 ( 
.A(n_1476),
.B(n_1462),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1472),
.A2(n_1435),
.B(n_1551),
.C(n_1443),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1549),
.A2(n_1445),
.B1(n_1480),
.B2(n_1473),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1436),
.B(n_1532),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1465),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1446),
.B(n_1439),
.Y(n_1566)
);

OR2x6_ASAP7_75t_L g1567 ( 
.A(n_1445),
.B(n_1523),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_R g1568 ( 
.A(n_1510),
.B(n_1539),
.Y(n_1568)
);

NOR3xp33_ASAP7_75t_SL g1569 ( 
.A(n_1453),
.B(n_1549),
.C(n_1500),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1466),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1457),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1507),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1457),
.B(n_1492),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1487),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1471),
.B(n_1494),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1435),
.A2(n_1451),
.B1(n_1452),
.B2(n_1479),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1552),
.A2(n_1460),
.B(n_1475),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_R g1578 ( 
.A(n_1483),
.B(n_1525),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1506),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1492),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1445),
.B(n_1523),
.Y(n_1581)
);

BUFx4f_ASAP7_75t_SL g1582 ( 
.A(n_1511),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1513),
.Y(n_1583)
);

INVxp33_ASAP7_75t_SL g1584 ( 
.A(n_1433),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1497),
.B(n_1505),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1451),
.A2(n_1485),
.B1(n_1479),
.B2(n_1437),
.Y(n_1586)
);

BUFx4f_ASAP7_75t_SL g1587 ( 
.A(n_1547),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1512),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1491),
.B(n_1503),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1526),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_SL g1593 ( 
.A(n_1550),
.B(n_1546),
.C(n_1496),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1432),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1499),
.B(n_1515),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1489),
.B(n_1524),
.Y(n_1596)
);

NAND2xp33_ASAP7_75t_R g1597 ( 
.A(n_1541),
.B(n_1444),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1528),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1434),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1543),
.B(n_1520),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1507),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_R g1602 ( 
.A(n_1525),
.B(n_1493),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1518),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1441),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1524),
.B(n_1522),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_R g1606 ( 
.A(n_1541),
.B(n_1464),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1468),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1495),
.Y(n_1608)
);

CKINVDCx16_ASAP7_75t_R g1609 ( 
.A(n_1486),
.Y(n_1609)
);

NOR2x1p5_ASAP7_75t_L g1610 ( 
.A(n_1438),
.B(n_1508),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1538),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1517),
.B(n_1535),
.C(n_1509),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1486),
.B(n_1490),
.Y(n_1613)
);

OR2x2_ASAP7_75t_SL g1614 ( 
.A(n_1527),
.B(n_1516),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1485),
.A2(n_1501),
.B1(n_1527),
.B2(n_1498),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_R g1616 ( 
.A(n_1442),
.B(n_1444),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1542),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1459),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1517),
.B(n_1521),
.Y(n_1619)
);

BUFx10_ASAP7_75t_L g1620 ( 
.A(n_1516),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1530),
.A2(n_1531),
.A3(n_1463),
.B(n_1467),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1469),
.A2(n_1488),
.B1(n_1516),
.B2(n_1482),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1474),
.A2(n_1467),
.B(n_1502),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1540),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_R g1625 ( 
.A(n_1442),
.B(n_1464),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1482),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_SL g1627 ( 
.A(n_1531),
.B(n_1468),
.C(n_1448),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1617),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1603),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1592),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1619),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1585),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1619),
.B(n_1521),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1558),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1565),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1567),
.B(n_1488),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1585),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1570),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1598),
.B(n_1519),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1567),
.B(n_1519),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1595),
.B(n_1559),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1574),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1607),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1579),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1583),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1567),
.B(n_1581),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1581),
.B(n_1504),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1581),
.B(n_1535),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1575),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1621),
.B(n_1536),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1621),
.B(n_1536),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1575),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1618),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1577),
.B(n_1455),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1591),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1594),
.Y(n_1656)
);

OR2x6_ASAP7_75t_L g1657 ( 
.A(n_1577),
.B(n_1449),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1621),
.Y(n_1658)
);

NAND2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1449),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1605),
.B(n_1537),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1599),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1605),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1596),
.B(n_1537),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1604),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1595),
.B(n_1545),
.Y(n_1665)
);

AND2x4_ASAP7_75t_SL g1666 ( 
.A(n_1627),
.B(n_1544),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1571),
.B(n_1580),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1589),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1620),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1608),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1556),
.A2(n_1469),
.B1(n_1482),
.B2(n_1508),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1571),
.B(n_1447),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1559),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1591),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1641),
.B(n_1611),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_1586),
.B1(n_1562),
.B2(n_1576),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1632),
.B(n_1560),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1641),
.B(n_1588),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1671),
.B(n_1569),
.C(n_1615),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1673),
.B(n_1563),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1673),
.B(n_1588),
.Y(n_1681)
);

OAI21xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1660),
.A2(n_1663),
.B(n_1632),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1665),
.B(n_1590),
.C(n_1622),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1666),
.A2(n_1590),
.B1(n_1612),
.B2(n_1553),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1665),
.B(n_1596),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1665),
.B(n_1553),
.C(n_1597),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1631),
.B(n_1557),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_SL g1688 ( 
.A1(n_1666),
.A2(n_1572),
.B1(n_1601),
.B2(n_1587),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1631),
.B(n_1613),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1662),
.B(n_1609),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1606),
.C(n_1484),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1649),
.B(n_1566),
.Y(n_1692)
);

OAI21xp33_ASAP7_75t_L g1693 ( 
.A1(n_1663),
.A2(n_1593),
.B(n_1612),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1632),
.B(n_1564),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1649),
.B(n_1593),
.Y(n_1695)
);

NOR3xp33_ASAP7_75t_SL g1696 ( 
.A(n_1652),
.B(n_1561),
.C(n_1555),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1643),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1660),
.A2(n_1448),
.B1(n_1544),
.B2(n_1533),
.C(n_1534),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1666),
.A2(n_1580),
.B1(n_1624),
.B2(n_1600),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1630),
.B(n_1573),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1666),
.A2(n_1438),
.B(n_1482),
.Y(n_1702)
);

OAI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1660),
.A2(n_1578),
.B(n_1600),
.Y(n_1703)
);

NAND2xp33_ASAP7_75t_SL g1704 ( 
.A(n_1669),
.B(n_1602),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1633),
.A2(n_1625),
.B1(n_1616),
.B2(n_1568),
.C(n_1626),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1630),
.B(n_1610),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1633),
.A2(n_1614),
.B1(n_1582),
.B2(n_1554),
.C(n_1620),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_1668),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1648),
.A2(n_1650),
.B(n_1651),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1670),
.B(n_1668),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1670),
.B(n_1662),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1662),
.B(n_1653),
.Y(n_1712)
);

OAI221xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1650),
.A2(n_1651),
.B1(n_1648),
.B2(n_1658),
.C(n_1633),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1662),
.B(n_1653),
.Y(n_1714)
);

NAND4xp25_ASAP7_75t_L g1715 ( 
.A(n_1650),
.B(n_1651),
.C(n_1639),
.D(n_1658),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1662),
.B(n_1653),
.Y(n_1716)
);

OAI31xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1646),
.A2(n_1648),
.A3(n_1636),
.B(n_1647),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1646),
.A2(n_1636),
.B(n_1647),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1678),
.B(n_1662),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1681),
.B(n_1662),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1717),
.B(n_1646),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1711),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1712),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1662),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1708),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1685),
.B(n_1637),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1690),
.B(n_1647),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1697),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1690),
.B(n_1640),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1677),
.B(n_1640),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1693),
.A2(n_1658),
.B1(n_1636),
.B2(n_1639),
.C(n_1640),
.Y(n_1732)
);

NAND2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1680),
.B(n_1639),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1714),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1710),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1718),
.B(n_1674),
.Y(n_1737)
);

OA211x2_ASAP7_75t_L g1738 ( 
.A1(n_1693),
.A2(n_1669),
.B(n_1657),
.C(n_1659),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1715),
.B(n_1656),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1677),
.B(n_1674),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1713),
.B(n_1656),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1680),
.B(n_1669),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1691),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1716),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1687),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1689),
.B(n_1674),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1692),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1675),
.Y(n_1748)
);

NAND2x1p5_ASAP7_75t_L g1749 ( 
.A(n_1702),
.B(n_1669),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1686),
.B(n_1655),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1694),
.B(n_1655),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1683),
.B(n_1657),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1694),
.B(n_1655),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1703),
.B(n_1669),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1706),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1725),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1739),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1725),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1735),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1721),
.B(n_1729),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1721),
.B(n_1709),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1743),
.A2(n_1679),
.B1(n_1684),
.B2(n_1688),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1729),
.B(n_1667),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1735),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1747),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1736),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1747),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1728),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1742),
.B(n_1704),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1739),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1707),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1741),
.B(n_1698),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1741),
.B(n_1661),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1733),
.B(n_1661),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1736),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1733),
.A2(n_1676),
.B(n_1705),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1733),
.B(n_1656),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1722),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1722),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1737),
.B(n_1667),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1724),
.B(n_1661),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1723),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1745),
.B(n_1744),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1745),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1750),
.B(n_1699),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1737),
.B(n_1672),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1748),
.B(n_1751),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1748),
.B(n_1644),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1727),
.B(n_1730),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_L g1791 ( 
.A(n_1727),
.B(n_1642),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1727),
.B(n_1667),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1730),
.B(n_1667),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1730),
.B(n_1667),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1755),
.B(n_1726),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1672),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1731),
.B(n_1672),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1744),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1776),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1790),
.Y(n_1800)
);

OAI21xp33_ASAP7_75t_L g1801 ( 
.A1(n_1786),
.A2(n_1753),
.B(n_1732),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1763),
.B(n_1742),
.Y(n_1802)
);

OAI222xp33_ASAP7_75t_L g1803 ( 
.A1(n_1762),
.A2(n_1753),
.B1(n_1742),
.B2(n_1773),
.C1(n_1770),
.C2(n_1761),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1761),
.B(n_1753),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1776),
.B(n_1753),
.Y(n_1805)
);

OAI33xp33_ASAP7_75t_L g1806 ( 
.A1(n_1771),
.A2(n_1719),
.A3(n_1720),
.B1(n_1634),
.B2(n_1644),
.B3(n_1645),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1762),
.B(n_1731),
.Y(n_1807)
);

OAI211xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1777),
.A2(n_1696),
.B(n_1700),
.C(n_1746),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1790),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1766),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1771),
.B(n_1704),
.C(n_1723),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1781),
.B(n_1740),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1768),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1773),
.A2(n_1738),
.B1(n_1749),
.B2(n_1740),
.Y(n_1816)
);

AO22x1_ASAP7_75t_L g1817 ( 
.A1(n_1772),
.A2(n_1669),
.B1(n_1752),
.B2(n_1754),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1795),
.A2(n_1749),
.B1(n_1734),
.B2(n_1754),
.Y(n_1818)
);

OAI322xp33_ASAP7_75t_L g1819 ( 
.A1(n_1758),
.A2(n_1749),
.A3(n_1734),
.B1(n_1634),
.B2(n_1645),
.C1(n_1628),
.C2(n_1629),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1758),
.A2(n_1752),
.B(n_1657),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1768),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1767),
.A2(n_1669),
.B1(n_1657),
.B2(n_1654),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1767),
.A2(n_1669),
.B(n_1672),
.C(n_1628),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1774),
.B(n_1664),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1757),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1774),
.A2(n_1657),
.B1(n_1654),
.B2(n_1659),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1757),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1759),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1775),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1781),
.B(n_1672),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1788),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1791),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1775),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1799),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1807),
.B(n_1793),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1799),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1811),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1807),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1800),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1800),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1809),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1809),
.Y(n_1842)
);

OR2x6_ASAP7_75t_L g1843 ( 
.A(n_1810),
.B(n_1812),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1831),
.B(n_1785),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1829),
.B(n_1785),
.Y(n_1845)
);

OAI31xp33_ASAP7_75t_L g1846 ( 
.A1(n_1801),
.A2(n_1778),
.A3(n_1765),
.B(n_1760),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1804),
.B(n_1793),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1805),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1802),
.B(n_1760),
.Y(n_1849)
);

NOR3xp33_ASAP7_75t_L g1850 ( 
.A(n_1803),
.B(n_1765),
.C(n_1759),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1805),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1813),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1832),
.B(n_1791),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1808),
.A2(n_1798),
.B(n_1784),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1829),
.B(n_1789),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1833),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1815),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1814),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1856),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1839),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1834),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1846),
.A2(n_1854),
.B1(n_1850),
.B2(n_1844),
.C(n_1849),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1835),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1843),
.A2(n_1818),
.B1(n_1816),
.B2(n_1822),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1843),
.A2(n_1817),
.B(n_1819),
.Y(n_1865)
);

OAI32xp33_ASAP7_75t_L g1866 ( 
.A1(n_1838),
.A2(n_1804),
.A3(n_1820),
.B1(n_1821),
.B2(n_1828),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1834),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1839),
.B(n_1833),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1835),
.B(n_1794),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1836),
.Y(n_1870)
);

NAND2xp33_ASAP7_75t_L g1871 ( 
.A(n_1848),
.B(n_1823),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1843),
.A2(n_1823),
.B1(n_1787),
.B2(n_1794),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1836),
.Y(n_1873)
);

AOI322xp5_ASAP7_75t_L g1874 ( 
.A1(n_1858),
.A2(n_1826),
.A3(n_1827),
.B1(n_1825),
.B2(n_1787),
.C1(n_1764),
.C2(n_1792),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1845),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1837),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1863),
.B(n_1848),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1860),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1862),
.A2(n_1846),
.B1(n_1843),
.B2(n_1851),
.C(n_1840),
.Y(n_1880)
);

NAND2x1_ASAP7_75t_SL g1881 ( 
.A(n_1860),
.B(n_1853),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1862),
.A2(n_1843),
.B1(n_1851),
.B2(n_1858),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1868),
.Y(n_1883)
);

NOR2x1_ASAP7_75t_L g1884 ( 
.A(n_1859),
.B(n_1842),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1868),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1875),
.B(n_1840),
.Y(n_1886)
);

AO22x2_ASAP7_75t_L g1887 ( 
.A1(n_1877),
.A2(n_1841),
.B1(n_1842),
.B2(n_1857),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1876),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1879),
.Y(n_1889)
);

AOI221x1_ASAP7_75t_L g1890 ( 
.A1(n_1882),
.A2(n_1865),
.B1(n_1873),
.B2(n_1861),
.C(n_1870),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1887),
.Y(n_1891)
);

OAI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1880),
.A2(n_1865),
.B1(n_1872),
.B2(n_1864),
.Y(n_1892)
);

NOR3xp33_ASAP7_75t_L g1893 ( 
.A(n_1884),
.B(n_1866),
.C(n_1867),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1883),
.B(n_1874),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1887),
.Y(n_1895)
);

XNOR2xp5_ASAP7_75t_L g1896 ( 
.A(n_1885),
.B(n_1847),
.Y(n_1896)
);

AOI32xp33_ASAP7_75t_L g1897 ( 
.A1(n_1888),
.A2(n_1871),
.A3(n_1841),
.B1(n_1853),
.B2(n_1847),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1881),
.B(n_1886),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1878),
.A2(n_1869),
.B1(n_1853),
.B2(n_1855),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1898),
.Y(n_1900)
);

NOR3xp33_ASAP7_75t_L g1901 ( 
.A(n_1892),
.B(n_1857),
.C(n_1852),
.Y(n_1901)
);

AO21x1_ASAP7_75t_L g1902 ( 
.A1(n_1891),
.A2(n_1852),
.B(n_1837),
.Y(n_1902)
);

OAI21xp33_ASAP7_75t_L g1903 ( 
.A1(n_1894),
.A2(n_1853),
.B(n_1830),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1896),
.B(n_1798),
.Y(n_1904)
);

AOI211x1_ASAP7_75t_L g1905 ( 
.A1(n_1895),
.A2(n_1826),
.B(n_1830),
.C(n_1792),
.Y(n_1905)
);

NOR3xp33_ASAP7_75t_L g1906 ( 
.A(n_1900),
.B(n_1889),
.C(n_1893),
.Y(n_1906)
);

NOR3x1_ASAP7_75t_L g1907 ( 
.A(n_1904),
.B(n_1897),
.C(n_1890),
.Y(n_1907)
);

NOR3x1_ASAP7_75t_L g1908 ( 
.A(n_1901),
.B(n_1899),
.C(n_1784),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1903),
.B(n_1783),
.Y(n_1909)
);

O2A1O1Ixp5_ASAP7_75t_L g1910 ( 
.A1(n_1902),
.A2(n_1806),
.B(n_1779),
.C(n_1780),
.Y(n_1910)
);

OAI21xp33_ASAP7_75t_L g1911 ( 
.A1(n_1905),
.A2(n_1787),
.B(n_1797),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1906),
.B(n_1783),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1909),
.Y(n_1913)
);

NOR2x1_ASAP7_75t_L g1914 ( 
.A(n_1907),
.B(n_1911),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1908),
.B(n_1779),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1910),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1914),
.A2(n_1787),
.B1(n_1764),
.B2(n_1797),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1916),
.B(n_1780),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1915),
.Y(n_1919)
);

NOR2xp67_ASAP7_75t_L g1920 ( 
.A(n_1918),
.B(n_1913),
.Y(n_1920)
);

CKINVDCx16_ASAP7_75t_R g1921 ( 
.A(n_1920),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1921),
.Y(n_1922)
);

NAND2xp33_ASAP7_75t_SL g1923 ( 
.A(n_1921),
.B(n_1912),
.Y(n_1923)
);

XNOR2xp5_ASAP7_75t_L g1924 ( 
.A(n_1922),
.B(n_1919),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1923),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1917),
.B1(n_1824),
.B2(n_1778),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1924),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1927),
.B(n_1796),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1928),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1929),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1930),
.A2(n_1926),
.B1(n_1796),
.B2(n_1782),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1931),
.A2(n_1659),
.B1(n_1629),
.B2(n_1635),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1782),
.B1(n_1635),
.B2(n_1638),
.C(n_1642),
.Y(n_1933)
);

AOI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1642),
.B(n_1638),
.C(n_1635),
.Y(n_1934)
);


endmodule