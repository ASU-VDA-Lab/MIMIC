module fake_jpeg_10724_n_131 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVxp67_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_1),
.B(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_28),
.Y(n_71)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_30),
.B(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_11),
.B(n_0),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_43),
.Y(n_76)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_3),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_3),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_12),
.B(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_12),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_13),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_24),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_29),
.B1(n_40),
.B2(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_28),
.B2(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_11),
.B(n_23),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_21),
.A3(n_44),
.B1(n_38),
.B2(n_11),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_73),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_27),
.B1(n_32),
.B2(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_37),
.B1(n_39),
.B2(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_42),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_27),
.B1(n_32),
.B2(n_15),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_48),
.B1(n_47),
.B2(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_77),
.B1(n_69),
.B2(n_58),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_38),
.B(n_28),
.C(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_73),
.B1(n_67),
.B2(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_59),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_64),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_77),
.B1(n_57),
.B2(n_64),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_93),
.B(n_92),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_86),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_79),
.C(n_84),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_111),
.C(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_102),
.B1(n_103),
.B2(n_89),
.Y(n_113)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_110),
.B(n_80),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_87),
.C(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_107),
.B(n_110),
.C(n_97),
.D(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_103),
.B(n_121),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.C(n_116),
.Y(n_128)
);

OAI31xp33_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_115),
.A3(n_107),
.B(n_111),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_128),
.B(n_112),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_124),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_126),
.Y(n_131)
);


endmodule