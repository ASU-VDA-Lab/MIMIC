module fake_jpeg_8879_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_33),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_1),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_13),
.B1(n_25),
.B2(n_17),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_25),
.B1(n_44),
.B2(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_33),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_35),
.Y(n_56)
);

MAJx2_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_34),
.C(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_51),
.C(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_12),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_71),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_24),
.B(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_12),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_57),
.B1(n_49),
.B2(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_81),
.B1(n_68),
.B2(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_3),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_70),
.B(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_48),
.B1(n_59),
.B2(n_18),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_16),
.B(n_21),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_84),
.B(n_68),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_74),
.C(n_69),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.C(n_91),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_73),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_24),
.B(n_18),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_76),
.B1(n_85),
.B2(n_87),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_77),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_84),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_94),
.B(n_92),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_94),
.B(n_67),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_102),
.B(n_103),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_5),
.B(n_6),
.Y(n_106)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_6),
.B(n_9),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_109),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_108),
.Y(n_111)
);


endmodule