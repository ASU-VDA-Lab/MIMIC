module fake_jpeg_6181_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx10_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_12),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_16),
.B1(n_19),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_51),
.B1(n_53),
.B2(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_30),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_19),
.B1(n_30),
.B2(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_60),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_10),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_65),
.Y(n_98)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_64),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_32),
.C(n_36),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_30),
.B1(n_26),
.B2(n_16),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_47),
.B1(n_46),
.B2(n_29),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_23),
.B(n_36),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_31),
.B(n_36),
.C(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_81),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_46),
.B1(n_29),
.B2(n_24),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_40),
.C(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_44),
.B1(n_47),
.B2(n_55),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_92),
.B1(n_110),
.B2(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_47),
.B1(n_46),
.B2(n_22),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_76),
.B1(n_63),
.B2(n_22),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_114),
.B1(n_76),
.B2(n_31),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_59),
.B1(n_31),
.B2(n_36),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_59),
.B1(n_24),
.B2(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_138),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_61),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_66),
.B(n_64),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_120),
.A2(n_123),
.B(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_59),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_83),
.B1(n_75),
.B2(n_88),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_105),
.B1(n_89),
.B2(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_66),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_105),
.B(n_35),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_130),
.B1(n_97),
.B2(n_99),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_135),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_61),
.B(n_75),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_76),
.B1(n_67),
.B2(n_41),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_99),
.B1(n_98),
.B2(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_67),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_63),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_85),
.C(n_34),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_142),
.C(n_112),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_40),
.B(n_35),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_40),
.C(n_35),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_21),
.C(n_80),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.Y(n_174)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_153),
.Y(n_185)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_89),
.B1(n_106),
.B2(n_29),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_141),
.B(n_0),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_34),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_21),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_34),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_125),
.B(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_164),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_171),
.Y(n_187)
);

CKINVDCx10_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_131),
.B1(n_122),
.B2(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_81),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_117),
.Y(n_186)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_177),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_173),
.B(n_178),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_192),
.C(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_181),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_167),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_184),
.B1(n_144),
.B2(n_143),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_123),
.B1(n_125),
.B2(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_133),
.B1(n_140),
.B2(n_132),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_159),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_21),
.C(n_23),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_21),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_185),
.Y(n_203)
);

AO22x2_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_166),
.B1(n_157),
.B2(n_148),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_213),
.B1(n_176),
.B2(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_175),
.C(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_216),
.B1(n_210),
.B2(n_208),
.Y(n_224)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_166),
.B1(n_160),
.B2(n_150),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_156),
.C(n_147),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_200),
.C(n_207),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_161),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_204),
.B1(n_198),
.B2(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_230),
.C(n_231),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_225),
.B1(n_233),
.B2(n_211),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_196),
.B1(n_174),
.B2(n_177),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_213),
.B(n_156),
.Y(n_226)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_227),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_193),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_197),
.B(n_203),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_180),
.C(n_190),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_183),
.C(n_171),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_1),
.C(n_2),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_212),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_242),
.B1(n_4),
.B2(n_5),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_202),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_219),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_198),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_216),
.B(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_199),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_228),
.B1(n_232),
.B2(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_229),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_237),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_253),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_209),
.C(n_2),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.C(n_15),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_1),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_242),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_262),
.C(n_6),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_235),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.Y(n_269)
);

OAI321xp33_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_246),
.A3(n_249),
.B1(n_237),
.B2(n_235),
.C(n_12),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_261),
.A2(n_8),
.B(n_11),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_6),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

OAI21x1_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_259),
.B(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_13),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_269),
.C(n_14),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_271),
.C(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_13),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_278),
.B(n_15),
.Y(n_279)
);


endmodule