module real_aes_11691_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_1352;
wire n_394;
wire n_1280;
wire n_1323;
wire n_729;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_0), .A2(n_210), .B1(n_346), .B2(n_484), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_0), .A2(n_210), .B1(n_382), .B2(n_477), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_1), .A2(n_13), .B1(n_469), .B2(n_891), .Y(n_941) );
INVx1_ASAP7_75t_L g950 ( .A(n_1), .Y(n_950) );
INVx1_ASAP7_75t_L g468 ( .A(n_2), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_2), .A2(n_130), .B1(n_295), .B2(n_398), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_3), .A2(n_22), .B1(n_618), .B2(n_619), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_3), .A2(n_230), .B1(n_317), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_4), .A2(n_10), .B1(n_410), .B2(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g502 ( .A(n_4), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g1038 ( .A1(n_5), .A2(n_7), .B1(n_1033), .B2(n_1039), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_6), .A2(n_164), .B1(n_629), .B2(n_635), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_6), .A2(n_164), .B1(n_737), .B2(n_792), .Y(n_795) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_8), .Y(n_261) );
INVx1_ASAP7_75t_L g403 ( .A(n_8), .Y(n_403) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_8), .B(n_282), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_8), .B(n_184), .Y(n_1237) );
INVx1_ASAP7_75t_L g920 ( .A(n_9), .Y(n_920) );
INVx1_ASAP7_75t_L g504 ( .A(n_10), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_11), .A2(n_218), .B1(n_1022), .B2(n_1025), .Y(n_1043) );
AOI222xp33_ASAP7_75t_L g1212 ( .A1(n_11), .A2(n_1213), .B1(n_1311), .B2(n_1313), .C1(n_1357), .C2(n_1361), .Y(n_1212) );
XNOR2x2_ASAP7_75t_L g1213 ( .A(n_11), .B(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g807 ( .A(n_12), .Y(n_807) );
INVx1_ASAP7_75t_L g948 ( .A(n_13), .Y(n_948) );
INVx1_ASAP7_75t_L g1322 ( .A(n_14), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_15), .A2(n_36), .B1(n_784), .B2(n_1227), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_15), .A2(n_36), .B1(n_896), .B2(n_1350), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_16), .A2(n_193), .B1(n_295), .B2(n_382), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_16), .A2(n_193), .B1(n_406), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_17), .A2(n_237), .B1(n_424), .B2(n_572), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_17), .A2(n_237), .B1(n_629), .B2(n_635), .Y(n_694) );
INVxp33_ASAP7_75t_SL g862 ( .A(n_18), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_18), .A2(n_243), .B1(n_654), .B2(n_663), .Y(n_881) );
CKINVDCx14_ASAP7_75t_R g1047 ( .A(n_19), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_20), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_21), .Y(n_461) );
INVx1_ASAP7_75t_L g607 ( .A(n_22), .Y(n_607) );
INVx1_ASAP7_75t_L g466 ( .A(n_23), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_23), .A2(n_245), .B1(n_393), .B2(n_480), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g560 ( .A(n_24), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g330 ( .A(n_25), .Y(n_330) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_25), .B(n_1268), .Y(n_1304) );
INVxp33_ASAP7_75t_SL g817 ( .A(n_26), .Y(n_817) );
AOI22xp5_ASAP7_75t_SL g850 ( .A1(n_26), .A2(n_59), .B1(n_851), .B2(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g326 ( .A(n_27), .Y(n_326) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_27), .A2(n_198), .B1(n_398), .B2(n_399), .Y(n_397) );
BUFx2_ASAP7_75t_L g323 ( .A(n_28), .Y(n_323) );
BUFx2_ASAP7_75t_L g374 ( .A(n_28), .Y(n_374) );
INVx1_ASAP7_75t_L g674 ( .A(n_28), .Y(n_674) );
AO22x1_ASAP7_75t_L g799 ( .A1(n_29), .A2(n_800), .B1(n_801), .B2(n_855), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_29), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_30), .A2(n_100), .B1(n_424), .B2(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_L g549 ( .A(n_30), .Y(n_549) );
INVx1_ASAP7_75t_L g867 ( .A(n_31), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_31), .A2(n_70), .B1(n_875), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_32), .A2(n_199), .B1(n_821), .B2(n_875), .Y(n_927) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_32), .A2(n_199), .B1(n_469), .B2(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1325 ( .A(n_33), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_33), .A2(n_90), .B1(n_295), .B2(n_1342), .Y(n_1341) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_34), .A2(n_161), .B1(n_827), .B2(n_829), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_34), .A2(n_161), .B1(n_845), .B2(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g1327 ( .A(n_35), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_35), .A2(n_140), .B1(n_546), .B2(n_973), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_37), .A2(n_45), .B1(n_393), .B2(n_1345), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_37), .A2(n_45), .B1(n_489), .B2(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g626 ( .A(n_38), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_39), .A2(n_137), .B1(n_653), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_39), .A2(n_137), .B1(n_792), .B2(n_888), .Y(n_887) );
INVxp67_ASAP7_75t_L g975 ( .A(n_40), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_40), .A2(n_116), .B1(n_999), .B2(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_41), .A2(n_44), .B1(n_777), .B2(n_1224), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_41), .A2(n_63), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
OAI211xp5_ASAP7_75t_L g917 ( .A1(n_42), .A2(n_452), .B(n_733), .C(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g932 ( .A1(n_42), .A2(n_197), .B1(n_821), .B2(n_876), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_43), .A2(n_234), .B1(n_572), .B2(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_43), .A2(n_169), .B1(n_317), .B2(n_629), .Y(n_748) );
INVxp67_ASAP7_75t_SL g1305 ( .A(n_44), .Y(n_1305) );
XNOR2xp5_ASAP7_75t_L g753 ( .A(n_46), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g869 ( .A(n_47), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_47), .A2(n_208), .B1(n_500), .B2(n_546), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_48), .A2(n_168), .B1(n_924), .B2(n_925), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_48), .A2(n_168), .B1(n_899), .B2(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1254 ( .A(n_49), .Y(n_1254) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_50), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_51), .A2(n_212), .B1(n_533), .B2(n_534), .Y(n_532) );
INVxp33_ASAP7_75t_L g551 ( .A(n_51), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_52), .A2(n_124), .B1(n_836), .B2(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_52), .A2(n_124), .B1(n_469), .B2(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g820 ( .A(n_53), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_53), .A2(n_131), .B1(n_516), .B2(n_845), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_54), .A2(n_81), .B1(n_614), .B2(n_618), .Y(n_643) );
INVx1_ASAP7_75t_L g667 ( .A(n_54), .Y(n_667) );
INVx1_ASAP7_75t_L g720 ( .A(n_55), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_55), .A2(n_169), .B1(n_614), .B2(n_618), .Y(n_739) );
INVx1_ASAP7_75t_L g963 ( .A(n_56), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_56), .A2(n_75), .B1(n_821), .B2(n_982), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_57), .A2(n_226), .B1(n_616), .B2(n_619), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_57), .A2(n_226), .B1(n_661), .B2(n_663), .C(n_666), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_58), .A2(n_84), .B1(n_1033), .B2(n_1039), .Y(n_1044) );
INVxp33_ASAP7_75t_SL g818 ( .A(n_59), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_60), .A2(n_176), .B1(n_262), .B2(n_317), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_60), .A2(n_174), .B1(n_484), .B2(n_790), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_61), .A2(n_231), .B1(n_346), .B2(n_484), .Y(n_491) );
INVx1_ASAP7_75t_L g497 ( .A(n_61), .Y(n_497) );
AOI22xp5_ASAP7_75t_SL g1028 ( .A1(n_62), .A2(n_78), .B1(n_1029), .B2(n_1033), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_63), .A2(n_172), .B1(n_784), .B2(n_1227), .C(n_1229), .Y(n_1226) );
INVx1_ASAP7_75t_L g625 ( .A(n_64), .Y(n_625) );
INVx1_ASAP7_75t_L g960 ( .A(n_65), .Y(n_960) );
INVx1_ASAP7_75t_L g762 ( .A(n_66), .Y(n_762) );
INVx1_ASAP7_75t_L g578 ( .A(n_67), .Y(n_578) );
INVx1_ASAP7_75t_L g765 ( .A(n_68), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_68), .A2(n_113), .B1(n_393), .B2(n_782), .Y(n_781) );
CKINVDCx16_ASAP7_75t_R g1067 ( .A(n_69), .Y(n_1067) );
INVxp33_ASAP7_75t_SL g861 ( .A(n_70), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_71), .A2(n_241), .B1(n_379), .B2(n_380), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_71), .A2(n_241), .B1(n_410), .B2(n_411), .Y(n_409) );
INVxp67_ASAP7_75t_SL g1335 ( .A(n_72), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_72), .A2(n_136), .B1(n_851), .B2(n_999), .Y(n_1355) );
INVx1_ASAP7_75t_L g717 ( .A(n_73), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_73), .A2(n_155), .B1(n_616), .B2(n_619), .Y(n_746) );
INVx1_ASAP7_75t_L g583 ( .A(n_74), .Y(n_583) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_74), .A2(n_318), .B(n_631), .C(n_633), .Y(n_630) );
INVxp33_ASAP7_75t_SL g957 ( .A(n_75), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_76), .A2(n_205), .B1(n_394), .B2(n_663), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_76), .A2(n_205), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g814 ( .A(n_77), .Y(n_814) );
INVxp33_ASAP7_75t_SL g1320 ( .A(n_79), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_79), .A2(n_153), .B1(n_393), .B2(n_782), .Y(n_1340) );
AO22x2_ASAP7_75t_L g274 ( .A1(n_80), .A2(n_275), .B1(n_429), .B2(n_430), .Y(n_274) );
INVxp67_ASAP7_75t_L g429 ( .A(n_80), .Y(n_429) );
INVx1_ASAP7_75t_L g693 ( .A(n_81), .Y(n_693) );
INVx1_ASAP7_75t_L g518 ( .A(n_82), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_82), .A2(n_85), .B1(n_500), .B2(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g372 ( .A(n_83), .Y(n_372) );
INVx1_ASAP7_75t_L g1268 ( .A(n_83), .Y(n_1268) );
INVx1_ASAP7_75t_L g519 ( .A(n_85), .Y(n_519) );
INVx1_ASAP7_75t_L g735 ( .A(n_86), .Y(n_735) );
OAI211xp5_ASAP7_75t_SL g749 ( .A1(n_86), .A2(n_318), .B(n_631), .C(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g656 ( .A(n_87), .Y(n_656) );
INVx1_ASAP7_75t_L g570 ( .A(n_88), .Y(n_570) );
INVxp67_ASAP7_75t_SL g971 ( .A(n_89), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_89), .A2(n_122), .B1(n_406), .B2(n_992), .Y(n_997) );
INVxp33_ASAP7_75t_SL g1319 ( .A(n_90), .Y(n_1319) );
INVx1_ASAP7_75t_L g1256 ( .A(n_91), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g1275 ( .A1(n_91), .A2(n_233), .B1(n_1276), .B2(n_1278), .C(n_1279), .Y(n_1275) );
INVx1_ASAP7_75t_L g611 ( .A(n_92), .Y(n_611) );
INVx1_ASAP7_75t_L g472 ( .A(n_93), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_93), .A2(n_175), .B1(n_301), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g278 ( .A(n_94), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_94), .A2(n_206), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_95), .A2(n_219), .B1(n_1022), .B2(n_1081), .Y(n_1080) );
CKINVDCx20_ASAP7_75t_R g1090 ( .A(n_96), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_97), .A2(n_192), .B1(n_382), .B2(n_386), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_97), .A2(n_192), .B1(n_406), .B2(n_407), .Y(n_405) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_98), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_98), .A2(n_181), .B1(n_410), .B2(n_572), .Y(n_729) );
INVxp33_ASAP7_75t_SL g804 ( .A(n_99), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_99), .A2(n_246), .B1(n_827), .B2(n_836), .Y(n_835) );
INVxp33_ASAP7_75t_L g548 ( .A(n_100), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_101), .A2(n_214), .B1(n_898), .B2(n_899), .Y(n_897) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_101), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_102), .A2(n_209), .B1(n_379), .B2(n_380), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_102), .A2(n_209), .B1(n_487), .B2(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g582 ( .A(n_103), .Y(n_582) );
OAI22xp33_ASAP7_75t_SL g634 ( .A1(n_103), .A2(n_138), .B1(n_262), .B2(n_635), .Y(n_634) );
AO22x2_ASAP7_75t_L g508 ( .A1(n_104), .A2(n_509), .B1(n_554), .B2(n_555), .Y(n_508) );
INVx1_ASAP7_75t_L g554 ( .A(n_104), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_105), .A2(n_1314), .B1(n_1315), .B2(n_1356), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_105), .Y(n_1356) );
INVx1_ASAP7_75t_L g253 ( .A(n_106), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_107), .A2(n_160), .B1(n_898), .B2(n_943), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_107), .A2(n_160), .B1(n_629), .B2(n_635), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_108), .A2(n_194), .B1(n_653), .B2(n_654), .C(n_655), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_108), .A2(n_194), .B1(n_424), .B2(n_425), .Y(n_681) );
INVx1_ASAP7_75t_L g649 ( .A(n_109), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_110), .Y(n_315) );
INVx1_ASAP7_75t_L g811 ( .A(n_111), .Y(n_811) );
INVx1_ASAP7_75t_L g521 ( .A(n_112), .Y(n_521) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_113), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_114), .A2(n_236), .B1(n_894), .B2(n_896), .Y(n_893) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_114), .Y(n_904) );
XNOR2xp5_ASAP7_75t_L g912 ( .A(n_115), .B(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_115), .A2(n_202), .B1(n_1022), .B2(n_1025), .Y(n_1021) );
INVxp67_ASAP7_75t_L g976 ( .A(n_116), .Y(n_976) );
INVxp67_ASAP7_75t_SL g966 ( .A(n_117), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_117), .A2(n_247), .B1(n_546), .B2(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g1262 ( .A(n_118), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_119), .A2(n_120), .B1(n_1029), .B2(n_1083), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_121), .A2(n_126), .B1(n_425), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_121), .A2(n_126), .B1(n_379), .B2(n_380), .Y(n_540) );
INVxp67_ASAP7_75t_SL g969 ( .A(n_122), .Y(n_969) );
CKINVDCx14_ASAP7_75t_R g640 ( .A(n_123), .Y(n_640) );
XOR2xp5_ASAP7_75t_L g703 ( .A(n_125), .B(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g1037 ( .A1(n_125), .A2(n_147), .B1(n_1022), .B2(n_1025), .Y(n_1037) );
INVx1_ASAP7_75t_L g648 ( .A(n_127), .Y(n_648) );
INVx1_ASAP7_75t_L g864 ( .A(n_128), .Y(n_864) );
INVxp33_ASAP7_75t_SL g512 ( .A(n_129), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_129), .A2(n_141), .B1(n_477), .B2(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g465 ( .A(n_130), .Y(n_465) );
INVxp33_ASAP7_75t_SL g823 ( .A(n_131), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_132), .A2(n_221), .B1(n_618), .B2(n_619), .Y(n_916) );
INVxp33_ASAP7_75t_SL g951 ( .A(n_132), .Y(n_951) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_133), .A2(n_176), .B1(n_614), .B2(n_618), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_133), .A2(n_203), .B1(n_398), .B2(n_784), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_134), .A2(n_197), .B1(n_614), .B2(n_616), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_134), .A2(n_221), .B1(n_924), .B2(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g574 ( .A(n_135), .Y(n_574) );
INVxp33_ASAP7_75t_L g1334 ( .A(n_136), .Y(n_1334) );
INVx1_ASAP7_75t_L g586 ( .A(n_138), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_139), .A2(n_157), .B1(n_1231), .B2(n_1238), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1287 ( .A1(n_139), .A2(n_157), .B1(n_1288), .B2(n_1295), .C(n_1298), .Y(n_1287) );
INVx1_ASAP7_75t_L g1326 ( .A(n_140), .Y(n_1326) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_141), .Y(n_515) );
INVxp33_ASAP7_75t_SL g522 ( .A(n_142), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_142), .A2(n_165), .B1(n_379), .B2(n_380), .Y(n_528) );
INVxp33_ASAP7_75t_SL g958 ( .A(n_143), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_143), .A2(n_227), .B1(n_980), .B2(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g606 ( .A(n_144), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_144), .A2(n_163), .B1(n_614), .B2(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g710 ( .A(n_145), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_146), .A2(n_222), .B1(n_382), .B2(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_146), .A2(n_222), .B1(n_346), .B2(n_484), .Y(n_483) );
AO221x2_ASAP7_75t_L g1045 ( .A1(n_148), .A2(n_229), .B1(n_1033), .B2(n_1039), .C(n_1046), .Y(n_1045) );
CKINVDCx16_ASAP7_75t_R g1069 ( .A(n_149), .Y(n_1069) );
XNOR2xp5_ASAP7_75t_L g953 ( .A(n_150), .B(n_954), .Y(n_953) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_151), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_151), .B(n_253), .Y(n_1010) );
AND3x2_ASAP7_75t_L g1032 ( .A(n_151), .B(n_253), .C(n_1013), .Y(n_1032) );
AOI22xp5_ASAP7_75t_SL g1086 ( .A1(n_152), .A2(n_171), .B1(n_1029), .B2(n_1033), .Y(n_1086) );
INVxp33_ASAP7_75t_SL g1323 ( .A(n_153), .Y(n_1323) );
INVxp33_ASAP7_75t_SL g1337 ( .A(n_154), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_154), .A2(n_207), .B1(n_896), .B2(n_1350), .Y(n_1354) );
INVx1_ASAP7_75t_L g718 ( .A(n_155), .Y(n_718) );
INVx1_ASAP7_75t_L g761 ( .A(n_156), .Y(n_761) );
INVx2_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
AOI22xp5_ASAP7_75t_SL g1085 ( .A1(n_159), .A2(n_225), .B1(n_1022), .B2(n_1025), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_162), .A2(n_216), .B1(n_931), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_162), .A2(n_216), .B1(n_569), .B2(n_792), .Y(n_994) );
INVx1_ASAP7_75t_L g610 ( .A(n_163), .Y(n_610) );
INVxp33_ASAP7_75t_SL g513 ( .A(n_165), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_166), .A2(n_177), .B1(n_982), .B2(n_984), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_166), .A2(n_177), .B1(n_935), .B2(n_992), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_167), .A2(n_186), .B1(n_775), .B2(n_777), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_167), .A2(n_186), .B1(n_737), .B2(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g1013 ( .A(n_170), .Y(n_1013) );
INVxp67_ASAP7_75t_SL g1307 ( .A(n_172), .Y(n_1307) );
INVx1_ASAP7_75t_L g1253 ( .A(n_173), .Y(n_1253) );
OAI211xp5_ASAP7_75t_L g769 ( .A1(n_174), .A2(n_318), .B(n_631), .C(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g470 ( .A(n_175), .Y(n_470) );
INVx1_ASAP7_75t_L g361 ( .A(n_178), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_178), .A2(n_213), .B1(n_393), .B2(n_394), .Y(n_392) );
AO221x2_ASAP7_75t_L g1087 ( .A1(n_179), .A2(n_248), .B1(n_1083), .B2(n_1088), .C(n_1089), .Y(n_1087) );
OAI211xp5_ASAP7_75t_L g1216 ( .A1(n_180), .A2(n_1217), .B(n_1222), .C(n_1240), .Y(n_1216) );
AOI221xp5_ASAP7_75t_L g1280 ( .A1(n_180), .A2(n_190), .B1(n_1281), .B2(n_1283), .C(n_1284), .Y(n_1280) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_181), .Y(n_712) );
INVx1_ASAP7_75t_L g709 ( .A(n_182), .Y(n_709) );
INVx1_ASAP7_75t_L g685 ( .A(n_183), .Y(n_685) );
INVx1_ASAP7_75t_L g268 ( .A(n_184), .Y(n_268) );
INVx2_ASAP7_75t_L g282 ( .A(n_184), .Y(n_282) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_185), .A2(n_452), .B(n_645), .C(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g670 ( .A(n_185), .Y(n_670) );
XOR2x2_ASAP7_75t_L g857 ( .A(n_187), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g1241 ( .A(n_188), .Y(n_1241) );
CKINVDCx14_ASAP7_75t_R g1091 ( .A(n_189), .Y(n_1091) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_190), .A2(n_1248), .B1(n_1250), .B2(n_1255), .C(n_1258), .Y(n_1247) );
INVx1_ASAP7_75t_L g294 ( .A(n_191), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_191), .A2(n_239), .B1(n_419), .B2(n_421), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_191), .A2(n_318), .B(n_434), .C(n_439), .Y(n_433) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_195), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g658 ( .A(n_196), .Y(n_658) );
INVx1_ASAP7_75t_L g349 ( .A(n_198), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_198), .A2(n_447), .B(n_452), .C(n_453), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g1064 ( .A(n_200), .Y(n_1064) );
INVx1_ASAP7_75t_L g732 ( .A(n_201), .Y(n_732) );
OAI22xp33_ASAP7_75t_SL g751 ( .A1(n_201), .A2(n_234), .B1(n_262), .B2(n_635), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_203), .Y(n_758) );
INVxp33_ASAP7_75t_SL g808 ( .A(n_204), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_204), .A2(n_224), .B1(n_663), .B2(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
INVxp67_ASAP7_75t_SL g1331 ( .A(n_207), .Y(n_1331) );
INVx1_ASAP7_75t_L g870 ( .A(n_208), .Y(n_870) );
INVx1_ASAP7_75t_L g567 ( .A(n_211), .Y(n_567) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_212), .Y(n_544) );
INVx1_ASAP7_75t_L g338 ( .A(n_213), .Y(n_338) );
INVxp33_ASAP7_75t_SL g907 ( .A(n_214), .Y(n_907) );
INVx1_ASAP7_75t_L g919 ( .A(n_215), .Y(n_919) );
INVx1_ASAP7_75t_L g1014 ( .A(n_217), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_217), .B(n_1012), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_220), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_223), .Y(n_744) );
INVxp33_ASAP7_75t_SL g805 ( .A(n_224), .Y(n_805) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_227), .Y(n_961) );
INVx2_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
INVx1_ASAP7_75t_L g588 ( .A(n_230), .Y(n_588) );
INVx1_ASAP7_75t_L g506 ( .A(n_231), .Y(n_506) );
INVx1_ASAP7_75t_L g1243 ( .A(n_232), .Y(n_1243) );
AOI21xp33_ASAP7_75t_L g1257 ( .A1(n_233), .A2(n_597), .B(n_1227), .Y(n_1257) );
CKINVDCx20_ASAP7_75t_R g1061 ( .A(n_235), .Y(n_1061) );
INVxp33_ASAP7_75t_SL g910 ( .A(n_236), .Y(n_910) );
BUFx3_ASAP7_75t_L g335 ( .A(n_238), .Y(n_335) );
INVx1_ASAP7_75t_L g365 ( .A(n_238), .Y(n_365) );
INVx1_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
BUFx3_ASAP7_75t_L g337 ( .A(n_240), .Y(n_337) );
INVx1_ASAP7_75t_L g343 ( .A(n_240), .Y(n_343) );
INVx1_ASAP7_75t_L g686 ( .A(n_242), .Y(n_686) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_243), .Y(n_865) );
INVx1_ASAP7_75t_L g722 ( .A(n_244), .Y(n_722) );
INVx1_ASAP7_75t_L g462 ( .A(n_245), .Y(n_462) );
INVx1_ASAP7_75t_L g810 ( .A(n_246), .Y(n_810) );
INVxp67_ASAP7_75t_SL g965 ( .A(n_247), .Y(n_965) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_269), .B(n_1004), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
AND2x4_ASAP7_75t_L g1312 ( .A(n_251), .B(n_257), .Y(n_1312) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_SL g1360 ( .A(n_252), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_252), .B(n_254), .Y(n_1362) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_254), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x6_ASAP7_75t_L g322 ( .A(n_259), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g553 ( .A(n_259), .B(n_323), .Y(n_553) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g390 ( .A(n_260), .B(n_268), .Y(n_390) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g597 ( .A(n_261), .B(n_281), .Y(n_597) );
INVx8_ASAP7_75t_L g314 ( .A(n_262), .Y(n_314) );
OR2x6_ASAP7_75t_L g262 ( .A(n_263), .B(n_267), .Y(n_262) );
OR2x6_ASAP7_75t_L g317 ( .A(n_263), .B(n_280), .Y(n_317) );
INVx2_ASAP7_75t_SL g593 ( .A(n_263), .Y(n_593) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_263), .Y(n_657) );
INVx2_ASAP7_75t_SL g669 ( .A(n_263), .Y(n_669) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_263), .Y(n_708) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g284 ( .A(n_265), .Y(n_284) );
AND2x4_ASAP7_75t_L g291 ( .A(n_265), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
INVx1_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
AND2x2_ASAP7_75t_L g385 ( .A(n_265), .B(n_266), .Y(n_385) );
INVx1_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
INVx2_ASAP7_75t_L g292 ( .A(n_266), .Y(n_292) );
INVx1_ASAP7_75t_L g303 ( .A(n_266), .Y(n_303) );
INVx1_ASAP7_75t_L g438 ( .A(n_266), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_266), .B(n_284), .Y(n_601) );
AND2x4_ASAP7_75t_L g302 ( .A(n_267), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g500 ( .A(n_268), .B(n_307), .Y(n_500) );
OR2x2_ASAP7_75t_L g973 ( .A(n_268), .B(n_307), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_696), .Y(n_269) );
XOR2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_507), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AO22x2_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_455), .B2(n_456), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI221x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_321), .B1(n_324), .B2(n_369), .C(n_375), .Y(n_275) );
NAND4xp25_ASAP7_75t_L g276 ( .A(n_277), .B(n_293), .C(n_312), .D(n_318), .Y(n_276) );
INVx1_ASAP7_75t_L g443 ( .A(n_277), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B1(n_287), .B2(n_288), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_279), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_279), .A2(n_503), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_279), .A2(n_288), .B1(n_817), .B2(n_818), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_279), .A2(n_288), .B1(n_907), .B2(n_908), .Y(n_906) );
AOI22xp5_ASAP7_75t_SL g974 ( .A1(n_279), .A2(n_288), .B1(n_975), .B2(n_976), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_279), .A2(n_503), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
AND2x4_ASAP7_75t_L g288 ( .A(n_280), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g503 ( .A(n_280), .B(n_289), .Y(n_503) );
INVx1_ASAP7_75t_L g636 ( .A(n_280), .Y(n_636) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_283), .Y(n_379) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_283), .Y(n_393) );
BUFx2_ASAP7_75t_L g653 ( .A(n_283), .Y(n_653) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_283), .Y(n_665) );
INVx1_ASAP7_75t_L g776 ( .A(n_283), .Y(n_776) );
BUFx2_ASAP7_75t_L g924 ( .A(n_283), .Y(n_924) );
INVx1_ASAP7_75t_L g1225 ( .A(n_283), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_283), .B(n_1221), .Y(n_1242) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g1239 ( .A(n_284), .Y(n_1239) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx5_ASAP7_75t_SL g629 ( .A(n_288), .Y(n_629) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_290), .Y(n_834) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_291), .Y(n_380) );
INVx3_ASAP7_75t_L g396 ( .A(n_291), .Y(n_396) );
INVx1_ASAP7_75t_L g1246 ( .A(n_291), .Y(n_1246) );
AND2x4_ASAP7_75t_L g297 ( .A(n_292), .B(n_298), .Y(n_297) );
AOI222xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B1(n_299), .B2(n_300), .C1(n_304), .C2(n_305), .Y(n_293) );
HB1xp67_ASAP7_75t_L g1330 ( .A(n_295), .Y(n_1330) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g1218 ( .A(n_296), .B(n_1219), .Y(n_1218) );
BUFx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g319 ( .A(n_297), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g387 ( .A(n_297), .Y(n_387) );
BUFx3_ASAP7_75t_L g399 ( .A(n_297), .Y(n_399) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_297), .Y(n_477) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_297), .Y(n_786) );
BUFx2_ASAP7_75t_L g885 ( .A(n_297), .Y(n_885) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_299), .A2(n_304), .B1(n_345), .B2(n_349), .C1(n_350), .C2(n_357), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_299), .A2(n_304), .B1(n_440), .B2(n_442), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_299), .A2(n_304), .B1(n_351), .B2(n_357), .Y(n_453) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g441 ( .A(n_302), .Y(n_441) );
INVx2_ASAP7_75t_L g546 ( .A(n_302), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_302), .A2(n_442), .B1(n_625), .B2(n_626), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g690 ( .A1(n_302), .A2(n_442), .B1(n_648), .B2(n_649), .C1(n_686), .C2(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_302), .A2(n_442), .B1(n_744), .B2(n_745), .Y(n_750) );
AOI222xp33_ASAP7_75t_L g819 ( .A1(n_302), .A2(n_442), .B1(n_811), .B2(n_814), .C1(n_820), .C2(n_821), .Y(n_819) );
AOI222xp33_ASAP7_75t_L g947 ( .A1(n_302), .A2(n_305), .B1(n_786), .B2(n_919), .C1(n_920), .C2(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1233 ( .A(n_303), .Y(n_1233) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
AND2x4_ASAP7_75t_L g442 ( .A(n_306), .B(n_309), .Y(n_442) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g437 ( .A(n_308), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_308), .B(n_438), .Y(n_595) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g320 ( .A(n_310), .Y(n_320) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g402 ( .A(n_311), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g432 ( .A(n_312), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_315), .B2(n_316), .Y(n_312) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_314), .A2(n_316), .B1(n_461), .B2(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_314), .A2(n_521), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_314), .A2(n_316), .B1(n_685), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_314), .A2(n_552), .B1(n_807), .B2(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_314), .A2(n_316), .B1(n_864), .B2(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_314), .A2(n_316), .B1(n_950), .B2(n_951), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_314), .A2(n_552), .B1(n_960), .B2(n_969), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_314), .A2(n_552), .B1(n_1322), .B2(n_1337), .Y(n_1336) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_315), .A2(n_360), .B1(n_361), .B2(n_362), .Y(n_359) );
INVx4_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx5_ASAP7_75t_L g552 ( .A(n_317), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_318), .B(n_690), .C(n_692), .Y(n_689) );
NAND4xp25_ASAP7_75t_SL g815 ( .A(n_318), .B(n_816), .C(n_819), .D(n_822), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g946 ( .A(n_318), .B(n_947), .C(n_949), .Y(n_946) );
CKINVDCx11_ASAP7_75t_R g318 ( .A(n_319), .Y(n_318) );
AOI211xp5_ASAP7_75t_L g496 ( .A1(n_319), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
AOI211xp5_ASAP7_75t_L g543 ( .A1(n_319), .A2(n_498), .B(n_544), .C(n_545), .Y(n_543) );
AOI211xp5_ASAP7_75t_SL g903 ( .A1(n_319), .A2(n_386), .B(n_904), .C(n_905), .Y(n_903) );
AOI211xp5_ASAP7_75t_L g970 ( .A1(n_319), .A2(n_386), .B(n_971), .C(n_972), .Y(n_970) );
AOI211xp5_ASAP7_75t_L g1329 ( .A1(n_319), .A2(n_1330), .B(n_1331), .C(n_1332), .Y(n_1329) );
OAI31xp33_ASAP7_75t_L g431 ( .A1(n_321), .A2(n_432), .A3(n_433), .B(n_443), .Y(n_431) );
OAI31xp33_ASAP7_75t_SL g627 ( .A1(n_321), .A2(n_628), .A3(n_630), .B(n_634), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_321), .A2(n_689), .B(n_694), .Y(n_688) );
OAI31xp33_ASAP7_75t_SL g747 ( .A1(n_321), .A2(n_748), .A3(n_749), .B(n_751), .Y(n_747) );
OAI31xp33_ASAP7_75t_L g767 ( .A1(n_321), .A2(n_768), .A3(n_769), .B(n_771), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_321), .A2(n_370), .B1(n_802), .B2(n_815), .C(n_824), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g945 ( .A1(n_321), .A2(n_946), .B(n_952), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g1316 ( .A1(n_321), .A2(n_370), .B1(n_1317), .B2(n_1328), .C(n_1338), .Y(n_1316) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_322), .Y(n_321) );
AOI31xp33_ASAP7_75t_L g495 ( .A1(n_322), .A2(n_496), .A3(n_501), .B(n_505), .Y(n_495) );
AOI31xp33_ASAP7_75t_L g902 ( .A1(n_322), .A2(n_903), .A3(n_906), .B(n_909), .Y(n_902) );
AOI31xp33_ASAP7_75t_L g967 ( .A1(n_322), .A2(n_968), .A3(n_970), .B(n_974), .Y(n_967) );
AND2x4_ASAP7_75t_L g426 ( .A(n_323), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g683 ( .A(n_323), .B(n_427), .Y(n_683) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_323), .B(n_1265), .Y(n_1264) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_325), .B(n_344), .C(n_359), .D(n_366), .Y(n_324) );
INVxp67_ASAP7_75t_L g445 ( .A(n_325), .Y(n_445) );
AOI22xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B1(n_338), .B2(n_339), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_327), .A2(n_339), .B1(n_861), .B2(n_862), .Y(n_860) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
AND2x6_ASAP7_75t_L g362 ( .A(n_328), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g464 ( .A(n_328), .B(n_331), .Y(n_464) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g623 ( .A(n_329), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g341 ( .A(n_330), .Y(n_341) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
AND2x2_ASAP7_75t_L g416 ( .A(n_330), .B(n_372), .Y(n_416) );
INVx2_ASAP7_75t_L g428 ( .A(n_330), .Y(n_428) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_332), .Y(n_420) );
INVx2_ASAP7_75t_L g847 ( .A(n_332), .Y(n_847) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_332), .Y(n_892) );
INVx2_ASAP7_75t_L g895 ( .A(n_332), .Y(n_895) );
INVx6_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g360 ( .A(n_333), .B(n_352), .Y(n_360) );
BUFx2_ASAP7_75t_L g406 ( .A(n_333), .Y(n_406) );
INVx2_ASAP7_75t_L g485 ( .A(n_333), .Y(n_485) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_333), .B(n_1266), .Y(n_1265) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g358 ( .A(n_334), .Y(n_358) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g342 ( .A(n_335), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g348 ( .A(n_335), .B(n_337), .Y(n_348) );
INVx1_ASAP7_75t_L g356 ( .A(n_336), .Y(n_356) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g364 ( .A(n_337), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_339), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_339), .A2(n_464), .B1(n_512), .B2(n_513), .Y(n_511) );
CKINVDCx6p67_ASAP7_75t_R g616 ( .A(n_339), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_339), .A2(n_362), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_339), .A2(n_464), .B1(n_804), .B2(n_805), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_339), .A2(n_464), .B1(n_957), .B2(n_958), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_339), .A2(n_464), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
AND2x6_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
INVx1_ASAP7_75t_L g615 ( .A(n_340), .Y(n_615) );
AND2x2_ASAP7_75t_L g646 ( .A(n_340), .B(n_346), .Y(n_646) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x6_ASAP7_75t_L g357 ( .A(n_341), .B(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_342), .Y(n_410) );
BUFx3_ASAP7_75t_L g424 ( .A(n_342), .Y(n_424) );
INVx2_ASAP7_75t_SL g488 ( .A(n_342), .Y(n_488) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_342), .Y(n_526) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_342), .Y(n_569) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_342), .Y(n_737) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_342), .Y(n_1352) );
INVx1_ASAP7_75t_L g451 ( .A(n_343), .Y(n_451) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_346), .Y(n_868) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g367 ( .A(n_347), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g422 ( .A(n_347), .Y(n_422) );
INVx2_ASAP7_75t_L g535 ( .A(n_347), .Y(n_535) );
BUFx6f_ASAP7_75t_L g993 ( .A(n_347), .Y(n_993) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_348), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g866 ( .A1(n_350), .A2(n_357), .B1(n_867), .B2(n_868), .C1(n_869), .C2(n_870), .Y(n_866) );
BUFx4f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_351), .A2(n_357), .B1(n_648), .B2(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g813 ( .A(n_351), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g918 ( .A1(n_351), .A2(n_357), .B1(n_919), .B2(n_920), .Y(n_918) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_352), .B(n_354), .Y(n_471) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g624 ( .A(n_355), .Y(n_624) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g1292 ( .A(n_356), .Y(n_1292) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_357), .A2(n_468), .B1(n_469), .B2(n_470), .C1(n_471), .C2(n_472), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g514 ( .A1(n_357), .A2(n_471), .B1(n_515), .B2(n_516), .C1(n_518), .C2(n_519), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_357), .A2(n_611), .B1(n_622), .B2(n_623), .C1(n_625), .C2(n_626), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g741 ( .A1(n_357), .A2(n_623), .B1(n_722), .B2(n_742), .C1(n_744), .C2(n_745), .Y(n_741) );
AOI222xp33_ASAP7_75t_L g757 ( .A1(n_357), .A2(n_471), .B1(n_758), .B2(n_759), .C1(n_761), .C2(n_762), .Y(n_757) );
AOI222xp33_ASAP7_75t_L g809 ( .A1(n_357), .A2(n_469), .B1(n_810), .B2(n_811), .C1(n_812), .C2(n_814), .Y(n_809) );
AOI222xp33_ASAP7_75t_L g962 ( .A1(n_357), .A2(n_471), .B1(n_963), .B2(n_964), .C1(n_965), .C2(n_966), .Y(n_962) );
AOI222xp33_ASAP7_75t_L g1324 ( .A1(n_357), .A2(n_471), .B1(n_992), .B2(n_1325), .C1(n_1326), .C2(n_1327), .Y(n_1324) );
BUFx3_ASAP7_75t_L g1297 ( .A(n_358), .Y(n_1297) );
INVxp67_ASAP7_75t_L g454 ( .A(n_359), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_360), .A2(n_362), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_360), .A2(n_362), .B1(n_521), .B2(n_522), .Y(n_520) );
INVx4_ASAP7_75t_L g618 ( .A(n_360), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_360), .A2(n_362), .B1(n_807), .B2(n_808), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_360), .A2(n_362), .B1(n_864), .B2(n_865), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_360), .A2(n_362), .B1(n_960), .B2(n_961), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_360), .A2(n_362), .B1(n_1322), .B2(n_1323), .Y(n_1321) );
INVx4_ASAP7_75t_L g619 ( .A(n_362), .Y(n_619) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_363), .Y(n_425) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_363), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_363), .Y(n_494) );
INVx2_ASAP7_75t_L g587 ( .A(n_363), .Y(n_587) );
INVx1_ASAP7_75t_L g1001 ( .A(n_363), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g412 ( .A(n_364), .Y(n_412) );
INVx2_ASAP7_75t_L g539 ( .A(n_364), .Y(n_539) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_364), .Y(n_572) );
INVx1_ASAP7_75t_L g944 ( .A(n_364), .Y(n_944) );
INVx1_ASAP7_75t_L g450 ( .A(n_365), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_366), .B(n_460), .C(n_463), .D(n_467), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g802 ( .A(n_366), .B(n_803), .C(n_806), .D(n_809), .Y(n_802) );
NAND4xp25_ASAP7_75t_SL g859 ( .A(n_366), .B(n_860), .C(n_863), .D(n_866), .Y(n_859) );
INVx5_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
CKINVDCx8_ASAP7_75t_R g452 ( .A(n_367), .Y(n_452) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_369), .A2(n_445), .A3(n_446), .B(n_454), .Y(n_444) );
AOI211xp5_ASAP7_75t_SL g858 ( .A1(n_369), .A2(n_859), .B(n_871), .C(n_902), .Y(n_858) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AO211x2_ASAP7_75t_L g954 ( .A1(n_370), .A2(n_955), .B(n_967), .C(n_977), .Y(n_954) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x4_ASAP7_75t_L g458 ( .A(n_371), .B(n_373), .Y(n_458) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g427 ( .A(n_372), .B(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g389 ( .A(n_374), .Y(n_389) );
OR2x6_ASAP7_75t_L g596 ( .A(n_374), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_376), .B(n_431), .C(n_444), .Y(n_430) );
AND4x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_391), .C(n_404), .D(n_417), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .C(n_388), .Y(n_377) );
BUFx3_ASAP7_75t_L g654 ( .A(n_380), .Y(n_654) );
INVx2_ASAP7_75t_SL g662 ( .A(n_380), .Y(n_662) );
INVx2_ASAP7_75t_SL g880 ( .A(n_380), .Y(n_880) );
INVx4_ASAP7_75t_L g926 ( .A(n_380), .Y(n_926) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g530 ( .A(n_383), .Y(n_530) );
INVx2_ASAP7_75t_L g1342 ( .A(n_383), .Y(n_1342) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g398 ( .A(n_384), .Y(n_398) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_384), .Y(n_828) );
AND2x4_ASAP7_75t_L g1249 ( .A(n_384), .B(n_1221), .Y(n_1249) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g877 ( .A(n_385), .Y(n_877) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_388), .B(n_475), .C(n_476), .Y(n_474) );
AOI33xp33_ASAP7_75t_L g531 ( .A1(n_388), .A2(n_426), .A3(n_532), .B1(n_536), .B2(n_540), .B3(n_541), .Y(n_531) );
BUFx3_ASAP7_75t_L g659 ( .A(n_388), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_388), .B(n_774), .C(n_779), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g978 ( .A(n_388), .B(n_979), .C(n_981), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_388), .B(n_1344), .C(n_1347), .Y(n_1343) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
AND2x2_ASAP7_75t_L g400 ( .A(n_389), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g414 ( .A(n_389), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g564 ( .A(n_389), .B(n_565), .Y(n_564) );
OR2x6_ASAP7_75t_L g839 ( .A(n_389), .B(n_565), .Y(n_839) );
AND2x4_ASAP7_75t_L g873 ( .A(n_389), .B(n_390), .Y(n_873) );
BUFx2_ASAP7_75t_L g1260 ( .A(n_389), .Y(n_1260) );
INVx2_ASAP7_75t_L g1270 ( .A(n_389), .Y(n_1270) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .C(n_400), .Y(n_391) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_SL g480 ( .A(n_395), .Y(n_480) );
INVx2_ASAP7_75t_L g782 ( .A(n_395), .Y(n_782) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g603 ( .A(n_396), .Y(n_603) );
INVx3_ASAP7_75t_L g715 ( .A(n_396), .Y(n_715) );
BUFx2_ASAP7_75t_L g691 ( .A(n_399), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_400), .B(n_479), .C(n_481), .Y(n_478) );
AOI33xp33_ASAP7_75t_L g524 ( .A1(n_400), .A2(n_413), .A3(n_525), .B1(n_527), .B2(n_528), .B3(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g608 ( .A(n_400), .Y(n_608) );
INVx2_ASAP7_75t_SL g1229 ( .A(n_401), .Y(n_1229) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x6_ASAP7_75t_L g672 ( .A(n_402), .B(n_673), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .C(n_413), .Y(n_404) );
INVx1_ASAP7_75t_L g849 ( .A(n_407), .Y(n_849) );
INVx1_ASAP7_75t_L g1282 ( .A(n_407), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_407), .B(n_1299), .Y(n_1298) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx3_ASAP7_75t_L g469 ( .A(n_408), .Y(n_469) );
INVx1_ASAP7_75t_L g517 ( .A(n_408), .Y(n_517) );
INVx2_ASAP7_75t_SL g743 ( .A(n_408), .Y(n_743) );
INVx1_ASAP7_75t_L g760 ( .A(n_408), .Y(n_760) );
BUFx4f_ASAP7_75t_L g896 ( .A(n_408), .Y(n_896) );
INVx2_ASAP7_75t_L g938 ( .A(n_410), .Y(n_938) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_412), .B(n_1303), .Y(n_1309) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_413), .B(n_483), .C(n_486), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_413), .B(n_789), .C(n_791), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g1348 ( .A(n_413), .B(n_1349), .C(n_1351), .Y(n_1348) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_414), .A2(n_682), .B1(n_724), .B2(n_730), .Y(n_723) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g565 ( .A(n_416), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .C(n_426), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx4_ASAP7_75t_L g935 ( .A(n_420), .Y(n_935) );
INVx2_ASAP7_75t_L g1350 ( .A(n_420), .Y(n_1350) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g841 ( .A(n_424), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_426), .B(n_491), .C(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g589 ( .A(n_426), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_426), .B(n_794), .C(n_795), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g1353 ( .A(n_426), .B(n_1354), .C(n_1355), .Y(n_1353) );
AND2x4_ASAP7_75t_L g1266 ( .A(n_428), .B(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_436), .A2(n_592), .B1(n_610), .B2(n_611), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_436), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
OAI22xp33_ASAP7_75t_SL g666 ( .A1(n_436), .A2(n_667), .B1(n_668), .B2(n_670), .Y(n_666) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g632 ( .A(n_437), .Y(n_632) );
INVx2_ASAP7_75t_L g721 ( .A(n_437), .Y(n_721) );
INVx2_ASAP7_75t_L g1259 ( .A(n_437), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_440), .A2(n_442), .B1(n_761), .B2(n_762), .Y(n_770) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_449), .Y(n_580) );
INVx2_ASAP7_75t_L g680 ( .A(n_449), .Y(n_680) );
INVx1_ASAP7_75t_L g728 ( .A(n_449), .Y(n_728) );
BUFx2_ASAP7_75t_L g734 ( .A(n_449), .Y(n_734) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
OR2x2_ASAP7_75t_L g577 ( .A(n_450), .B(n_451), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_452), .B(n_511), .C(n_514), .D(n_520), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_452), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_452), .B(n_741), .Y(n_740) );
NAND3xp33_ASAP7_75t_SL g756 ( .A(n_452), .B(n_757), .C(n_763), .Y(n_756) );
NAND4xp25_ASAP7_75t_SL g955 ( .A(n_452), .B(n_956), .C(n_959), .D(n_962), .Y(n_955) );
NAND4xp25_ASAP7_75t_L g1317 ( .A(n_452), .B(n_1318), .C(n_1321), .D(n_1324), .Y(n_1317) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_473), .C(n_495), .Y(n_457) );
AOI211x1_ASAP7_75t_L g509 ( .A1(n_458), .A2(n_510), .B(n_523), .C(n_542), .Y(n_509) );
OAI31xp33_ASAP7_75t_L g612 ( .A1(n_458), .A2(n_613), .A3(n_617), .B(n_620), .Y(n_612) );
OAI31xp33_ASAP7_75t_L g642 ( .A1(n_458), .A2(n_643), .A3(n_644), .B(n_650), .Y(n_642) );
OAI31xp33_ASAP7_75t_SL g738 ( .A1(n_458), .A2(n_739), .A3(n_740), .B(n_746), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_458), .A2(n_756), .B(n_766), .Y(n_755) );
OAI31xp33_ASAP7_75t_L g914 ( .A1(n_458), .A2(n_915), .A3(n_916), .B(n_917), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .C(n_482), .D(n_490), .Y(n_473) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx2_ASAP7_75t_SL g830 ( .A(n_477), .Y(n_830) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g533 ( .A(n_485), .Y(n_533) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_487), .B(n_1302), .Y(n_1301) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g853 ( .A(n_488), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_488), .A2(n_1001), .B1(n_1253), .B2(n_1254), .Y(n_1279) );
INVx1_ASAP7_75t_L g843 ( .A(n_489), .Y(n_843) );
INVx1_ASAP7_75t_L g1286 ( .A(n_493), .Y(n_1286) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_556), .B1(n_557), .B2(n_695), .Y(n_507) );
INVx2_ASAP7_75t_L g695 ( .A(n_508), .Y(n_695) );
INVx1_ASAP7_75t_L g555 ( .A(n_509), .Y(n_555) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_531), .Y(n_523) );
INVx1_ASAP7_75t_L g585 ( .A(n_526), .Y(n_585) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_533), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_533), .B(n_1302), .Y(n_1306) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g622 ( .A(n_535), .Y(n_622) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g852 ( .A(n_538), .Y(n_852) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI31xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_547), .A3(n_550), .B(n_553), .Y(n_542) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
XNOR2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_638), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_612), .C(n_627), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_590), .Y(n_562) );
OAI33xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .A3(n_573), .B1(n_581), .B2(n_584), .B3(n_589), .Y(n_563) );
OAI22xp5_ASAP7_75t_SL g675 ( .A1(n_564), .A2(n_676), .B1(n_682), .B2(n_684), .Y(n_675) );
INVx1_ASAP7_75t_SL g939 ( .A(n_564), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_570), .B2(n_571), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_567), .A2(n_570), .B1(n_599), .B2(n_602), .Y(n_598) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx4f_ASAP7_75t_L g999 ( .A(n_569), .Y(n_999) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_572), .Y(n_792) );
INVx1_ASAP7_75t_L g900 ( .A(n_572), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_578), .B2(n_579), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_574), .A2(n_578), .B1(n_592), .B2(n_594), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_575), .A2(n_579), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g614 ( .A(n_577), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g678 ( .A(n_577), .Y(n_678) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_584) );
OAI33xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_596), .A3(n_598), .B1(n_604), .B2(n_608), .B3(n_609), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_594), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI33xp33_ASAP7_75t_L g706 ( .A1(n_596), .A2(n_608), .A3(n_707), .B1(n_711), .B2(n_716), .B3(n_719), .Y(n_706) );
OAI22xp33_ASAP7_75t_SL g711 ( .A1(n_599), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_599), .A2(n_602), .B1(n_717), .B2(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g605 ( .A(n_600), .Y(n_605) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_600), .Y(n_1252) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx2_ASAP7_75t_L g637 ( .A(n_601), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_602), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_602), .A2(n_1251), .B1(n_1253), .B2(n_1254), .Y(n_1250) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx3_ASAP7_75t_L g931 ( .A(n_603), .Y(n_931) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_640), .A2(n_1009), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
NAND3x1_ASAP7_75t_SL g641 ( .A(n_642), .B(n_651), .C(n_688), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_659), .B1(n_660), .B2(n_671), .C(n_675), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_656), .A2(n_658), .B1(n_677), .B2(n_679), .C(n_681), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_657), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
AOI33xp33_ASAP7_75t_L g825 ( .A1(n_659), .A2(n_671), .A3(n_826), .B1(n_831), .B2(n_832), .B3(n_835), .Y(n_825) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI33xp33_ASAP7_75t_L g872 ( .A1(n_671), .A2(n_873), .A3(n_874), .B1(n_878), .B2(n_881), .B3(n_882), .Y(n_872) );
INVx6_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx5_ASAP7_75t_L g787 ( .A(n_672), .Y(n_787) );
NAND2x1p5_ASAP7_75t_L g1294 ( .A(n_673), .B(n_1266), .Y(n_1294) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_674), .B(n_1304), .Y(n_1303) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_677), .A2(n_679), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_684) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g725 ( .A(n_678), .Y(n_725) );
INVx2_ASAP7_75t_L g731 ( .A(n_678), .Y(n_731) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x6_ASAP7_75t_L g1310 ( .A(n_680), .B(n_1303), .Y(n_1310) );
INVx4_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI33xp33_ASAP7_75t_L g837 ( .A1(n_683), .A2(n_838), .A3(n_840), .B1(n_844), .B2(n_850), .B3(n_854), .Y(n_837) );
BUFx4f_ASAP7_75t_L g901 ( .A(n_683), .Y(n_901) );
BUFx4f_ASAP7_75t_L g1002 ( .A(n_683), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1274 ( .A1(n_683), .A2(n_995), .B1(n_1275), .B2(n_1280), .C(n_1287), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_911), .B2(n_1003), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_797), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_752), .B2(n_796), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_738), .C(n_747), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_723), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_709), .A2(n_710), .B1(n_725), .B2(n_726), .C(n_729), .Y(n_724) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g778 ( .A(n_715), .Y(n_778) );
INVx2_ASAP7_75t_L g988 ( .A(n_715), .Y(n_988) );
OAI21xp5_ASAP7_75t_SL g1255 ( .A1(n_721), .A2(n_1256), .B(n_1257), .Y(n_1255) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_730) );
INVx2_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g889 ( .A(n_737), .Y(n_889) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g790 ( .A(n_743), .Y(n_790) );
INVx1_ASAP7_75t_L g796 ( .A(n_752), .Y(n_796) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND3x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_767), .C(n_772), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AND4x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_780), .C(n_788), .D(n_793), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g980 ( .A(n_776), .Y(n_980) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .C(n_787), .Y(n_780) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g821 ( .A(n_785), .Y(n_821) );
INVx2_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
BUFx2_ASAP7_75t_L g984 ( .A(n_786), .Y(n_984) );
NAND3xp33_ASAP7_75t_L g929 ( .A(n_787), .B(n_930), .C(n_932), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g985 ( .A(n_787), .B(n_986), .C(n_989), .Y(n_985) );
NAND3xp33_ASAP7_75t_L g1339 ( .A(n_787), .B(n_1340), .C(n_1341), .Y(n_1339) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_856), .B2(n_857), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g855 ( .A(n_801), .Y(n_855) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_837), .Y(n_824) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_SL g836 ( .A(n_830), .Y(n_836) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
AOI33xp33_ASAP7_75t_L g886 ( .A1(n_838), .A2(n_887), .A3(n_890), .B1(n_893), .B2(n_897), .B3(n_901), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g995 ( .A(n_839), .Y(n_995) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g964 ( .A(n_849), .Y(n_964) );
INVx2_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_886), .Y(n_871) );
BUFx2_ASAP7_75t_L g928 ( .A(n_873), .Y(n_928) );
BUFx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_SL g983 ( .A(n_877), .Y(n_983) );
INVx2_ASAP7_75t_SL g1273 ( .A(n_877), .Y(n_1273) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_SL g898 ( .A(n_889), .Y(n_898) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
BUFx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
HB1xp67_ASAP7_75t_L g1278 ( .A(n_895), .Y(n_1278) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g940 ( .A(n_901), .B(n_941), .C(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g1003 ( .A(n_911), .Y(n_1003) );
XOR2x2_ASAP7_75t_L g911 ( .A(n_912), .B(n_953), .Y(n_911) );
NAND3x1_ASAP7_75t_L g913 ( .A(n_914), .B(n_921), .C(n_945), .Y(n_913) );
AND4x1_ASAP7_75t_L g921 ( .A(n_922), .B(n_929), .C(n_933), .D(n_940), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_927), .C(n_928), .Y(n_922) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
NAND3xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_936), .C(n_939), .Y(n_933) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NAND4xp25_ASAP7_75t_L g977 ( .A(n_978), .B(n_985), .C(n_990), .D(n_996), .Y(n_977) );
BUFx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g1228 ( .A(n_983), .Y(n_1228) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_991), .B(n_994), .C(n_995), .Y(n_990) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1277 ( .A(n_993), .Y(n_1277) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .C(n_1002), .Y(n_996) );
INVx1_ASAP7_75t_L g1285 ( .A(n_999), .Y(n_1285) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI21xp33_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1015), .B(n_1212), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_1007), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1089) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_1008), .A2(n_1061), .B1(n_1062), .B2(n_1064), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1010), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_1010), .B(n_1027), .Y(n_1048) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1011), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1014), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1014), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1093), .B1(n_1156), .B2(n_1157), .C(n_1185), .Y(n_1015) );
A2O1A1Ixp33_ASAP7_75t_SL g1016 ( .A1(n_1017), .A2(n_1049), .B(n_1076), .C(n_1087), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1034), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1019), .B(n_1106), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1019), .B(n_1074), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1019), .B(n_1114), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1019), .B(n_1166), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1019), .B(n_1135), .Y(n_1200) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_1020), .B(n_1054), .Y(n_1053) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1020), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1020), .B(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1020), .B(n_1124), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1020), .B(n_1055), .Y(n_1128) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1020), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1020), .B(n_1035), .Y(n_1181) );
AOI211xp5_ASAP7_75t_L g1188 ( .A1(n_1020), .A2(n_1100), .B(n_1189), .C(n_1190), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1020), .B(n_1131), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1028), .Y(n_1020) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
OAI21xp33_ASAP7_75t_SL g1361 ( .A1(n_1023), .A2(n_1360), .B(n_1362), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_1024), .B(n_1026), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_1025), .Y(n_1081) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1029), .Y(n_1066) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_1029), .Y(n_1088) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1032), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1030), .B(n_1032), .Y(n_1039) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_1031), .B(n_1032), .Y(n_1033) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1033), .Y(n_1068) );
O2A1O1Ixp33_ASAP7_75t_L g1175 ( .A1(n_1034), .A2(n_1138), .B(n_1176), .C(n_1179), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1040), .Y(n_1034) );
NOR2x1_ASAP7_75t_L g1100 ( .A(n_1035), .B(n_1075), .Y(n_1100) );
AOI21xp5_ASAP7_75t_L g1129 ( .A1(n_1035), .A2(n_1130), .B(n_1133), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1135 ( .A(n_1035), .B(n_1041), .Y(n_1135) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_1036), .Y(n_1054) );
INVxp67_ASAP7_75t_L g1098 ( .A(n_1036), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1036), .B(n_1142), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1040), .B(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1040), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1045), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_1041), .A2(n_1159), .B1(n_1163), .B2(n_1165), .Y(n_1158) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1042), .B(n_1045), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1042), .B(n_1075), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1042), .B(n_1054), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1042), .B(n_1045), .Y(n_1143) );
NOR2xp33_ASAP7_75t_L g1207 ( .A(n_1042), .B(n_1054), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1045), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1045), .B(n_1054), .Y(n_1124) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1048), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1056), .B(n_1070), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1055), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1053), .B(n_1143), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1054), .B(n_1074), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1054), .B(n_1148), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1054), .B(n_1149), .Y(n_1189) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1055), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1055), .B(n_1181), .Y(n_1180) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1057), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_1057), .A2(n_1119), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1057), .B(n_1071), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1057), .B(n_1193), .Y(n_1192) );
INVx2_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1119 ( .A(n_1058), .B(n_1115), .Y(n_1119) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1058), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1140 ( .A(n_1058), .B(n_1141), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1058), .B(n_1110), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1058), .B(n_1084), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_1058), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_1059), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1059), .B(n_1084), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1059), .B(n_1115), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1065), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1062), .Y(n_1092) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1067), .B1(n_1068), .B2(n_1069), .Y(n_1065) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1068), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1071), .B(n_1113), .Y(n_1112) );
O2A1O1Ixp33_ASAP7_75t_L g1116 ( .A1(n_1071), .A2(n_1075), .B(n_1117), .C(n_1118), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1071), .B(n_1142), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1071), .B(n_1119), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1071), .B(n_1124), .Y(n_1184) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1073), .B(n_1141), .Y(n_1198) );
OAI21xp5_ASAP7_75t_L g1204 ( .A1(n_1073), .A2(n_1132), .B(n_1184), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1074), .B(n_1098), .Y(n_1122) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1074), .Y(n_1161) );
OAI32xp33_ASAP7_75t_L g1107 ( .A1(n_1075), .A2(n_1108), .A3(n_1109), .B1(n_1111), .B2(n_1114), .Y(n_1107) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1084), .Y(n_1077) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1078), .Y(n_1104) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1078), .Y(n_1110) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1079), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1079), .B(n_1084), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1079), .B(n_1115), .Y(n_1178) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1079), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1082), .Y(n_1079) );
INVx3_ASAP7_75t_L g1115 ( .A(n_1084), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1087), .Y(n_1144) );
OAI21xp5_ASAP7_75t_L g1195 ( .A1(n_1087), .A2(n_1166), .B(n_1196), .Y(n_1195) );
NAND5xp2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1099), .C(n_1120), .D(n_1129), .E(n_1145), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1096), .Y(n_1094) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1097), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1098), .B(n_1128), .Y(n_1127) );
AOI211xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1101), .B(n_1107), .C(n_1116), .Y(n_1099) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1102), .B(n_1147), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1105), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1104), .Y(n_1137) );
O2A1O1Ixp33_ASAP7_75t_L g1191 ( .A1(n_1104), .A2(n_1127), .B(n_1192), .C(n_1194), .Y(n_1191) );
OAI22xp5_ASAP7_75t_SL g1152 ( .A1(n_1105), .A2(n_1153), .B1(n_1154), .B2(n_1155), .Y(n_1152) );
A2O1A1Ixp33_ASAP7_75t_L g1179 ( .A1(n_1105), .A2(n_1180), .B(n_1182), .C(n_1183), .Y(n_1179) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1105), .A2(n_1174), .B(n_1203), .C(n_1204), .Y(n_1202) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_1106), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_1109), .A2(n_1121), .B1(n_1125), .B2(n_1127), .Y(n_1120) );
OAI211xp5_ASAP7_75t_SL g1157 ( .A1(n_1109), .A2(n_1158), .B(n_1167), .C(n_1175), .Y(n_1157) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1110), .B(n_1119), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1110), .B(n_1126), .Y(n_1196) );
OAI322xp33_ASAP7_75t_L g1205 ( .A1(n_1111), .A2(n_1118), .A3(n_1154), .B1(n_1155), .B2(n_1206), .C1(n_1208), .C2(n_1210), .Y(n_1205) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1113), .Y(n_1154) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
NAND3xp33_ASAP7_75t_L g1139 ( .A(n_1115), .B(n_1140), .C(n_1142), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1115), .B(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1122), .Y(n_1169) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1126), .B(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1130), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1132), .Y(n_1130) );
OAI211xp5_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1136), .B(n_1139), .C(n_1144), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1138), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1142), .B(n_1181), .Y(n_1193) );
NOR2xp33_ASAP7_75t_SL g1206 ( .A(n_1142), .B(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1144), .Y(n_1156) );
O2A1O1Ixp33_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1149), .B(n_1150), .C(n_1152), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
OAI21xp5_ASAP7_75t_L g1199 ( .A1(n_1149), .A2(n_1190), .B(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
O2A1O1Ixp33_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1169), .B(n_1170), .C(n_1172), .Y(n_1167) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1168), .Y(n_1182) );
OAI21xp5_ASAP7_75t_L g1183 ( .A1(n_1169), .A2(n_1178), .B(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
OAI211xp5_ASAP7_75t_SL g1185 ( .A1(n_1186), .A2(n_1188), .B(n_1191), .C(n_1201), .Y(n_1185) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1193), .Y(n_1203) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1197), .B(n_1199), .Y(n_1194) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
NOR3xp33_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1205), .C(n_1211), .Y(n_1201) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
NAND4xp25_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1261), .C(n_1274), .D(n_1300), .Y(n_1214) );
OAI21xp5_ASAP7_75t_SL g1215 ( .A1(n_1216), .A2(n_1247), .B(n_1260), .Y(n_1215) );
INVx8_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x4_ASAP7_75t_L g1244 ( .A(n_1219), .B(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
AOI21xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1226), .B(n_1230), .Y(n_1222) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
NAND2x1p5_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1234), .Y(n_1231) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
OR2x6_ASAP7_75t_L g1238 ( .A(n_1235), .B(n_1239), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1235), .B(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1235), .Y(n_1272) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_1241), .A2(n_1242), .B1(n_1243), .B2(n_1244), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_1241), .A2(n_1243), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1245), .Y(n_1346) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
CKINVDCx6p67_ASAP7_75t_R g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1263), .Y(n_1261) );
OR2x6_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1269), .Y(n_1263) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
NOR2xp67_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1271), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1273), .Y(n_1271) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
NAND2x1p5_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1293), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_SL g1293 ( .A(n_1294), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1294), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1294), .Y(n_1299) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1305), .B1(n_1306), .B2(n_1307), .C(n_1308), .Y(n_1300) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1333), .C(n_1336), .Y(n_1328) );
NAND4xp25_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1343), .C(n_1348), .D(n_1353), .Y(n_1338) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_1359), .Y(n_1358) );
endmodule