module fake_jpeg_9102_n_101 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_28),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_37),
.B(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_38),
.B1(n_40),
.B2(n_8),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_3),
.Y(n_71)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_14),
.B1(n_16),
.B2(n_19),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_86),
.B1(n_87),
.B2(n_68),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.A3(n_63),
.B1(n_79),
.B2(n_85),
.C1(n_80),
.C2(n_65),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_78),
.B1(n_79),
.B2(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_73),
.C(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_83),
.C(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_20),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_23),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_31),
.B(n_33),
.Y(n_101)
);


endmodule