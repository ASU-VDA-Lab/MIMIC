module fake_jpeg_615_n_389 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_9),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_55),
.B(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_57),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_63),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_69),
.Y(n_124)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_8),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_73),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_80),
.Y(n_130)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_31),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_32),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_89),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_12),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_15),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_15),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_98),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_16),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_33),
.B(n_13),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_14),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_54),
.B1(n_50),
.B2(n_45),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_37),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_52),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_39),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_26),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

BUFx2_ASAP7_75t_R g175 ( 
.A(n_110),
.Y(n_175)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_114),
.A2(n_144),
.B1(n_172),
.B2(n_164),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_116),
.A2(n_120),
.B1(n_155),
.B2(n_156),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_40),
.B1(n_46),
.B2(n_44),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_118),
.B(n_135),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_132),
.B1(n_137),
.B2(n_178),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_59),
.B1(n_66),
.B2(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_125),
.B(n_161),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_70),
.A2(n_43),
.B1(n_41),
.B2(n_54),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_41),
.B1(n_45),
.B2(n_50),
.Y(n_137)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_29),
.B1(n_26),
.B2(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_13),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_68),
.B(n_14),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_0),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_87),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_91),
.B(n_0),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_170),
.B(n_173),
.Y(n_214)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_2),
.Y(n_173)
);

CKINVDCx12_ASAP7_75t_R g177 ( 
.A(n_78),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g237 ( 
.A(n_177),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_94),
.A2(n_26),
.B1(n_42),
.B2(n_49),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_93),
.A2(n_42),
.B1(n_49),
.B2(n_3),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_60),
.B1(n_92),
.B2(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_184),
.B(n_192),
.Y(n_272)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_185),
.Y(n_279)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_140),
.A2(n_97),
.B1(n_96),
.B2(n_110),
.Y(n_186)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_62),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_194),
.Y(n_255)
);

BUFx2_ASAP7_75t_SL g191 ( 
.A(n_113),
.Y(n_191)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_90),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_126),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_193),
.B(n_209),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_111),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_132),
.B(n_178),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_195),
.A2(n_204),
.B(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_99),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_196),
.B(n_218),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_201),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_110),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_212),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_130),
.A2(n_82),
.B(n_84),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_120),
.A2(n_119),
.B1(n_134),
.B2(n_164),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_221),
.B1(n_225),
.B2(n_233),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_210),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_213),
.A2(n_227),
.B1(n_185),
.B2(n_235),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_215),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_149),
.B(n_4),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_217),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_49),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_58),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_219),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_220),
.A2(n_228),
.B1(n_230),
.B2(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_124),
.B(n_121),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_143),
.B(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_148),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_216),
.C(n_211),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_129),
.A2(n_139),
.B(n_147),
.C(n_180),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_231),
.B(n_186),
.C(n_237),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_148),
.B(n_174),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_231),
.Y(n_265)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_R g231 ( 
.A(n_129),
.B(n_121),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_127),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_133),
.A2(n_166),
.B1(n_157),
.B2(n_135),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_225),
.B1(n_198),
.B2(n_227),
.Y(n_247)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_226),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_128),
.B(n_160),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_237),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_165),
.A2(n_128),
.B1(n_160),
.B2(n_115),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_122),
.B1(n_165),
.B2(n_115),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_240),
.A2(n_251),
.B1(n_256),
.B2(n_260),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_165),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_278),
.C(n_280),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_247),
.A2(n_249),
.B1(n_265),
.B2(n_264),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_197),
.B1(n_196),
.B2(n_214),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_190),
.A2(n_208),
.B1(n_222),
.B2(n_182),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_242),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_208),
.A2(n_186),
.B1(n_189),
.B2(n_202),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_269),
.B(n_255),
.Y(n_291)
);

AO21x1_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_265),
.B(n_275),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_204),
.A2(n_208),
.B(n_183),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_208),
.A2(n_199),
.B1(n_230),
.B2(n_207),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_273),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_207),
.A2(n_212),
.B1(n_224),
.B2(n_228),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_224),
.A2(n_223),
.B1(n_206),
.B2(n_203),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_273),
.Y(n_305)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_200),
.B(n_220),
.C(n_232),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_188),
.B(n_194),
.C(n_218),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_245),
.A2(n_187),
.B1(n_249),
.B2(n_258),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_289),
.B1(n_300),
.B2(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_187),
.C(n_243),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_299),
.C(n_301),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_285),
.B(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_286),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_287),
.A2(n_296),
.B1(n_262),
.B2(n_268),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_272),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_288),
.B(n_290),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_245),
.A2(n_258),
.B1(n_251),
.B2(n_255),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_272),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_291),
.A2(n_299),
.B(n_292),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_248),
.B(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_260),
.B1(n_259),
.B2(n_263),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_248),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_259),
.C(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_253),
.B1(n_240),
.B2(n_244),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_278),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_274),
.B(n_241),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_303),
.C(n_281),
.Y(n_330)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_310),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_244),
.A2(n_270),
.B1(n_241),
.B2(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_252),
.B(n_242),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_252),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_254),
.Y(n_311)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_309),
.B(n_286),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_313),
.A2(n_318),
.B1(n_329),
.B2(n_300),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_254),
.A3(n_262),
.B1(n_268),
.B2(n_279),
.C1(n_310),
.C2(n_289),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_316),
.B(n_306),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_309),
.A2(n_283),
.B(n_285),
.Y(n_322)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_330),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_294),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_292),
.A2(n_297),
.B1(n_283),
.B2(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_281),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_336),
.C(n_339),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_284),
.C(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_303),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_302),
.C(n_282),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_341),
.C(n_322),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_297),
.C(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_345),
.C(n_347),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_321),
.B(n_307),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_324),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_317),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_333),
.A2(n_329),
.B1(n_312),
.B2(n_335),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_349),
.A2(n_313),
.B1(n_331),
.B2(n_332),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_335),
.A2(n_312),
.B1(n_320),
.B2(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_317),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_351),
.B(n_355),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_326),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_356),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_334),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_320),
.B1(n_323),
.B2(n_332),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_359),
.A2(n_350),
.B1(n_352),
.B2(n_357),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_364),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_352),
.A2(n_331),
.B(n_318),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_365),
.A2(n_359),
.B(n_356),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_338),
.B1(n_327),
.B2(n_337),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_368),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_367),
.A2(n_348),
.B1(n_339),
.B2(n_336),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_366),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_348),
.B1(n_363),
.B2(n_353),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_358),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_375),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_324),
.Y(n_375)
);

AOI31xp67_ASAP7_75t_SL g376 ( 
.A1(n_364),
.A2(n_353),
.A3(n_360),
.B(n_354),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_376),
.B(n_365),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_374),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_377),
.A2(n_380),
.B1(n_362),
.B2(n_361),
.Y(n_382)
);

AOI21xp33_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_381),
.B(n_371),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_383),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_379),
.A2(n_367),
.B(n_372),
.Y(n_383)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_384),
.Y(n_385)
);

AOI321xp33_ASAP7_75t_SL g387 ( 
.A1(n_385),
.A2(n_377),
.A3(n_370),
.B1(n_361),
.B2(n_362),
.C(n_354),
.Y(n_387)
);

OAI321xp33_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_360),
.A3(n_342),
.B1(n_328),
.B2(n_319),
.C(n_386),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_319),
.Y(n_389)
);


endmodule