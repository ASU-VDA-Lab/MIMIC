module real_aes_6834_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_792;
wire n_386;
wire n_905;
wire n_503;
wire n_518;
wire n_673;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_1123;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_744;
wire n_384;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_976;
wire n_466;
wire n_636;
wire n_872;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_780;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_1025;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_725;
wire n_455;
wire n_504;
wire n_973;
wire n_671;
wire n_1081;
wire n_960;
wire n_1084;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_817;
wire n_565;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_703;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_1006;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_1136;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_1033;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_831;
wire n_487;
wire n_653;
wire n_637;
wire n_526;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_717;
wire n_982;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_1114;
wire n_465;
wire n_566;
wire n_473;
wire n_837;
wire n_967;
wire n_871;
wire n_1045;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_1040;
wire n_393;
wire n_1097;
wire n_652;
wire n_500;
wire n_1101;
wire n_1102;
wire n_601;
wire n_463;
wire n_661;
wire n_396;
wire n_804;
wire n_1076;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_0), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_1), .A2(n_300), .B1(n_559), .B2(n_561), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_2), .A2(n_163), .B1(n_443), .B2(n_446), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_3), .A2(n_166), .B1(n_528), .B2(n_530), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_4), .Y(n_966) );
INVx1_ASAP7_75t_L g418 ( .A(n_5), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_6), .A2(n_349), .B1(n_524), .B2(n_610), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_7), .A2(n_131), .B1(n_446), .B2(n_659), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_8), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_9), .A2(n_103), .B1(n_596), .B2(n_597), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_10), .A2(n_139), .B1(n_468), .B2(n_523), .Y(n_1129) );
AO22x2_ASAP7_75t_L g407 ( .A1(n_11), .A2(n_223), .B1(n_408), .B2(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g1073 ( .A(n_11), .Y(n_1073) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_12), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_13), .A2(n_150), .B1(n_572), .B2(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g880 ( .A1(n_14), .A2(n_325), .B1(n_334), .B2(n_548), .C1(n_583), .C2(n_706), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_15), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_16), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_17), .A2(n_216), .B1(n_597), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_18), .A2(n_50), .B1(n_475), .B2(n_478), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_19), .A2(n_118), .B1(n_723), .B2(n_898), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_20), .A2(n_291), .B1(n_548), .B2(n_706), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_21), .A2(n_246), .B1(n_571), .B2(n_573), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_22), .A2(n_255), .B1(n_559), .B2(n_635), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_23), .B(n_977), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_24), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_25), .A2(n_263), .B1(n_573), .B2(n_718), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_26), .A2(n_361), .B1(n_461), .B2(n_889), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_27), .A2(n_95), .B1(n_548), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_28), .A2(n_204), .B1(n_571), .B2(n_573), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_29), .A2(n_192), .B1(n_420), .B2(n_426), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_30), .A2(n_317), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_31), .A2(n_157), .B1(n_602), .B2(n_785), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_32), .A2(n_321), .B1(n_478), .B2(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_33), .A2(n_136), .B1(n_600), .B2(n_603), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_34), .A2(n_85), .B1(n_664), .B2(n_992), .Y(n_1046) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_35), .A2(n_117), .B1(n_408), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_36), .A2(n_270), .B1(n_468), .B2(n_572), .Y(n_680) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_37), .A2(n_189), .B1(n_303), .B2(n_404), .C1(n_426), .C2(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_38), .B(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_39), .A2(n_76), .B1(n_468), .B2(n_751), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_40), .A2(n_262), .B1(n_602), .B2(n_722), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_41), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_42), .B(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_43), .A2(n_119), .B1(n_682), .B2(n_715), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g1049 ( .A1(n_44), .A2(n_365), .B1(n_779), .B2(n_785), .Y(n_1049) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_45), .A2(n_127), .B1(n_630), .B2(n_664), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_46), .A2(n_79), .B1(n_637), .B2(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_47), .A2(n_319), .B1(n_641), .B2(n_715), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_48), .A2(n_100), .B1(n_468), .B2(n_635), .Y(n_741) );
AOI222xp33_ASAP7_75t_L g975 ( .A1(n_49), .A2(n_81), .B1(n_135), .B2(n_857), .C1(n_976), .C2(n_977), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_51), .A2(n_142), .B1(n_836), .B2(n_986), .Y(n_1002) );
INVx1_ASAP7_75t_L g1013 ( .A(n_52), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_53), .B(n_857), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_54), .A2(n_110), .B1(n_515), .B2(n_517), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_55), .A2(n_285), .B1(n_836), .B2(n_838), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_56), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g1053 ( .A1(n_57), .A2(n_120), .B1(n_559), .B2(n_782), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_58), .A2(n_230), .B1(n_468), .B2(n_471), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g1099 ( .A1(n_59), .A2(n_175), .B1(n_344), .B2(n_405), .C1(n_803), .C2(n_1100), .Y(n_1099) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_60), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_61), .A2(n_96), .B1(n_719), .B2(n_759), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_62), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_63), .A2(n_184), .B1(n_597), .B2(n_992), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_64), .A2(n_87), .B1(n_632), .B2(n_657), .Y(n_761) );
INVx1_ASAP7_75t_L g687 ( .A(n_65), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_66), .B(n_657), .Y(n_875) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_67), .A2(n_380), .B1(n_607), .B2(n_608), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_68), .Y(n_974) );
AOI22xp33_ASAP7_75t_SL g828 ( .A1(n_69), .A2(n_164), .B1(n_600), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_70), .A2(n_227), .B1(n_517), .B2(n_635), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_71), .A2(n_302), .B1(n_635), .B2(n_834), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_72), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_73), .A2(n_292), .B1(n_987), .B2(n_1134), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_74), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_75), .A2(n_338), .B1(n_838), .B2(n_1090), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_77), .A2(n_373), .B1(n_664), .B2(n_992), .Y(n_1008) );
INVx1_ASAP7_75t_L g1112 ( .A(n_78), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_78), .A2(n_1112), .B1(n_1114), .B2(n_1136), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_80), .Y(n_780) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_82), .A2(n_258), .B1(n_464), .B2(n_682), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_83), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_84), .A2(n_206), .B1(n_523), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_86), .A2(n_281), .B1(n_446), .B2(n_630), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_88), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_89), .A2(n_198), .B1(n_571), .B2(n_573), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g1082 ( .A(n_90), .Y(n_1082) );
AO22x2_ASAP7_75t_L g417 ( .A1(n_91), .A2(n_261), .B1(n_408), .B2(n_409), .Y(n_417) );
INVx1_ASAP7_75t_L g1070 ( .A(n_91), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_92), .A2(n_108), .B1(n_751), .B2(n_753), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_93), .A2(n_147), .B1(n_596), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_94), .A2(n_237), .B1(n_569), .B2(n_682), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_97), .A2(n_286), .B1(n_470), .B2(n_471), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_98), .A2(n_128), .B1(n_437), .B2(n_632), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_99), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_101), .A2(n_273), .B1(n_420), .B2(n_443), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_102), .A2(n_186), .B1(n_591), .B2(n_824), .Y(n_990) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_104), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_105), .A2(n_538), .B1(n_574), .B2(n_575), .Y(n_537) );
INVx1_ASAP7_75t_L g574 ( .A(n_105), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_106), .A2(n_371), .B1(n_549), .B2(n_659), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g743 ( .A1(n_107), .A2(n_114), .B1(n_177), .B2(n_545), .C1(n_706), .C2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_109), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_111), .A2(n_265), .B1(n_515), .B2(n_517), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_112), .Y(n_891) );
XOR2x2_ASAP7_75t_L g842 ( .A(n_113), .B(n_843), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_115), .A2(n_279), .B1(n_715), .B2(n_716), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_116), .Y(n_671) );
INVx1_ASAP7_75t_L g1074 ( .A(n_117), .Y(n_1074) );
XOR2x2_ASAP7_75t_L g1021 ( .A(n_121), .B(n_1022), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_122), .B(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_123), .A2(n_277), .B1(n_613), .B2(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_124), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_125), .Y(n_906) );
AO22x1_ASAP7_75t_L g745 ( .A1(n_126), .A2(n_746), .B1(n_747), .B2(n_765), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_126), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_129), .B(n_853), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_130), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_132), .A2(n_348), .B1(n_470), .B2(n_524), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g1126 ( .A(n_133), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_134), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_137), .A2(n_140), .B1(n_715), .B2(n_716), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_138), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_141), .A2(n_284), .B1(n_530), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_143), .A2(n_162), .B1(n_523), .B2(n_525), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_144), .A2(n_346), .B1(n_718), .B2(n_866), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_145), .A2(n_226), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_146), .A2(n_160), .B1(n_530), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_148), .A2(n_358), .B1(n_838), .B2(n_862), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_149), .A2(n_1077), .B1(n_1101), .B2(n_1102), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_149), .Y(n_1101) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_151), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_152), .A2(n_197), .B1(n_420), .B2(n_803), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_153), .A2(n_203), .B1(n_659), .B2(n_664), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_154), .A2(n_306), .B1(n_560), .B2(n_753), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_155), .A2(n_342), .B1(n_561), .B2(n_862), .Y(n_1054) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_156), .A2(n_252), .B1(n_718), .B2(n_719), .Y(n_717) );
AND2x6_ASAP7_75t_L g387 ( .A(n_158), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_158), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_159), .A2(n_289), .B1(n_528), .B2(n_866), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_161), .A2(n_266), .B1(n_552), .B2(n_586), .Y(n_585) );
AOI222xp33_ASAP7_75t_L g1018 ( .A1(n_165), .A2(n_241), .B1(n_260), .B2(n_405), .C1(n_549), .C2(n_552), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g881 ( .A(n_167), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_168), .A2(n_315), .B1(n_986), .B2(n_987), .Y(n_985) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_169), .A2(n_340), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g1019 ( .A(n_170), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g902 ( .A(n_171), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_172), .A2(n_359), .B1(n_461), .B2(n_464), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_173), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_174), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_176), .A2(n_250), .B1(n_528), .B2(n_566), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_178), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_179), .Y(n_790) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_180), .A2(n_251), .B1(n_408), .B2(n_412), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_180), .B(n_1072), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_181), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_182), .A2(n_213), .B1(n_526), .B2(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_183), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_185), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_187), .A2(n_370), .B1(n_566), .B2(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g584 ( .A(n_188), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_190), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_191), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g763 ( .A1(n_193), .A2(n_329), .B1(n_339), .B2(n_420), .C1(n_545), .C2(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_194), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_195), .A2(n_254), .B1(n_452), .B2(n_753), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_196), .A2(n_343), .B1(n_530), .B2(n_1051), .Y(n_1050) );
XOR2x2_ASAP7_75t_L g730 ( .A(n_199), .B(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_200), .A2(n_278), .B1(n_437), .B2(n_825), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_201), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_202), .Y(n_1097) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_205), .Y(n_1118) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_207), .A2(n_208), .B1(n_559), .B2(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g1015 ( .A(n_209), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_210), .A2(n_305), .B1(n_431), .B2(n_675), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_211), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_212), .B(n_803), .Y(n_802) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_214), .A2(n_383), .B(n_392), .C(n_1075), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_215), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_217), .A2(n_267), .B1(n_461), .B2(n_524), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_218), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g912 ( .A(n_219), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_220), .A2(n_299), .B1(n_682), .B2(n_738), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_221), .A2(n_248), .B1(n_501), .B2(n_597), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g1120 ( .A(n_222), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_224), .A2(n_288), .B1(n_464), .B2(n_603), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_225), .A2(n_301), .B1(n_744), .B2(n_992), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_228), .A2(n_290), .B1(n_517), .B2(n_641), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_229), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_231), .A2(n_368), .B1(n_531), .B2(n_610), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g1084 ( .A(n_232), .Y(n_1084) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_233), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_234), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_235), .Y(n_807) );
INVx1_ASAP7_75t_L g1011 ( .A(n_236), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_238), .A2(n_333), .B1(n_549), .B2(n_659), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_239), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_240), .A2(n_264), .B1(n_461), .B2(n_531), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_242), .A2(n_381), .B1(n_632), .B2(n_824), .C(n_971), .Y(n_970) );
AOI222xp33_ASAP7_75t_L g998 ( .A1(n_243), .A2(n_350), .B1(n_362), .B2(n_405), .C1(n_420), .C2(n_764), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_244), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_245), .A2(n_379), .B1(n_824), .B2(n_825), .Y(n_823) );
INVx2_ASAP7_75t_L g391 ( .A(n_247), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_249), .A2(n_282), .B1(n_501), .B2(n_848), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g812 ( .A(n_253), .B(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_256), .A2(n_693), .B1(n_694), .B2(n_725), .Y(n_692) );
CKINVDCx14_ASAP7_75t_R g725 ( .A(n_256), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_257), .A2(n_364), .B1(n_515), .B2(n_569), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_259), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_268), .A2(n_297), .B1(n_613), .B2(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_269), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_271), .A2(n_919), .B1(n_942), .B2(n_943), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g942 ( .A(n_271), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_272), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_274), .A2(n_377), .B1(n_519), .B2(n_653), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_275), .A2(n_369), .B1(n_528), .B2(n_530), .Y(n_1130) );
XOR2x2_ASAP7_75t_L g578 ( .A(n_276), .B(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_280), .Y(n_972) );
OA22x2_ASAP7_75t_L g619 ( .A1(n_283), .A2(n_620), .B1(n_621), .B2(n_645), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_283), .Y(n_620) );
INVx1_ASAP7_75t_L g408 ( .A(n_287), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_287), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_293), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_294), .B(n_657), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_295), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_296), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_298), .B(n_431), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_304), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_307), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_308), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_309), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_310), .A2(n_330), .B1(n_478), .B2(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g1086 ( .A(n_311), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_312), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_313), .B(n_437), .Y(n_436) );
OA22x2_ASAP7_75t_L g1038 ( .A1(n_314), .A2(n_1039), .B1(n_1040), .B2(n_1055), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_314), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_316), .A2(n_376), .B1(n_432), .B2(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g390 ( .A(n_318), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_320), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_322), .B(n_931), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_323), .Y(n_497) );
INVx1_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_326), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_327), .A2(n_332), .B1(n_517), .B2(n_610), .Y(n_661) );
INVx1_ASAP7_75t_L g1017 ( .A(n_328), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_331), .Y(n_963) );
AO22x2_ASAP7_75t_L g949 ( .A1(n_335), .A2(n_950), .B1(n_978), .B2(n_979), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_335), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_336), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_337), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_341), .A2(n_360), .B1(n_528), .B2(n_831), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_345), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_347), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_351), .Y(n_911) );
INVx1_ASAP7_75t_L g1005 ( .A(n_352), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g1117 ( .A(n_353), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_354), .B(n_431), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_355), .A2(n_372), .B1(n_452), .B2(n_456), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_356), .B(n_591), .Y(n_1028) );
XOR2x2_ASAP7_75t_L g982 ( .A(n_357), .B(n_983), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_363), .B(n_1007), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_366), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_367), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_374), .A2(n_483), .B1(n_533), .B2(n_534), .Y(n_482) );
INVx1_ASAP7_75t_L g533 ( .A(n_374), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_375), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_378), .A2(n_773), .B1(n_810), .B2(n_811), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_378), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_384), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_388), .Y(n_1066) );
OAI21xp5_ASAP7_75t_L g1110 ( .A1(n_389), .A2(n_1065), .B(n_1111), .Y(n_1110) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_917), .B1(n_1060), .B2(n_1061), .C(n_1062), .Y(n_392) );
INVx1_ASAP7_75t_L g1060 ( .A(n_393), .Y(n_1060) );
XNOR2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_769), .Y(n_393) );
XOR2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_615), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_535), .B2(n_614), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_399), .B1(n_481), .B2(n_482), .Y(n_397) );
INVx3_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
XNOR2xp5_ASAP7_75t_L g577 ( .A(n_399), .B(n_578), .Y(n_577) );
XOR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_480), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_449), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_429), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_418), .B(n_419), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g1042 ( .A1(n_403), .A2(n_1043), .B(n_1044), .Y(n_1042) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx4_ASAP7_75t_L g496 ( .A(n_405), .Y(n_496) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_405), .Y(n_545) );
INVx2_ASAP7_75t_L g670 ( .A(n_405), .Y(n_670) );
INVx2_ASAP7_75t_SL g799 ( .A(n_405), .Y(n_799) );
AND2x6_ASAP7_75t_L g405 ( .A(n_406), .B(n_413), .Y(n_405) );
AND2x4_ASAP7_75t_L g446 ( .A(n_406), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g510 ( .A(n_406), .Y(n_510) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_407), .B(n_415), .Y(n_425) );
INVx2_ASAP7_75t_L g434 ( .A(n_407), .Y(n_434) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_410), .Y(n_412) );
INVx2_ASAP7_75t_L g424 ( .A(n_411), .Y(n_424) );
AND2x2_ASAP7_75t_L g433 ( .A(n_411), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g441 ( .A(n_411), .B(n_434), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
AND2x6_ASAP7_75t_L g470 ( .A(n_413), .B(n_440), .Y(n_470) );
AND2x4_ASAP7_75t_L g473 ( .A(n_413), .B(n_433), .Y(n_473) );
AND2x2_ASAP7_75t_L g477 ( .A(n_413), .B(n_455), .Y(n_477) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
AND2x2_ASAP7_75t_L g435 ( .A(n_414), .B(n_417), .Y(n_435) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g454 ( .A(n_415), .B(n_448), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_415), .B(n_417), .Y(n_459) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_417), .Y(n_423) );
INVx1_ASAP7_75t_L g448 ( .A(n_417), .Y(n_448) );
INVx1_ASAP7_75t_L g498 ( .A(n_420), .Y(n_498) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_421), .Y(n_549) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_421), .Y(n_588) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_421), .Y(n_857) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_421), .Y(n_1100) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g428 ( .A(n_423), .Y(n_428) );
AND2x2_ASAP7_75t_L g455 ( .A(n_424), .B(n_434), .Y(n_455) );
INVx1_ASAP7_75t_L g465 ( .A(n_424), .Y(n_465) );
AND2x4_ASAP7_75t_L g427 ( .A(n_425), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g443 ( .A(n_425), .B(n_444), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g506 ( .A(n_425), .B(n_465), .Y(n_506) );
INVx2_ASAP7_75t_L g707 ( .A(n_426), .Y(n_707) );
BUFx4f_ASAP7_75t_SL g764 ( .A(n_426), .Y(n_764) );
BUFx12f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_427), .Y(n_552) );
INVx1_ASAP7_75t_L g819 ( .A(n_427), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_436), .C(n_442), .Y(n_429) );
BUFx4f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g592 ( .A(n_432), .Y(n_592) );
BUFx2_ASAP7_75t_L g632 ( .A(n_432), .Y(n_632) );
BUFx2_ASAP7_75t_L g855 ( .A(n_432), .Y(n_855) );
AND2x6_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
AND2x2_ASAP7_75t_L g463 ( .A(n_433), .B(n_454), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_433), .B(n_435), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g958 ( .A(n_433), .B(n_454), .Y(n_958) );
AND2x4_ASAP7_75t_L g439 ( .A(n_435), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g479 ( .A(n_435), .B(n_455), .Y(n_479) );
INVx1_ASAP7_75t_L g489 ( .A(n_435), .Y(n_489) );
BUFx2_ASAP7_75t_L g1007 ( .A(n_437), .Y(n_1007) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g594 ( .A(n_438), .Y(n_594) );
INVx5_ASAP7_75t_L g657 ( .A(n_438), .Y(n_657) );
INVx2_ASAP7_75t_L g675 ( .A(n_438), .Y(n_675) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g488 ( .A(n_441), .B(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g596 ( .A(n_443), .Y(n_596) );
BUFx2_ASAP7_75t_L g630 ( .A(n_443), .Y(n_630) );
BUFx3_ASAP7_75t_L g659 ( .A(n_443), .Y(n_659) );
INVx1_ASAP7_75t_L g993 ( .A(n_443), .Y(n_993) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x6_ASAP7_75t_L g532 ( .A(n_445), .B(n_459), .Y(n_532) );
BUFx2_ASAP7_75t_SL g597 ( .A(n_446), .Y(n_597) );
BUFx3_ASAP7_75t_L g664 ( .A(n_446), .Y(n_664) );
BUFx2_ASAP7_75t_SL g744 ( .A(n_446), .Y(n_744) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_446), .Y(n_850) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_466), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
INVx1_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
BUFx2_ASAP7_75t_L g834 ( .A(n_452), .Y(n_834) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g560 ( .A(n_453), .Y(n_560) );
BUFx3_ASAP7_75t_L g610 ( .A(n_453), .Y(n_610) );
BUFx3_ASAP7_75t_L g723 ( .A(n_453), .Y(n_723) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_454), .B(n_455), .Y(n_789) );
AND2x4_ASAP7_75t_L g457 ( .A(n_455), .B(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
BUFx3_ASAP7_75t_L g562 ( .A(n_457), .Y(n_562) );
BUFx2_ASAP7_75t_SL g613 ( .A(n_457), .Y(n_613) );
INVx1_ASAP7_75t_L g739 ( .A(n_457), .Y(n_739) );
BUFx3_ASAP7_75t_L g753 ( .A(n_457), .Y(n_753) );
BUFx3_ASAP7_75t_L g838 ( .A(n_457), .Y(n_838) );
BUFx2_ASAP7_75t_SL g898 ( .A(n_457), .Y(n_898) );
AND2x2_ASAP7_75t_L g464 ( .A(n_458), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_461), .Y(n_1051) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g529 ( .A(n_462), .Y(n_529) );
INVx5_ASAP7_75t_L g572 ( .A(n_462), .Y(n_572) );
INVx1_ASAP7_75t_L g638 ( .A(n_462), .Y(n_638) );
INVx3_ASAP7_75t_L g759 ( .A(n_462), .Y(n_759) );
INVx8_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_474), .Y(n_466) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g519 ( .A(n_469), .Y(n_519) );
INVx3_ASAP7_75t_L g641 ( .A(n_469), .Y(n_641) );
INVx4_ASAP7_75t_L g782 ( .A(n_469), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_469), .A2(n_784), .B1(n_963), .B2(n_964), .Y(n_962) );
INVx11_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx11_ASAP7_75t_L g565 ( .A(n_470), .Y(n_565) );
INVx1_ASAP7_75t_L g892 ( .A(n_471), .Y(n_892) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
INVx2_ASAP7_75t_L g566 ( .A(n_472), .Y(n_566) );
INVx2_ASAP7_75t_L g612 ( .A(n_472), .Y(n_612) );
INVx6_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g635 ( .A(n_473), .Y(n_635) );
BUFx3_ASAP7_75t_L g653 ( .A(n_473), .Y(n_653) );
BUFx3_ASAP7_75t_L g785 ( .A(n_473), .Y(n_785) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g862 ( .A(n_476), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_476), .A2(n_778), .B1(n_953), .B2(n_954), .Y(n_952) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_477), .Y(n_524) );
BUFx2_ASAP7_75t_SL g715 ( .A(n_477), .Y(n_715) );
BUFx2_ASAP7_75t_SL g986 ( .A(n_477), .Y(n_986) );
INVx1_ASAP7_75t_L g644 ( .A(n_478), .Y(n_644) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g526 ( .A(n_479), .Y(n_526) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_479), .Y(n_603) );
INVx2_ASAP7_75t_L g683 ( .A(n_479), .Y(n_683) );
BUFx3_ASAP7_75t_L g716 ( .A(n_479), .Y(n_716) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g534 ( .A(n_483), .Y(n_534) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_484), .B(n_512), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .C(n_502), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_490), .B2(n_491), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_487), .A2(n_491), .B1(n_541), .B2(n_542), .Y(n_540) );
OAI221xp5_ASAP7_75t_SL g1095 ( .A1(n_487), .A2(n_925), .B1(n_1096), .B2(n_1097), .C(n_1098), .Y(n_1095) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g699 ( .A(n_488), .Y(n_699) );
BUFx3_ASAP7_75t_L g910 ( .A(n_488), .Y(n_910) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g797 ( .A(n_492), .Y(n_797) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx3_ASAP7_75t_L g702 ( .A(n_493), .Y(n_702) );
OAI221xp5_ASAP7_75t_SL g494 ( .A1(n_495), .A2(n_497), .B1(n_498), .B2(n_499), .C(n_500), .Y(n_494) );
OAI21xp5_ASAP7_75t_SL g703 ( .A1(n_495), .A2(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g976 ( .A(n_495), .Y(n_976) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_496), .A2(n_904), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_903) );
OAI222xp33_ASAP7_75t_L g623 ( .A1(n_498), .A2(n_582), .B1(n_624), .B2(n_625), .C1(n_626), .C2(n_627), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g798 ( .A1(n_498), .A2(n_799), .B1(n_800), .B2(n_801), .C(n_802), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g927 ( .A1(n_498), .A2(n_544), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_927) );
BUFx2_ASAP7_75t_L g803 ( .A(n_501), .Y(n_803) );
INVx2_ASAP7_75t_L g905 ( .A(n_501), .Y(n_905) );
BUFx3_ASAP7_75t_L g977 ( .A(n_501), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_507), .B2(n_508), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_504), .A2(n_509), .B1(n_901), .B2(n_902), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_504), .A2(n_808), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
INVx3_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g806 ( .A(n_505), .Y(n_806) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_506), .A2(n_508), .B1(n_554), .B2(n_555), .Y(n_553) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_506), .Y(n_710) );
BUFx3_ASAP7_75t_L g973 ( .A(n_506), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_508), .A2(n_972), .B1(n_973), .B2(n_974), .Y(n_971) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_509), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
CKINVDCx16_ASAP7_75t_R g809 ( .A(n_509), .Y(n_809) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g1135 ( .A(n_517), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g569 ( .A(n_524), .Y(n_569) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_524), .Y(n_607) );
INVx3_ASAP7_75t_L g776 ( .A(n_524), .Y(n_776) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g960 ( .A(n_530), .Y(n_960) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g573 ( .A(n_531), .Y(n_573) );
BUFx2_ASAP7_75t_L g719 ( .A(n_531), .Y(n_719) );
BUFx2_ASAP7_75t_L g866 ( .A(n_531), .Y(n_866) );
INVx6_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g792 ( .A(n_532), .Y(n_792) );
INVx1_ASAP7_75t_SL g831 ( .A(n_532), .Y(n_831) );
INVx1_ASAP7_75t_L g889 ( .A(n_532), .Y(n_889) );
INVx1_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B1(n_576), .B2(n_577), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g575 ( .A(n_538), .Y(n_575) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_556), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .C(n_553), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_546), .B1(n_547), .B2(n_550), .C(n_551), .Y(n_543) );
OAI222xp33_ASAP7_75t_L g815 ( .A1(n_544), .A2(n_816), .B1(n_817), .B2(n_818), .C1(n_819), .C2(n_820), .Y(n_815) );
OAI21xp5_ASAP7_75t_SL g1024 ( .A1(n_544), .A2(n_1025), .B(n_1026), .Y(n_1024) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g626 ( .A(n_552), .Y(n_626) );
BUFx4f_ASAP7_75t_L g931 ( .A(n_552), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_567), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .Y(n_557) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g969 ( .A(n_561), .Y(n_969) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_SL g602 ( .A(n_565), .Y(n_602) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_565), .Y(n_757) );
INVx1_ASAP7_75t_L g997 ( .A(n_565), .Y(n_997) );
INVx5_ASAP7_75t_SL g1092 ( .A(n_565), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_572), .Y(n_718) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND3x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_598), .C(n_605), .Y(n_579) );
NOR2x1_ASAP7_75t_SL g580 ( .A(n_581), .B(n_589), .Y(n_580) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_584), .B(n_585), .Y(n_581) );
OAI221xp5_ASAP7_75t_SL g1119 ( .A1(n_582), .A2(n_1120), .B1(n_1121), .B2(n_1122), .C(n_1123), .Y(n_1119) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g817 ( .A(n_588), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .C(n_595), .Y(n_589) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g825 ( .A(n_592), .Y(n_825) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx4_ASAP7_75t_L g837 ( .A(n_603), .Y(n_837) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_611), .Y(n_605) );
INVx1_ASAP7_75t_SL g1085 ( .A(n_607), .Y(n_1085) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g1081 ( .A(n_612), .Y(n_1081) );
XNOR2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_689), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_646), .B2(n_647), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g645 ( .A(n_621), .Y(n_645) );
NAND3x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_633), .C(n_639), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g1016 ( .A(n_641), .Y(n_1016) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AO22x2_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_666), .B2(n_688), .Y(n_647) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
XOR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_665), .Y(n_649) );
NAND4xp75_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .C(n_660), .D(n_663), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx3_ASAP7_75t_L g752 ( .A(n_653), .Y(n_752) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_656), .B(n_658), .Y(n_655) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_657), .Y(n_824) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_657), .Y(n_853) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx2_ASAP7_75t_L g688 ( .A(n_666), .Y(n_688) );
XOR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_687), .Y(n_666) );
NAND2x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_678), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_671), .B(n_672), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .C(n_677), .Y(n_673) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_684), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_726), .B2(n_727), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_712), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_703), .C(n_708), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_700), .B2(n_701), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_698), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g923 ( .A(n_699), .Y(n_923) );
OA211x2_ASAP7_75t_L g873 ( .A1(n_701), .A2(n_874), .B(n_875), .C(n_876), .Y(n_873) );
OA211x2_ASAP7_75t_L g1004 ( .A1(n_701), .A2(n_1005), .B(n_1006), .C(n_1008), .Y(n_1004) );
BUFx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g926 ( .A(n_702), .Y(n_926) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_710), .A2(n_808), .B1(n_933), .B2(n_934), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_720), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
BUFx2_ASAP7_75t_L g779 ( .A(n_716), .Y(n_779) );
INVxp67_ASAP7_75t_L g1087 ( .A(n_716), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .Y(n_720) );
BUFx4f_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_745), .B1(n_766), .B2(n_768), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_730), .Y(n_767) );
XOR2x2_ASAP7_75t_L g882 ( .A(n_730), .B(n_883), .Y(n_882) );
NAND4xp75_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .C(n_740), .D(n_743), .Y(n_731) );
AND2x2_ASAP7_75t_SL g732 ( .A(n_733), .B(n_734), .Y(n_732) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g768 ( .A(n_745), .Y(n_768) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
NAND4xp75_ASAP7_75t_SL g747 ( .A(n_748), .B(n_754), .C(n_760), .D(n_763), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVxp67_ASAP7_75t_L g1012 ( .A(n_753), .Y(n_1012) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_SL g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVxp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
XOR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_841), .Y(n_769) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_812), .B1(n_839), .B2(n_840), .Y(n_770) );
INVx2_ASAP7_75t_L g839 ( .A(n_771), .Y(n_839) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g811 ( .A(n_773), .Y(n_811) );
AND2x2_ASAP7_75t_SL g773 ( .A(n_774), .B(n_793), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_783), .Y(n_774) );
OAI221xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_780), .C(n_781), .Y(n_775) );
INVx2_ASAP7_75t_L g829 ( .A(n_776), .Y(n_829) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI221xp5_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_786), .B1(n_787), .B2(n_790), .C(n_791), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_787), .A2(n_891), .B1(n_892), .B2(n_893), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_787), .A2(n_1011), .B1(n_1012), .B2(n_1013), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_787), .A2(n_1080), .B1(n_1081), .B2(n_1082), .Y(n_1079) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g967 ( .A(n_788), .Y(n_967) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_798), .C(n_804), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_797), .A2(n_909), .B1(n_910), .B2(n_911), .Y(n_908) );
OAI21xp5_ASAP7_75t_SL g845 ( .A1(n_799), .A2(n_846), .B(n_847), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_804) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g840 ( .A(n_812), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_826), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_821), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_832), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
INVx3_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_837), .A2(n_895), .B1(n_896), .B2(n_897), .Y(n_894) );
INVx4_ASAP7_75t_L g987 ( .A(n_837), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_867), .B1(n_915), .B2(n_916), .Y(n_841) );
INVx2_ASAP7_75t_L g915 ( .A(n_842), .Y(n_915) );
NAND2xp5_ASAP7_75t_SL g843 ( .A(n_844), .B(n_858), .Y(n_843) );
NOR2xp33_ASAP7_75t_SL g844 ( .A(n_845), .B(n_851), .Y(n_844) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_SL g849 ( .A(n_850), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_854), .C(n_856), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g1121 ( .A(n_857), .Y(n_1121) );
NOR2x1_ASAP7_75t_L g858 ( .A(n_859), .B(n_863), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
INVx1_ASAP7_75t_L g916 ( .A(n_867), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_882), .B1(n_913), .B2(n_914), .Y(n_867) );
INVx3_ASAP7_75t_SL g914 ( .A(n_868), .Y(n_914) );
XOR2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_881), .Y(n_868) );
NAND4xp75_ASAP7_75t_L g869 ( .A(n_870), .B(n_873), .C(n_877), .D(n_880), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
INVx1_ASAP7_75t_L g913 ( .A(n_882), .Y(n_913) );
XOR2xp5_ASAP7_75t_SL g883 ( .A(n_884), .B(n_912), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_899), .Y(n_884) );
NOR3xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_890), .C(n_894), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_892), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
INVx1_ASAP7_75t_SL g897 ( .A(n_898), .Y(n_897) );
NOR3xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_903), .C(n_908), .Y(n_899) );
INVx1_ASAP7_75t_L g1061 ( .A(n_917), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_944), .B1(n_945), .B2(n_1059), .Y(n_917) );
INVx1_ASAP7_75t_L g1059 ( .A(n_918), .Y(n_1059) );
INVx2_ASAP7_75t_L g943 ( .A(n_919), .Y(n_943) );
AND2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_935), .Y(n_919) );
NOR3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_927), .C(n_932), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_923), .A2(n_925), .B1(n_1117), .B2(n_1118), .Y(n_1116) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_936), .B(n_939), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
INVx1_ASAP7_75t_SL g944 ( .A(n_945), .Y(n_944) );
OAI22xp5_ASAP7_75t_SL g945 ( .A1(n_946), .A2(n_1020), .B1(n_1057), .B2(n_1058), .Y(n_945) );
INVx1_ASAP7_75t_L g1057 ( .A(n_946), .Y(n_1057) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_948), .A2(n_949), .B1(n_980), .B2(n_981), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g979 ( .A(n_950), .Y(n_979) );
AND4x1_ASAP7_75t_L g950 ( .A(n_951), .B(n_961), .C(n_970), .D(n_975), .Y(n_950) );
NOR2xp33_ASAP7_75t_SL g951 ( .A(n_952), .B(n_955), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_957), .B1(n_959), .B2(n_960), .Y(n_955) );
BUFx2_ASAP7_75t_R g957 ( .A(n_958), .Y(n_957) );
NOR2xp33_ASAP7_75t_SL g961 ( .A(n_962), .B(n_965), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_965) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
XOR2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_999), .Y(n_981) );
NAND4xp75_ASAP7_75t_L g983 ( .A(n_984), .B(n_989), .C(n_994), .D(n_998), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_985), .B(n_988), .Y(n_984) );
AND2x2_ASAP7_75t_SL g989 ( .A(n_990), .B(n_991), .Y(n_989) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AND2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
XOR2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1019), .Y(n_999) );
NAND4xp75_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1004), .C(n_1009), .D(n_1018), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1014), .Y(n_1009) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1020), .Y(n_1058) );
OAI22xp5_ASAP7_75t_SL g1020 ( .A1(n_1021), .A2(n_1037), .B1(n_1038), .B2(n_1056), .Y(n_1020) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1021), .Y(n_1056) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1031), .C(n_1034), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1027), .Y(n_1023) );
NAND3xp33_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .C(n_1030), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_SL g1055 ( .A(n_1040), .Y(n_1055) );
NAND3x1_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1048), .C(n_1052), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1045), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1047), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
NOR2x1_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1068), .Y(n_1063) );
OR2x2_ASAP7_75t_SL g1139 ( .A(n_1064), .B(n_1069), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1067), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_1065), .Y(n_1105) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1066), .B(n_1108), .Y(n_1111) );
CKINVDCx16_ASAP7_75t_R g1108 ( .A(n_1067), .Y(n_1108) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_1069), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1071), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1074), .Y(n_1072) );
OAI322xp33_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1103), .A3(n_1106), .B1(n_1109), .B2(n_1112), .C1(n_1113), .C2(n_1137), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_1077), .Y(n_1102) );
AND4x1_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1088), .C(n_1094), .D(n_1099), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1083), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1093), .Y(n_1088) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
CKINVDCx16_ASAP7_75t_R g1109 ( .A(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1114), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1127), .Y(n_1114) );
NOR3xp33_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1119), .C(n_1124), .Y(n_1115) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1131), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1130), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1137 ( .A(n_1138), .Y(n_1137) );
CKINVDCx20_ASAP7_75t_R g1138 ( .A(n_1139), .Y(n_1138) );
endmodule