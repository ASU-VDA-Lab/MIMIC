module fake_jpeg_7722_n_286 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_18),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_38),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_33),
.B(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_53),
.B1(n_46),
.B2(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_35),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_61),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_41),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_15),
.B(n_24),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_11),
.Y(n_118)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_59),
.B1(n_57),
.B2(n_50),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_94),
.B1(n_99),
.B2(n_45),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_20),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_59),
.B1(n_31),
.B2(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_22),
.B1(n_18),
.B2(n_40),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_18),
.B1(n_56),
.B2(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_31),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_32),
.B1(n_31),
.B2(n_49),
.Y(n_99)
);

AOI22x1_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_14),
.B1(n_29),
.B2(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_44),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_116),
.Y(n_130)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_105),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_111),
.B1(n_120),
.B2(n_126),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_39),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_114),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_80),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_121),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_14),
.B1(n_29),
.B2(n_26),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_49),
.B1(n_45),
.B2(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_43),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_39),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_83),
.B(n_100),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_39),
.B1(n_15),
.B2(n_28),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_94),
.B1(n_97),
.B2(n_92),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_134),
.B1(n_140),
.B2(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_143),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_90),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_137),
.C(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_99),
.B1(n_91),
.B2(n_85),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_85),
.C(n_103),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_54),
.C(n_74),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_52),
.B1(n_51),
.B2(n_42),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_19),
.B1(n_28),
.B2(n_42),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_19),
.B1(n_16),
.B2(n_68),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_26),
.B1(n_105),
.B2(n_20),
.Y(n_173)
);

XOR2x1_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_122),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_124),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_69),
.C(n_89),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_1),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_144),
.C(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_156),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_153),
.B(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_123),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_160),
.B(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_167),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_113),
.B(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_113),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_170),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_23),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_132),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_138),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_174),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_127),
.B1(n_142),
.B2(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_154),
.B1(n_159),
.B2(n_157),
.Y(n_201)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_184),
.B1(n_196),
.B2(n_197),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_152),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_127),
.B1(n_141),
.B2(n_135),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_159),
.B1(n_172),
.B2(n_173),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_165),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_142),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_195),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_192),
.C(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_27),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_105),
.C(n_107),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_27),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_29),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_211),
.C(n_215),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_168),
.B1(n_167),
.B2(n_158),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_157),
.B(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_204),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_107),
.B1(n_98),
.B2(n_68),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_98),
.B1(n_23),
.B2(n_17),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_1),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_98),
.C(n_25),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_1),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_25),
.B1(n_8),
.B2(n_3),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_193),
.B1(n_189),
.B2(n_177),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_8),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_228),
.C(n_203),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_185),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_195),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_205),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_187),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_178),
.B1(n_180),
.B2(n_187),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_183),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_175),
.B1(n_183),
.B2(n_197),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_217),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

OAI322xp33_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_222),
.A3(n_226),
.B1(n_212),
.B2(n_218),
.C1(n_200),
.C2(n_194),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_9),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_190),
.C(n_175),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_244),
.C(n_7),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_225),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_191),
.C(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_230),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_259),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_258),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_7),
.C(n_3),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_3),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_264),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_239),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_268),
.B(n_5),
.Y(n_273)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_270),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_243),
.C(n_251),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_266),
.Y(n_278)
);

OAI211xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_249),
.B(n_4),
.C(n_5),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_274),
.B(n_272),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_281),
.A2(n_280),
.B(n_277),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_282),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_10),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_10),
.B(n_12),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_2),
.Y(n_286)
);


endmodule