module real_aes_17712_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1730;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1691;
wire n_640;
wire n_1721;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g799 ( .A(n_0), .Y(n_799) );
OAI211xp5_ASAP7_75t_L g973 ( .A1(n_1), .A2(n_550), .B(n_666), .C(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g986 ( .A(n_1), .Y(n_986) );
INVx1_ASAP7_75t_L g1704 ( .A(n_2), .Y(n_1704) );
OAI211xp5_ASAP7_75t_L g1733 ( .A1(n_2), .A2(n_1734), .B(n_1735), .C(n_1739), .Y(n_1733) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_3), .A2(n_81), .B1(n_1412), .B2(n_1415), .Y(n_1437) );
AND2x2_ASAP7_75t_L g329 ( .A(n_4), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g345 ( .A(n_4), .Y(n_345) );
AND2x2_ASAP7_75t_L g355 ( .A(n_4), .B(n_223), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_4), .B(n_344), .Y(n_579) );
OAI211xp5_ASAP7_75t_SL g818 ( .A1(n_5), .A2(n_538), .B(n_689), .C(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g831 ( .A(n_5), .Y(n_831) );
INVx1_ASAP7_75t_L g1323 ( .A(n_6), .Y(n_1323) );
INVx1_ASAP7_75t_L g840 ( .A(n_7), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_8), .A2(n_133), .B1(n_510), .B2(n_515), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_8), .A2(n_133), .B1(n_564), .B2(n_566), .Y(n_563) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_9), .A2(n_256), .B1(n_785), .B2(n_903), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g909 ( .A1(n_9), .A2(n_256), .B1(n_771), .B2(n_772), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_10), .A2(n_247), .B1(n_522), .B2(n_524), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_10), .A2(n_247), .B1(n_543), .B2(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g1082 ( .A(n_11), .Y(n_1082) );
OAI211xp5_ASAP7_75t_L g1321 ( .A1(n_12), .A2(n_552), .B(n_964), .C(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1333 ( .A(n_12), .Y(n_1333) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_13), .A2(n_41), .B1(n_1106), .B2(n_1108), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_13), .A2(n_41), .B1(n_524), .B2(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g993 ( .A(n_14), .Y(n_993) );
INVx1_ASAP7_75t_L g1634 ( .A(n_15), .Y(n_1634) );
OA222x2_ASAP7_75t_L g1653 ( .A1(n_15), .A2(n_135), .B1(n_169), .B2(n_1654), .C1(n_1656), .C2(n_1660), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1724 ( .A1(n_16), .A2(n_161), .B1(n_1725), .B2(n_1727), .Y(n_1724) );
INVx1_ASAP7_75t_L g1736 ( .A(n_16), .Y(n_1736) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_17), .A2(n_26), .B1(n_1065), .B2(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1170 ( .A(n_17), .Y(n_1170) );
INVx1_ASAP7_75t_L g869 ( .A(n_18), .Y(n_869) );
OAI211xp5_ASAP7_75t_L g880 ( .A1(n_18), .A2(n_666), .B(n_881), .C(n_882), .Y(n_880) );
INVx1_ASAP7_75t_L g843 ( .A(n_19), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_20), .Y(n_730) );
INVx2_ASAP7_75t_L g412 ( .A(n_21), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_22), .A2(n_311), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
INVx1_ASAP7_75t_L g1060 ( .A(n_22), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1625 ( .A1(n_23), .A2(n_173), .B1(n_1139), .B2(n_1620), .Y(n_1625) );
INVxp67_ASAP7_75t_SL g1674 ( .A(n_23), .Y(n_1674) );
INVx1_ASAP7_75t_L g417 ( .A(n_24), .Y(n_417) );
INVx1_ASAP7_75t_L g802 ( .A(n_25), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g1149 ( .A1(n_26), .A2(n_40), .B1(n_1049), .B2(n_1150), .C(n_1153), .Y(n_1149) );
INVx1_ASAP7_75t_L g928 ( .A(n_27), .Y(n_928) );
INVx1_ASAP7_75t_L g849 ( .A(n_28), .Y(n_849) );
HB1xp67_ASAP7_75t_L g1395 ( .A(n_29), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_29), .B(n_1393), .Y(n_1406) );
INVx1_ASAP7_75t_L g682 ( .A(n_30), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_31), .A2(n_291), .B1(n_324), .B2(n_1152), .Y(n_1349) );
INVxp67_ASAP7_75t_SL g1365 ( .A(n_31), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_32), .A2(n_185), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_32), .A2(n_237), .B1(n_1070), .B2(n_1072), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_33), .A2(n_192), .B1(n_455), .B2(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1155 ( .A(n_33), .Y(n_1155) );
INVx1_ASAP7_75t_L g1002 ( .A(n_34), .Y(n_1002) );
INVx1_ASAP7_75t_L g1083 ( .A(n_35), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_36), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_37), .A2(n_65), .B1(n_1405), .B2(n_1422), .Y(n_1436) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_38), .A2(n_166), .B1(n_776), .B2(n_874), .Y(n_895) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_38), .A2(n_166), .B1(n_522), .B2(n_825), .Y(n_910) );
INVx1_ASAP7_75t_L g1251 ( .A(n_39), .Y(n_1251) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_40), .A2(n_286), .B1(n_474), .B2(n_1135), .Y(n_1141) );
INVx1_ASAP7_75t_L g1296 ( .A(n_42), .Y(n_1296) );
AOI22xp33_ASAP7_75t_SL g1619 ( .A1(n_43), .A2(n_243), .B1(n_448), .B2(n_1620), .Y(n_1619) );
INVxp67_ASAP7_75t_SL g1668 ( .A(n_43), .Y(n_1668) );
INVx1_ASAP7_75t_L g1259 ( .A(n_44), .Y(n_1259) );
INVx1_ASAP7_75t_L g1716 ( .A(n_45), .Y(n_1716) );
AOI21xp33_ASAP7_75t_L g1740 ( .A1(n_45), .A2(n_338), .B(n_389), .Y(n_1740) );
AOI22xp33_ASAP7_75t_SL g1354 ( .A1(n_46), .A2(n_233), .B1(n_1152), .B2(n_1355), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_46), .A2(n_214), .B1(n_1367), .B2(n_1368), .Y(n_1366) );
OAI22xp33_ASAP7_75t_L g1325 ( .A1(n_47), .A2(n_124), .B1(n_878), .B2(n_1326), .Y(n_1325) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_47), .A2(n_124), .B1(n_652), .B2(n_772), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_48), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_49), .A2(n_62), .B1(n_467), .B2(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1154 ( .A(n_49), .Y(n_1154) );
OAI22xp33_ASAP7_75t_SL g1345 ( .A1(n_50), .A2(n_221), .B1(n_921), .B2(n_925), .Y(n_1345) );
INVx1_ASAP7_75t_L g1381 ( .A(n_50), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_51), .A2(n_90), .B1(n_347), .B2(n_352), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_51), .A2(n_203), .B1(n_455), .B2(n_459), .Y(n_454) );
INVx1_ASAP7_75t_L g1712 ( .A(n_52), .Y(n_1712) );
OAI22xp5_ASAP7_75t_L g1731 ( .A1(n_52), .A2(n_280), .B1(n_1216), .B2(n_1732), .Y(n_1731) );
INVx1_ASAP7_75t_L g690 ( .A(n_53), .Y(n_690) );
INVx1_ASAP7_75t_L g581 ( .A(n_54), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g1208 ( .A1(n_55), .A2(n_1026), .B(n_1209), .Y(n_1208) );
AOI221xp5_ASAP7_75t_L g1223 ( .A1(n_55), .A2(n_239), .B1(n_1137), .B2(n_1224), .C(n_1226), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_56), .Y(n_1128) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_57), .A2(n_97), .B1(n_1405), .B2(n_1422), .Y(n_1421) );
XOR2x2_ASAP7_75t_L g318 ( .A(n_58), .B(n_319), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g1442 ( .A1(n_58), .A2(n_228), .B1(n_1405), .B2(n_1422), .Y(n_1442) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_59), .A2(n_105), .B1(n_522), .B2(n_657), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_59), .A2(n_105), .B1(n_543), .B2(n_776), .Y(n_775) );
OAI222xp33_ASAP7_75t_L g1187 ( .A1(n_60), .A2(n_67), .B1(n_73), .B2(n_430), .C1(n_1188), .C2(n_1189), .Y(n_1187) );
AOI21xp33_ASAP7_75t_L g1044 ( .A1(n_61), .A2(n_1045), .B(n_1046), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_61), .A2(n_185), .B1(n_1062), .B2(n_1065), .Y(n_1061) );
INVx1_ASAP7_75t_L g1174 ( .A(n_62), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_63), .A2(n_68), .B1(n_1122), .B2(n_1245), .Y(n_1244) );
OAI22xp33_ASAP7_75t_L g1283 ( .A1(n_63), .A2(n_68), .B1(n_566), .B2(n_877), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_64), .Y(n_1194) );
CKINVDCx5p33_ASAP7_75t_R g1018 ( .A(n_66), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_69), .A2(n_275), .B1(n_378), .B2(n_383), .Y(n_1163) );
INVx1_ASAP7_75t_L g1176 ( .A(n_69), .Y(n_1176) );
INVx1_ASAP7_75t_L g1267 ( .A(n_70), .Y(n_1267) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_71), .B(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_71), .A2(n_218), .B1(n_1405), .B2(n_1422), .Y(n_1449) );
INVx1_ASAP7_75t_L g929 ( .A(n_72), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_73), .A2(n_309), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1430 ( .A1(n_74), .A2(n_222), .B1(n_1412), .B2(n_1415), .Y(n_1430) );
INVx1_ASAP7_75t_L g793 ( .A(n_75), .Y(n_793) );
INVx1_ASAP7_75t_L g820 ( .A(n_76), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g1431 ( .A1(n_77), .A2(n_87), .B1(n_1405), .B2(n_1432), .Y(n_1431) );
AO22x1_ASAP7_75t_L g1411 ( .A1(n_78), .A2(n_229), .B1(n_1412), .B2(n_1415), .Y(n_1411) );
INVx1_ASAP7_75t_L g649 ( .A(n_79), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_80), .A2(n_147), .B1(n_1029), .B2(n_1048), .Y(n_1210) );
INVx1_ASAP7_75t_L g1222 ( .A(n_80), .Y(n_1222) );
XNOR2xp5_ASAP7_75t_L g1291 ( .A(n_82), .B(n_1292), .Y(n_1291) );
OAI211xp5_ASAP7_75t_L g526 ( .A1(n_83), .A2(n_527), .B(n_531), .C(n_538), .Y(n_526) );
INVx1_ASAP7_75t_L g559 ( .A(n_83), .Y(n_559) );
INVx1_ASAP7_75t_L g1300 ( .A(n_84), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1626 ( .A1(n_85), .A2(n_100), .B1(n_1378), .B2(n_1627), .C(n_1628), .Y(n_1626) );
AOI22xp33_ASAP7_75t_SL g1675 ( .A1(n_85), .A2(n_243), .B1(n_1049), .B2(n_1152), .Y(n_1675) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_86), .A2(n_144), .B1(n_545), .B2(n_776), .Y(n_972) );
OAI22xp33_ASAP7_75t_L g980 ( .A1(n_86), .A2(n_144), .B1(n_522), .B2(n_825), .Y(n_980) );
INVx1_ASAP7_75t_L g1178 ( .A(n_87), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_88), .A2(n_134), .B1(n_524), .B2(n_1242), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_88), .A2(n_134), .B1(n_828), .B2(n_874), .Y(n_1279) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_89), .A2(n_95), .B1(n_656), .B2(n_657), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_89), .A2(n_95), .B1(n_671), .B2(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_90), .A2(n_111), .B1(n_464), .B2(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g950 ( .A(n_91), .Y(n_950) );
INVx1_ASAP7_75t_L g1723 ( .A(n_92), .Y(n_1723) );
AOI22xp33_ASAP7_75t_L g1738 ( .A1(n_92), .A2(n_227), .B1(n_324), .B2(n_1152), .Y(n_1738) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_93), .Y(n_1016) );
INVx1_ASAP7_75t_L g1393 ( .A(n_94), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_96), .A2(n_158), .B1(n_419), .B2(n_430), .Y(n_418) );
XOR2x2_ASAP7_75t_L g892 ( .A(n_97), .B(n_893), .Y(n_892) );
AO221x2_ASAP7_75t_L g1503 ( .A1(n_98), .A2(n_302), .B1(n_1412), .B2(n_1415), .C(n_1504), .Y(n_1503) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_99), .A2(n_538), .B(n_647), .C(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g669 ( .A(n_99), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g1665 ( .A1(n_100), .A2(n_152), .B1(n_333), .B2(n_1666), .C(n_1667), .Y(n_1665) );
INVx1_ASAP7_75t_L g537 ( .A(n_101), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g549 ( .A1(n_101), .A2(n_550), .B(n_552), .C(n_554), .Y(n_549) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_102), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_102), .A2(n_250), .B1(n_450), .B2(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_103), .A2(n_140), .B1(n_584), .B2(n_1084), .Y(n_1344) );
NOR2xp33_ASAP7_75t_L g1385 ( .A(n_103), .B(n_564), .Y(n_1385) );
INVx1_ASAP7_75t_L g808 ( .A(n_104), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_106), .Y(n_1146) );
INVx1_ASAP7_75t_L g804 ( .A(n_107), .Y(n_804) );
INVx1_ASAP7_75t_L g960 ( .A(n_108), .Y(n_960) );
INVx1_ASAP7_75t_L g806 ( .A(n_109), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_110), .A2(n_120), .B1(n_512), .B2(n_517), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_110), .A2(n_120), .B1(n_661), .B2(n_783), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_111), .A2(n_203), .B1(n_338), .B2(n_387), .C(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g698 ( .A(n_112), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_113), .A2(n_266), .B1(n_517), .B2(n_652), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_113), .A2(n_266), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g924 ( .A(n_114), .Y(n_924) );
INVx1_ASAP7_75t_L g868 ( .A(n_115), .Y(n_868) );
INVx1_ASAP7_75t_L g822 ( .A(n_116), .Y(n_822) );
OAI211xp5_ASAP7_75t_L g829 ( .A1(n_116), .A2(n_664), .B(n_666), .C(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g795 ( .A(n_117), .Y(n_795) );
INVx1_ASAP7_75t_L g834 ( .A(n_118), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g1718 ( .A1(n_119), .A2(n_252), .B1(n_1719), .B2(n_1720), .Y(n_1718) );
AOI21xp33_ASAP7_75t_L g1737 ( .A1(n_119), .A2(n_1046), .B(n_1666), .Y(n_1737) );
INVx1_ASAP7_75t_L g1112 ( .A(n_121), .Y(n_1112) );
OAI211xp5_ASAP7_75t_L g1118 ( .A1(n_121), .A2(n_595), .B(n_982), .C(n_1119), .Y(n_1118) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_122), .A2(n_250), .B1(n_333), .B2(n_336), .C(n_342), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_122), .A2(n_207), .B1(n_448), .B2(n_451), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_123), .A2(n_298), .B1(n_652), .B2(n_653), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_123), .A2(n_298), .B1(n_564), .B2(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g953 ( .A(n_125), .Y(n_953) );
INVx1_ASAP7_75t_L g955 ( .A(n_126), .Y(n_955) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_127), .A2(n_538), .B(n_761), .C(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g781 ( .A(n_127), .Y(n_781) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_128), .A2(n_168), .B1(n_656), .B2(n_657), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_128), .A2(n_168), .B1(n_545), .B2(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g1090 ( .A(n_129), .Y(n_1090) );
AO22x1_ASAP7_75t_L g1427 ( .A1(n_130), .A2(n_304), .B1(n_1412), .B2(n_1415), .Y(n_1427) );
OAI22xp33_ASAP7_75t_L g824 ( .A1(n_131), .A2(n_215), .B1(n_656), .B2(n_825), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_131), .A2(n_215), .B1(n_545), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g1262 ( .A(n_132), .Y(n_1262) );
INVx1_ASAP7_75t_L g1649 ( .A(n_135), .Y(n_1649) );
OAI221xp5_ASAP7_75t_L g1358 ( .A1(n_136), .A2(n_294), .B1(n_647), .B2(n_1359), .C(n_1360), .Y(n_1358) );
INVx1_ASAP7_75t_L g1377 ( .A(n_136), .Y(n_1377) );
INVx1_ASAP7_75t_L g1347 ( .A(n_137), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_137), .A2(n_233), .B1(n_1367), .B2(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1308 ( .A(n_138), .Y(n_1308) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_139), .Y(n_1351) );
INVx1_ASAP7_75t_L g1380 ( .A(n_140), .Y(n_1380) );
INVx1_ASAP7_75t_L g1303 ( .A(n_141), .Y(n_1303) );
INVx1_ASAP7_75t_L g901 ( .A(n_142), .Y(n_901) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_142), .A2(n_855), .B(n_906), .C(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g846 ( .A(n_143), .Y(n_846) );
INVx1_ASAP7_75t_L g534 ( .A(n_145), .Y(n_534) );
INVx1_ASAP7_75t_L g922 ( .A(n_146), .Y(n_922) );
INVxp67_ASAP7_75t_SL g1227 ( .A(n_147), .Y(n_1227) );
INVx1_ASAP7_75t_L g975 ( .A(n_148), .Y(n_975) );
INVx1_ASAP7_75t_L g1304 ( .A(n_149), .Y(n_1304) );
OAI22xp33_ASAP7_75t_L g1320 ( .A1(n_150), .A2(n_301), .B1(n_776), .B2(n_1106), .Y(n_1320) );
OAI22xp33_ASAP7_75t_L g1328 ( .A1(n_150), .A2(n_301), .B1(n_522), .B2(n_657), .Y(n_1328) );
OAI211xp5_ASAP7_75t_L g862 ( .A1(n_151), .A2(n_595), .B(n_863), .C(n_867), .Y(n_862) );
INVx1_ASAP7_75t_L g883 ( .A(n_151), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g1621 ( .A1(n_152), .A2(n_181), .B1(n_451), .B2(n_1622), .C(n_1624), .Y(n_1621) );
AO22x1_ASAP7_75t_L g1404 ( .A1(n_153), .A2(n_305), .B1(n_1405), .B2(n_1409), .Y(n_1404) );
CKINVDCx16_ASAP7_75t_R g1505 ( .A(n_154), .Y(n_1505) );
INVx1_ASAP7_75t_L g1298 ( .A(n_155), .Y(n_1298) );
INVx1_ASAP7_75t_L g926 ( .A(n_156), .Y(n_926) );
INVx1_ASAP7_75t_L g957 ( .A(n_157), .Y(n_957) );
OAI211xp5_ASAP7_75t_L g321 ( .A1(n_158), .A2(n_322), .B(n_331), .C(n_356), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g1022 ( .A1(n_159), .A2(n_299), .B1(n_1023), .B2(n_1025), .C(n_1026), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_159), .A2(n_311), .B1(n_624), .B2(n_1068), .Y(n_1067) );
XOR2x2_ASAP7_75t_L g1077 ( .A(n_160), .B(n_1078), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1741 ( .A1(n_161), .A2(n_252), .B1(n_324), .B2(n_1152), .Y(n_1741) );
INVx1_ASAP7_75t_L g1111 ( .A(n_162), .Y(n_1111) );
INVx1_ASAP7_75t_L g1093 ( .A(n_163), .Y(n_1093) );
INVx1_ASAP7_75t_L g1338 ( .A(n_164), .Y(n_1338) );
INVx1_ASAP7_75t_L g688 ( .A(n_165), .Y(n_688) );
INVx1_ASAP7_75t_L g650 ( .A(n_167), .Y(n_650) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_167), .A2(n_664), .B(n_666), .C(n_667), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g1643 ( .A1(n_169), .A2(n_170), .B1(n_726), .B2(n_1644), .C(n_1645), .Y(n_1643) );
INVxp67_ASAP7_75t_SL g1662 ( .A(n_170), .Y(n_1662) );
INVx1_ASAP7_75t_L g916 ( .A(n_171), .Y(n_916) );
INVx1_ASAP7_75t_L g1207 ( .A(n_172), .Y(n_1207) );
AOI221x1_ASAP7_75t_SL g1220 ( .A1(n_172), .A2(n_234), .B1(n_464), .B2(n_1137), .C(n_1221), .Y(n_1220) );
INVxp33_ASAP7_75t_SL g1669 ( .A(n_173), .Y(n_1669) );
INVx1_ASAP7_75t_L g839 ( .A(n_174), .Y(n_839) );
INVx1_ASAP7_75t_L g357 ( .A(n_175), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_175), .A2(n_278), .B1(n_488), .B2(n_494), .Y(n_487) );
AOI21xp33_ASAP7_75t_L g1213 ( .A1(n_176), .A2(n_1045), .B(n_1046), .Y(n_1213) );
INVx1_ASAP7_75t_L g1228 ( .A(n_176), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_177), .A2(n_232), .B1(n_365), .B2(n_369), .C(n_375), .Y(n_364) );
INVx1_ASAP7_75t_L g477 ( .A(n_177), .Y(n_477) );
INVx2_ASAP7_75t_L g1408 ( .A(n_178), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_178), .B(n_272), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_178), .B(n_1414), .Y(n_1416) );
OAI22xp33_ASAP7_75t_L g1113 ( .A1(n_179), .A2(n_230), .B1(n_661), .B2(n_903), .Y(n_1113) );
OAI22xp33_ASAP7_75t_L g1121 ( .A1(n_179), .A2(n_230), .B1(n_652), .B2(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1239 ( .A(n_180), .Y(n_1239) );
INVx1_ASAP7_75t_L g1672 ( .A(n_181), .Y(n_1672) );
INVx1_ASAP7_75t_L g900 ( .A(n_182), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_183), .A2(n_991), .B1(n_1073), .B2(n_1074), .Y(n_990) );
INVxp67_ASAP7_75t_L g1074 ( .A(n_183), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1235 ( .A1(n_184), .A2(n_1236), .B(n_1237), .C(n_1238), .Y(n_1235) );
INVx1_ASAP7_75t_L g1282 ( .A(n_184), .Y(n_1282) );
XOR2x2_ASAP7_75t_L g502 ( .A(n_186), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g976 ( .A(n_187), .Y(n_976) );
OAI211xp5_ASAP7_75t_L g981 ( .A1(n_187), .A2(n_683), .B(n_982), .C(n_983), .Y(n_981) );
XOR2x2_ASAP7_75t_L g711 ( .A(n_188), .B(n_712), .Y(n_711) );
OAI221xp5_ASAP7_75t_SL g1010 ( .A1(n_189), .A2(n_267), .B1(n_1011), .B2(n_1013), .C(n_1015), .Y(n_1010) );
INVx1_ASAP7_75t_L g1037 ( .A(n_189), .Y(n_1037) );
INVx1_ASAP7_75t_L g1648 ( .A(n_190), .Y(n_1648) );
OAI22xp5_ASAP7_75t_L g1680 ( .A1(n_190), .A2(n_211), .B1(n_420), .B2(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1087 ( .A(n_191), .Y(n_1087) );
INVx1_ASAP7_75t_L g1172 ( .A(n_192), .Y(n_1172) );
INVx1_ASAP7_75t_L g1088 ( .A(n_193), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_194), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g440 ( .A(n_194), .Y(n_440) );
INVx1_ASAP7_75t_L g472 ( .A(n_194), .Y(n_472) );
INVx1_ASAP7_75t_L g1301 ( .A(n_195), .Y(n_1301) );
INVx1_ASAP7_75t_L g851 ( .A(n_196), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_197), .A2(n_201), .B1(n_771), .B2(n_772), .Y(n_770) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_197), .A2(n_201), .B1(n_783), .B2(n_785), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_198), .Y(n_725) );
INVx1_ASAP7_75t_L g1185 ( .A(n_199), .Y(n_1185) );
INVx1_ASAP7_75t_L g844 ( .A(n_200), .Y(n_844) );
BUFx3_ASAP7_75t_L g405 ( .A(n_202), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_204), .A2(n_208), .B1(n_1412), .B2(n_1415), .Y(n_1450) );
INVx1_ASAP7_75t_L g996 ( .A(n_205), .Y(n_996) );
INVx1_ASAP7_75t_L g1097 ( .A(n_206), .Y(n_1097) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_207), .Y(n_381) );
OAI22xp5_ASAP7_75t_SL g1196 ( .A1(n_209), .A2(n_253), .B1(n_401), .B2(n_425), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_209), .Y(n_1205) );
INVx1_ASAP7_75t_L g678 ( .A(n_210), .Y(n_678) );
INVx1_ASAP7_75t_L g1632 ( .A(n_211), .Y(n_1632) );
INVx1_ASAP7_75t_L g914 ( .A(n_212), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_213), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g1348 ( .A1(n_214), .A2(n_1045), .B(n_1046), .Y(n_1348) );
INVx1_ASAP7_75t_L g585 ( .A(n_216), .Y(n_585) );
INVx1_ASAP7_75t_L g1257 ( .A(n_217), .Y(n_1257) );
INVx1_ASAP7_75t_L g918 ( .A(n_219), .Y(n_918) );
INVx1_ASAP7_75t_L g1708 ( .A(n_220), .Y(n_1708) );
INVx1_ASAP7_75t_L g1384 ( .A(n_221), .Y(n_1384) );
INVx1_ASAP7_75t_L g330 ( .A(n_223), .Y(n_330) );
BUFx3_ASAP7_75t_L g344 ( .A(n_223), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g1507 ( .A(n_224), .Y(n_1507) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_225), .A2(n_241), .B1(n_1412), .B2(n_1415), .Y(n_1441) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_226), .A2(n_277), .B1(n_878), .B2(n_903), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_226), .A2(n_277), .B1(n_652), .B2(n_653), .Y(n_987) );
INVx1_ASAP7_75t_L g1717 ( .A(n_227), .Y(n_1717) );
XNOR2xp5_ASAP7_75t_L g788 ( .A(n_231), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g482 ( .A(n_232), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_234), .A2(n_239), .B1(n_1029), .B2(n_1048), .Y(n_1214) );
INVx1_ASAP7_75t_L g800 ( .A(n_235), .Y(n_800) );
INVx1_ASAP7_75t_L g602 ( .A(n_236), .Y(n_602) );
INVx1_ASAP7_75t_L g1043 ( .A(n_237), .Y(n_1043) );
INVx1_ASAP7_75t_L g1240 ( .A(n_238), .Y(n_1240) );
OAI211xp5_ASAP7_75t_L g1280 ( .A1(n_238), .A2(n_552), .B(n_619), .C(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g680 ( .A(n_240), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_242), .Y(n_732) );
INVx1_ASAP7_75t_L g1263 ( .A(n_244), .Y(n_1263) );
INVx1_ASAP7_75t_L g598 ( .A(n_245), .Y(n_598) );
INVx1_ASAP7_75t_L g958 ( .A(n_246), .Y(n_958) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_248), .Y(n_1147) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_249), .A2(n_308), .B1(n_1412), .B2(n_1415), .Y(n_1420) );
AO22x1_ASAP7_75t_L g1426 ( .A1(n_251), .A2(n_258), .B1(n_1405), .B2(n_1422), .Y(n_1426) );
INVx1_ASAP7_75t_L g1200 ( .A(n_253), .Y(n_1200) );
INVx1_ASAP7_75t_L g594 ( .A(n_254), .Y(n_594) );
INVx1_ASAP7_75t_L g406 ( .A(n_255), .Y(n_406) );
INVx1_ASAP7_75t_L g436 ( .A(n_255), .Y(n_436) );
INVx1_ASAP7_75t_L g1324 ( .A(n_257), .Y(n_1324) );
OAI211xp5_ASAP7_75t_L g1329 ( .A1(n_257), .A2(n_906), .B(n_1330), .C(n_1332), .Y(n_1329) );
INVx1_ASAP7_75t_L g610 ( .A(n_259), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_260), .Y(n_766) );
INVxp67_ASAP7_75t_SL g1705 ( .A(n_261), .Y(n_1705) );
OAI221xp5_ASAP7_75t_L g1743 ( .A1(n_261), .A2(n_300), .B1(n_370), .B2(n_416), .C(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1646 ( .A(n_262), .Y(n_1646) );
NOR2xp33_ASAP7_75t_L g1651 ( .A(n_262), .B(n_998), .Y(n_1651) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_263), .Y(n_723) );
INVx1_ASAP7_75t_L g961 ( .A(n_264), .Y(n_961) );
INVx1_ASAP7_75t_L g1212 ( .A(n_265), .Y(n_1212) );
INVx1_ASAP7_75t_L g1052 ( .A(n_267), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1709 ( .A(n_268), .Y(n_1709) );
INVx1_ASAP7_75t_L g1091 ( .A(n_269), .Y(n_1091) );
AOI22xp5_ASAP7_75t_L g1231 ( .A1(n_270), .A2(n_1232), .B1(n_1233), .B2(n_1285), .Y(n_1231) );
INVxp67_ASAP7_75t_SL g1285 ( .A(n_270), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_271), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_272), .B(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1414 ( .A(n_272), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_273), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_274), .A2(n_1696), .B1(n_1697), .B2(n_1746), .Y(n_1695) );
CKINVDCx5p33_ASAP7_75t_R g1746 ( .A(n_274), .Y(n_1746) );
INVx1_ASAP7_75t_L g1131 ( .A(n_275), .Y(n_1131) );
OAI211xp5_ASAP7_75t_L g1109 ( .A1(n_276), .A2(n_666), .B(n_703), .C(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1120 ( .A(n_276), .Y(n_1120) );
INVx1_ASAP7_75t_L g360 ( .A(n_278), .Y(n_360) );
INVx1_ASAP7_75t_L g676 ( .A(n_279), .Y(n_676) );
INVx1_ASAP7_75t_L g1713 ( .A(n_280), .Y(n_1713) );
INVx1_ASAP7_75t_L g1357 ( .A(n_281), .Y(n_1357) );
INVx1_ASAP7_75t_L g769 ( .A(n_282), .Y(n_769) );
OAI211xp5_ASAP7_75t_L g777 ( .A1(n_282), .A2(n_666), .B(n_778), .C(n_780), .Y(n_777) );
INVx1_ASAP7_75t_L g1306 ( .A(n_283), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g1722 ( .A(n_284), .Y(n_1722) );
INVx1_ASAP7_75t_L g609 ( .A(n_285), .Y(n_609) );
AOI211xp5_ASAP7_75t_SL g1167 ( .A1(n_286), .A2(n_1168), .B(n_1169), .C(n_1171), .Y(n_1167) );
INVx1_ASAP7_75t_L g847 ( .A(n_287), .Y(n_847) );
AOI21xp5_ASAP7_75t_SL g1352 ( .A1(n_288), .A2(n_1045), .B(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1364 ( .A(n_288), .Y(n_1364) );
INVx1_ASAP7_75t_L g947 ( .A(n_289), .Y(n_947) );
XOR2x2_ASAP7_75t_L g942 ( .A(n_290), .B(n_943), .Y(n_942) );
INVxp67_ASAP7_75t_L g1370 ( .A(n_291), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g896 ( .A1(n_292), .A2(n_666), .B(n_897), .C(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g908 ( .A(n_292), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_293), .Y(n_717) );
INVxp67_ASAP7_75t_SL g1383 ( .A(n_294), .Y(n_1383) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
INVx1_ASAP7_75t_L g1253 ( .A(n_296), .Y(n_1253) );
INVx1_ASAP7_75t_L g1268 ( .A(n_297), .Y(n_1268) );
INVx1_ASAP7_75t_L g1059 ( .A(n_299), .Y(n_1059) );
INVx1_ASAP7_75t_L g1707 ( .A(n_300), .Y(n_1707) );
INVx1_ASAP7_75t_L g695 ( .A(n_303), .Y(n_695) );
INVx1_ASAP7_75t_L g1684 ( .A(n_304), .Y(n_1684) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_304), .A2(n_1691), .B1(n_1694), .B2(n_1747), .Y(n_1690) );
INVx1_ASAP7_75t_L g596 ( .A(n_306), .Y(n_596) );
INVx2_ASAP7_75t_L g397 ( .A(n_307), .Y(n_397) );
INVx1_ASAP7_75t_L g410 ( .A(n_307), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_307), .Y(n_415) );
INVx1_ASAP7_75t_L g1195 ( .A(n_309), .Y(n_1195) );
CKINVDCx5p33_ASAP7_75t_R g1132 ( .A(n_310), .Y(n_1132) );
AOI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_1388), .B(n_1399), .Y(n_312) );
XNOR2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_887), .Y(n_313) );
OA22x2_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_640), .B1(n_641), .B2(n_886), .Y(n_314) );
INVx1_ASAP7_75t_L g886 ( .A(n_315), .Y(n_886) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
XNOR2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_502), .Y(n_317) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_398), .C(n_442), .Y(n_319) );
OAI21xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_364), .B(n_392), .Y(n_320) );
INVx2_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_329), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_325), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_325), .Y(n_1049) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g335 ( .A(n_326), .B(n_328), .Y(n_335) );
INVx2_ASAP7_75t_L g341 ( .A(n_326), .Y(n_341) );
INVx1_ASAP7_75t_L g351 ( .A(n_326), .Y(n_351) );
BUFx2_ASAP7_75t_L g373 ( .A(n_326), .Y(n_373) );
OR2x2_ASAP7_75t_L g380 ( .A(n_326), .B(n_328), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_326), .B(n_327), .Y(n_384) );
NAND2x1_ASAP7_75t_L g530 ( .A(n_326), .B(n_328), .Y(n_530) );
OR2x2_ASAP7_75t_L g593 ( .A(n_326), .B(n_350), .Y(n_593) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g340 ( .A(n_328), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g350 ( .A(n_328), .Y(n_350) );
INVx1_ASAP7_75t_L g423 ( .A(n_328), .Y(n_423) );
AND2x2_ASAP7_75t_L g359 ( .A(n_329), .B(n_349), .Y(n_359) );
AND2x4_ASAP7_75t_L g362 ( .A(n_329), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_329), .B(n_334), .Y(n_368) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_329), .B(n_363), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_329), .B(n_352), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1159 ( .A(n_329), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1659 ( .A(n_329), .B(n_415), .Y(n_1659) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_330), .Y(n_514) );
AOI21xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_346), .B(n_354), .Y(n_331) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x6_ASAP7_75t_L g354 ( .A(n_334), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
AND2x2_ASAP7_75t_L g539 ( .A(n_334), .B(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g1025 ( .A(n_334), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_334), .Y(n_1168) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g866 ( .A(n_335), .Y(n_866) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g1666 ( .A(n_339), .Y(n_1666) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
AND2x4_ASAP7_75t_L g525 ( .A(n_340), .B(n_514), .Y(n_525) );
BUFx3_ASAP7_75t_L g1209 ( .A(n_340), .Y(n_1209) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_343), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_343), .B(n_408), .Y(n_692) );
AND2x4_ASAP7_75t_L g755 ( .A(n_343), .B(n_606), .Y(n_755) );
INVx4_ASAP7_75t_L g1046 ( .A(n_343), .Y(n_1046) );
OAI21xp33_ASAP7_75t_L g1169 ( .A1(n_343), .A2(n_921), .B(n_1170), .Y(n_1169) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
BUFx2_ASAP7_75t_L g520 ( .A(n_344), .Y(n_520) );
AND2x4_ASAP7_75t_L g536 ( .A(n_344), .B(n_422), .Y(n_536) );
AND2x4_ASAP7_75t_L g390 ( .A(n_345), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g506 ( .A(n_345), .Y(n_506) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g1028 ( .A(n_348), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_348), .Y(n_1032) );
INVx1_ASAP7_75t_L g1048 ( .A(n_348), .Y(n_1048) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_349), .B(n_355), .Y(n_416) );
BUFx6f_ASAP7_75t_L g1152 ( .A(n_349), .Y(n_1152) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_350), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1657 ( .A(n_352), .B(n_1658), .Y(n_1657) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g1355 ( .A(n_353), .Y(n_1355) );
AOI211xp5_ASAP7_75t_SL g1742 ( .A1(n_354), .A2(n_1053), .B(n_1708), .C(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_355), .B(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_355), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_355), .B(n_397), .Y(n_1679) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_360), .B2(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g1732 ( .A(n_358), .Y(n_1732) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g999 ( .A(n_359), .B(n_1000), .Y(n_999) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g1734 ( .A(n_362), .Y(n_1734) );
INVx1_ASAP7_75t_L g1024 ( .A(n_363), .Y(n_1024) );
BUFx6f_ASAP7_75t_L g1045 ( .A(n_363), .Y(n_1045) );
INVx2_ASAP7_75t_L g1162 ( .A(n_363), .Y(n_1162) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g1217 ( .A(n_366), .Y(n_1217) );
INVx4_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_368), .Y(n_1053) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g1036 ( .A(n_372), .Y(n_1036) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g533 ( .A(n_373), .B(n_520), .Y(n_533) );
AND2x2_ASAP7_75t_L g765 ( .A(n_373), .B(n_520), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_373), .A2(n_1034), .B1(n_1128), .B2(n_1146), .Y(n_1166) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_373), .Y(n_1204) );
INVx1_ASAP7_75t_L g1683 ( .A(n_373), .Y(n_1683) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_381), .B1(n_382), .B2(n_385), .C(n_386), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_376), .A2(n_696), .B1(n_717), .B2(n_738), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_376), .A2(n_725), .B1(n_732), .B2(n_757), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g813 ( .A1(n_376), .A2(n_588), .B1(n_793), .B2(n_806), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_376), .A2(n_696), .B1(n_960), .B2(n_961), .Y(n_959) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g584 ( .A(n_378), .Y(n_584) );
OR2x6_ASAP7_75t_L g656 ( .A(n_378), .B(n_523), .Y(n_656) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_378), .Y(n_677) );
BUFx3_ASAP7_75t_L g915 ( .A(n_378), .Y(n_915) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g513 ( .A(n_379), .Y(n_513) );
BUFx4f_ASAP7_75t_L g1096 ( .A(n_379), .Y(n_1096) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_382), .A2(n_694), .B1(n_800), .B2(n_804), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_382), .A2(n_694), .B1(n_844), .B2(n_847), .Y(n_858) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g519 ( .A(n_383), .B(n_520), .Y(n_519) );
INVx8_ASAP7_75t_L g589 ( .A(n_383), .Y(n_589) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g1026 ( .A(n_390), .Y(n_1026) );
OAI221xp5_ASAP7_75t_L g1153 ( .A1(n_390), .A2(n_753), .B1(n_1154), .B2(n_1155), .C(n_1156), .Y(n_1153) );
INVx1_ASAP7_75t_L g1353 ( .A(n_390), .Y(n_1353) );
INVxp67_ASAP7_75t_L g523 ( .A(n_391), .Y(n_523) );
INVx1_ASAP7_75t_L g540 ( .A(n_391), .Y(n_540) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g1729 ( .A1(n_393), .A2(n_1730), .B(n_1742), .Y(n_1729) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_394), .Y(n_1218) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI31xp33_ASAP7_75t_L g1148 ( .A1(n_395), .A2(n_1149), .A3(n_1157), .B(n_1167), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_395), .Y(n_1341) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND3x4_ASAP7_75t_L g445 ( .A(n_396), .B(n_440), .C(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g470 ( .A(n_397), .Y(n_470) );
AOI21xp33_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_417), .B(n_418), .Y(n_398) );
INVx8_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_413), .Y(n_400) );
INVx1_ASAP7_75t_L g1017 ( .A(n_401), .Y(n_1017) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_407), .Y(n_401) );
BUFx3_ASAP7_75t_L g803 ( .A(n_402), .Y(n_803) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_403), .Y(n_627) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g568 ( .A(n_404), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_405), .Y(n_433) );
AND2x4_ASAP7_75t_L g452 ( .A(n_405), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g491 ( .A(n_405), .B(n_435), .Y(n_491) );
INVx1_ASAP7_75t_L g428 ( .A(n_406), .Y(n_428) );
INVx2_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
OR2x2_ASAP7_75t_L g425 ( .A(n_407), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g493 ( .A(n_407), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_407), .Y(n_496) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_408), .Y(n_574) );
INVx1_ASAP7_75t_L g607 ( .A(n_408), .Y(n_607) );
OR2x2_ASAP7_75t_L g613 ( .A(n_408), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g424 ( .A(n_409), .Y(n_424) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g1642 ( .A(n_411), .Y(n_1642) );
INVx3_ASAP7_75t_L g438 ( .A(n_412), .Y(n_438) );
BUFx3_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
NAND2xp33_ASAP7_75t_SL g614 ( .A(n_412), .B(n_440), .Y(n_614) );
INVx1_ASAP7_75t_L g1655 ( .A(n_413), .Y(n_1655) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
AND2x4_ASAP7_75t_L g481 ( .A(n_414), .B(n_437), .Y(n_481) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g639 ( .A(n_415), .Y(n_639) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_425), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g1745 ( .A(n_421), .Y(n_1745) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g441 ( .A(n_424), .Y(n_441) );
INVx1_ASAP7_75t_L g507 ( .A(n_424), .Y(n_507) );
INVx1_ASAP7_75t_L g1000 ( .A(n_424), .Y(n_1000) );
INVx2_ASAP7_75t_L g1019 ( .A(n_425), .Y(n_1019) );
INVx4_ASAP7_75t_L g551 ( .A(n_426), .Y(n_551) );
INVx3_ASAP7_75t_L g704 ( .A(n_426), .Y(n_704) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_426), .Y(n_807) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g621 ( .A(n_427), .Y(n_621) );
BUFx2_ASAP7_75t_L g741 ( .A(n_427), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
BUFx2_ASAP7_75t_L g562 ( .A(n_428), .Y(n_562) );
AND2x4_ASAP7_75t_L g461 ( .A(n_429), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
BUFx2_ASAP7_75t_L g558 ( .A(n_429), .Y(n_558) );
INVx3_ASAP7_75t_L g994 ( .A(n_430), .Y(n_994) );
INVx5_ASAP7_75t_L g1177 ( .A(n_430), .Y(n_1177) );
OR2x6_ASAP7_75t_L g430 ( .A(n_431), .B(n_441), .Y(n_430) );
INVx2_ASAP7_75t_L g1650 ( .A(n_431), .Y(n_1650) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_432), .B(n_437), .Y(n_431) );
BUFx3_ASAP7_75t_L g450 ( .A(n_432), .Y(n_450) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_432), .Y(n_1064) );
INVx8_ASAP7_75t_L g1071 ( .A(n_432), .Y(n_1071) );
AND2x4_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AND2x4_ASAP7_75t_L g457 ( .A(n_433), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g458 ( .A(n_436), .Y(n_458) );
AND2x6_ASAP7_75t_L g1631 ( .A(n_437), .B(n_479), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_437), .B(n_486), .Y(n_1633) );
INVx1_ASAP7_75t_L g1637 ( .A(n_437), .Y(n_1637) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_438), .B(n_472), .Y(n_471) );
OR2x4_ASAP7_75t_L g545 ( .A(n_438), .B(n_491), .Y(n_545) );
INVx1_ASAP7_75t_L g548 ( .A(n_438), .Y(n_548) );
AND2x4_ASAP7_75t_L g553 ( .A(n_438), .B(n_452), .Y(n_553) );
OR2x6_ASAP7_75t_L g567 ( .A(n_438), .B(n_568), .Y(n_567) );
NAND3x1_ASAP7_75t_L g638 ( .A(n_438), .B(n_472), .C(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_440), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_487), .C(n_498), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_444), .B(n_476), .Y(n_443) );
AOI33xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .A3(n_454), .B1(n_463), .B2(n_468), .B3(n_473), .Y(n_444) );
AOI33xp33_ASAP7_75t_L g1133 ( .A1(n_445), .A2(n_468), .A3(n_1134), .B1(n_1136), .B2(n_1138), .B3(n_1141), .Y(n_1133) );
BUFx3_ASAP7_75t_L g1229 ( .A(n_445), .Y(n_1229) );
INVx3_ASAP7_75t_L g557 ( .A(n_446), .Y(n_557) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g1719 ( .A(n_450), .Y(n_1719) );
INVx1_ASAP7_75t_L g1726 ( .A(n_450), .Y(n_1726) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
BUFx2_ASAP7_75t_L g501 ( .A(n_452), .Y(n_501) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_452), .Y(n_1065) );
BUFx2_ASAP7_75t_L g1372 ( .A(n_452), .Y(n_1372) );
BUFx3_ASAP7_75t_L g1378 ( .A(n_452), .Y(n_1378) );
BUFx2_ASAP7_75t_L g1710 ( .A(n_452), .Y(n_1710) );
INVx1_ASAP7_75t_L g462 ( .A(n_453), .Y(n_462) );
INVx1_ASAP7_75t_L g969 ( .A(n_455), .Y(n_969) );
INVx1_ASAP7_75t_L g1101 ( .A(n_455), .Y(n_1101) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g547 ( .A(n_456), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g724 ( .A(n_456), .Y(n_724) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_456), .Y(n_935) );
INVx2_ASAP7_75t_L g1058 ( .A(n_456), .Y(n_1058) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_457), .Y(n_466) );
BUFx8_ASAP7_75t_L g497 ( .A(n_457), .Y(n_497) );
INVx2_ASAP7_75t_L g625 ( .A(n_457), .Y(n_625) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx5_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
BUFx12f_ASAP7_75t_L g1068 ( .A(n_461), .Y(n_1068) );
BUFx3_ASAP7_75t_L g1137 ( .A(n_461), .Y(n_1137) );
BUFx2_ASAP7_75t_L g1620 ( .A(n_461), .Y(n_1620) );
INVx1_ASAP7_75t_L g486 ( .A(n_462), .Y(n_486) );
INVx2_ASAP7_75t_L g1258 ( .A(n_464), .Y(n_1258) );
INVx1_ASAP7_75t_L g1297 ( .A(n_464), .Y(n_1297) );
INVx8_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g731 ( .A(n_465), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_465), .A2(n_726), .B1(n_922), .B2(n_929), .Y(n_936) );
INVx5_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_466), .Y(n_630) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_466), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_466), .A2(n_1135), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
INVx2_ASAP7_75t_SL g1623 ( .A(n_466), .Y(n_1623) );
INVx3_ASAP7_75t_L g1644 ( .A(n_466), .Y(n_1644) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI33xp33_ASAP7_75t_L g699 ( .A1(n_469), .A2(n_700), .A3(n_701), .B1(n_705), .B2(n_708), .B3(n_710), .Y(n_699) );
OAI33xp33_ASAP7_75t_L g791 ( .A1(n_469), .A2(n_700), .A3(n_792), .B1(n_798), .B2(n_801), .B3(n_805), .Y(n_791) );
OAI33xp33_ASAP7_75t_L g837 ( .A1(n_469), .A2(n_700), .A3(n_838), .B1(n_842), .B2(n_845), .B3(n_848), .Y(n_837) );
OAI33xp33_ASAP7_75t_L g1098 ( .A1(n_469), .A2(n_715), .A3(n_1099), .B1(n_1100), .B2(n_1102), .B3(n_1103), .Y(n_1098) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x4_ASAP7_75t_L g578 ( .A(n_470), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g1055 ( .A(n_470), .Y(n_1055) );
INVx3_ASAP7_75t_L g1629 ( .A(n_471), .Y(n_1629) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g1072 ( .A(n_475), .Y(n_1072) );
INVx2_ASAP7_75t_L g1368 ( .A(n_475), .Y(n_1368) );
INVx1_ASAP7_75t_L g1720 ( .A(n_475), .Y(n_1720) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_482), .B2(n_483), .Y(n_476) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
AND2x4_ASAP7_75t_SL g1012 ( .A(n_479), .B(n_481), .Y(n_1012) );
NAND2x1_ASAP7_75t_L g1193 ( .A(n_479), .B(n_481), .Y(n_1193) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g483 ( .A(n_481), .B(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g500 ( .A(n_481), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_SL g1014 ( .A(n_481), .B(n_484), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_483), .A2(n_1192), .B1(n_1194), .B2(n_1195), .C(n_1196), .Y(n_1191) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
INVx2_ASAP7_75t_SL g634 ( .A(n_489), .Y(n_634) );
OR2x6_ASAP7_75t_L g1001 ( .A(n_489), .B(n_492), .Y(n_1001) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g702 ( .A(n_490), .Y(n_702) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x4_ASAP7_75t_L g565 ( .A(n_491), .B(n_548), .Y(n_565) );
BUFx4f_ASAP7_75t_L g618 ( .A(n_491), .Y(n_618) );
BUFx3_ASAP7_75t_L g720 ( .A(n_491), .Y(n_720) );
BUFx3_ASAP7_75t_L g850 ( .A(n_491), .Y(n_850) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_493), .B(n_967), .Y(n_1005) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_495), .B(n_1143), .Y(n_1142) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_496), .B(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_SL g709 ( .A(n_497), .Y(n_709) );
INVx2_ASAP7_75t_SL g1225 ( .A(n_497), .Y(n_1225) );
INVx3_ASAP7_75t_L g1261 ( .A(n_497), .Y(n_1261) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
OAI211xp5_ASAP7_75t_SL g1056 ( .A1(n_499), .A2(n_612), .B(n_1057), .C(n_1066), .Y(n_1056) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_500), .A2(n_1012), .B1(n_1014), .B2(n_1146), .C(n_1147), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_500), .A2(n_637), .B1(n_1220), .B2(n_1223), .C(n_1229), .Y(n_1219) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_508), .B1(n_541), .B2(n_569), .C(n_575), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_SL g658 ( .A(n_505), .Y(n_658) );
BUFx3_ASAP7_75t_L g773 ( .A(n_505), .Y(n_773) );
OAI31xp33_ASAP7_75t_L g817 ( .A1(n_505), .A2(n_818), .A3(n_823), .B(n_824), .Y(n_817) );
BUFx2_ASAP7_75t_L g871 ( .A(n_505), .Y(n_871) );
OAI31xp33_ASAP7_75t_L g1234 ( .A1(n_505), .A2(n_1235), .A3(n_1241), .B(n_1244), .Y(n_1234) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g1398 ( .A(n_506), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1689 ( .A(n_506), .B(n_1390), .Y(n_1689) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .C(n_526), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_512), .Y(n_652) );
BUFx2_ASAP7_75t_L g771 ( .A(n_512), .Y(n_771) );
HB1xp67_ASAP7_75t_L g1245 ( .A(n_512), .Y(n_1245) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
OR2x6_ASAP7_75t_L g522 ( .A(n_513), .B(n_523), .Y(n_522) );
BUFx4f_ASAP7_75t_L g694 ( .A(n_513), .Y(n_694) );
INVxp67_ASAP7_75t_L g949 ( .A(n_513), .Y(n_949) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g654 ( .A(n_519), .Y(n_654) );
INVx3_ASAP7_75t_L g1243 ( .A(n_522), .Y(n_1243) );
INVx3_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g657 ( .A(n_525), .Y(n_657) );
INVx4_ASAP7_75t_L g825 ( .A(n_525), .Y(n_825) );
OAI211xp5_ASAP7_75t_L g1206 ( .A1(n_527), .A2(n_1207), .B(n_1208), .C(n_1210), .Y(n_1206) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g683 ( .A(n_528), .Y(n_683) );
INVx2_ASAP7_75t_L g689 ( .A(n_528), .Y(n_689) );
INVx2_ASAP7_75t_L g753 ( .A(n_528), .Y(n_753) );
INVx2_ASAP7_75t_L g1673 ( .A(n_528), .Y(n_1673) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx4f_ASAP7_75t_L g595 ( .A(n_529), .Y(n_595) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_529), .Y(n_647) );
BUFx4f_ASAP7_75t_L g855 ( .A(n_529), .Y(n_855) );
BUFx4f_ASAP7_75t_L g925 ( .A(n_529), .Y(n_925) );
BUFx4f_ASAP7_75t_L g1236 ( .A(n_529), .Y(n_1236) );
OR2x6_ASAP7_75t_L g1676 ( .A(n_529), .B(n_1677), .Y(n_1676) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g601 ( .A(n_530), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_534), .B1(n_535), .B2(n_537), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_532), .A2(n_535), .B1(n_1239), .B2(n_1240), .Y(n_1238) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_533), .A2(n_536), .B1(n_649), .B2(n_650), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_533), .A2(n_536), .B1(n_1111), .B2(n_1120), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_534), .A2(n_555), .B1(n_559), .B2(n_560), .Y(n_554) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g768 ( .A(n_536), .Y(n_768) );
INVx2_ASAP7_75t_L g985 ( .A(n_536), .Y(n_985) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g906 ( .A(n_539), .Y(n_906) );
INVx1_ASAP7_75t_L g1237 ( .A(n_539), .Y(n_1237) );
AND2x2_ASAP7_75t_L g864 ( .A(n_540), .B(n_865), .Y(n_864) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .C(n_563), .Y(n_541) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g1711 ( .A1(n_544), .A2(n_784), .B1(n_1712), .B2(n_1713), .Y(n_1711) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g875 ( .A(n_545), .Y(n_875) );
INVx1_ASAP7_75t_L g1107 ( .A(n_545), .Y(n_1107) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g671 ( .A(n_547), .Y(n_671) );
INVx2_ASAP7_75t_L g776 ( .A(n_547), .Y(n_776) );
INVx2_ASAP7_75t_L g828 ( .A(n_547), .Y(n_828) );
INVxp67_ASAP7_75t_L g1108 ( .A(n_547), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1703 ( .A1(n_547), .A2(n_662), .B1(n_1704), .B2(n_1705), .Y(n_1703) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_550), .A2(n_718), .B1(n_950), .B2(n_958), .Y(n_970) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g665 ( .A(n_551), .Y(n_665) );
INVx1_ASAP7_75t_L g779 ( .A(n_551), .Y(n_779) );
INVx1_ASAP7_75t_L g932 ( .A(n_551), .Y(n_932) );
INVx2_ASAP7_75t_L g941 ( .A(n_551), .Y(n_941) );
NAND4xp25_ASAP7_75t_L g1702 ( .A(n_552), .B(n_1703), .C(n_1706), .D(n_1711), .Y(n_1702) );
CKINVDCx8_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
CKINVDCx8_ASAP7_75t_R g666 ( .A(n_553), .Y(n_666) );
OAI31xp33_ASAP7_75t_L g1374 ( .A1(n_553), .A2(n_1375), .A3(n_1385), .B(n_1386), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_555), .A2(n_560), .B1(n_1239), .B2(n_1282), .Y(n_1281) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g899 ( .A(n_556), .Y(n_899) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x4_ASAP7_75t_L g561 ( .A(n_557), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g668 ( .A(n_557), .B(n_558), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g1375 ( .A1(n_557), .A2(n_1376), .B(n_1379), .C(n_1382), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_560), .A2(n_899), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
AOI222xp33_ASAP7_75t_L g1706 ( .A1(n_560), .A2(n_899), .B1(n_1707), .B2(n_1708), .C1(n_1709), .C2(n_1710), .Y(n_1706) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_561), .A2(n_649), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_561), .A2(n_668), .B1(n_766), .B2(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_561), .A2(n_668), .B1(n_820), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_561), .A2(n_668), .B1(n_868), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_561), .A2(n_899), .B1(n_900), .B2(n_901), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_561), .A2(n_668), .B1(n_975), .B2(n_976), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_561), .A2(n_668), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1382 ( .A1(n_561), .A2(n_668), .B1(n_1383), .B2(n_1384), .Y(n_1382) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_SL g784 ( .A(n_565), .Y(n_784) );
BUFx3_ASAP7_75t_L g903 ( .A(n_565), .Y(n_903) );
BUFx2_ASAP7_75t_L g1326 ( .A(n_565), .Y(n_1326) );
BUFx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g662 ( .A(n_567), .Y(n_662) );
INVx1_ASAP7_75t_L g786 ( .A(n_567), .Y(n_786) );
INVx1_ASAP7_75t_L g879 ( .A(n_567), .Y(n_879) );
INVx1_ASAP7_75t_L g728 ( .A(n_568), .Y(n_728) );
BUFx3_ASAP7_75t_L g1307 ( .A(n_568), .Y(n_1307) );
CKINVDCx14_ASAP7_75t_R g569 ( .A(n_570), .Y(n_569) );
OAI31xp33_ASAP7_75t_L g774 ( .A1(n_570), .A2(n_775), .A3(n_777), .B(n_782), .Y(n_774) );
OAI31xp33_ASAP7_75t_L g894 ( .A1(n_570), .A2(n_895), .A3(n_896), .B(n_902), .Y(n_894) );
AOI211xp5_ASAP7_75t_L g1701 ( .A1(n_570), .A2(n_1702), .B(n_1714), .C(n_1729), .Y(n_1701) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
AND2x2_ASAP7_75t_L g672 ( .A(n_571), .B(n_573), .Y(n_672) );
AND2x2_ASAP7_75t_L g978 ( .A(n_571), .B(n_573), .Y(n_978) );
AND2x2_ASAP7_75t_SL g1284 ( .A(n_571), .B(n_573), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_571), .B(n_573), .Y(n_1386) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_611), .Y(n_575) );
OAI33xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .A3(n_590), .B1(n_597), .B2(n_603), .B3(n_608), .Y(n_576) );
OAI33xp33_ASAP7_75t_L g674 ( .A1(n_577), .A2(n_675), .A3(n_679), .B1(n_684), .B2(n_691), .B3(n_693), .Y(n_674) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g745 ( .A(n_578), .Y(n_745) );
INVx4_ASAP7_75t_L g812 ( .A(n_578), .Y(n_812) );
INVx2_ASAP7_75t_L g856 ( .A(n_578), .Y(n_856) );
INVx1_ASAP7_75t_L g1270 ( .A(n_578), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_585), .B2(n_586), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_581), .A2(n_598), .B1(n_616), .B2(n_619), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_582), .A2(n_586), .B1(n_609), .B2(n_610), .Y(n_608) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_585), .A2(n_602), .B1(n_633), .B2(n_635), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_586), .A2(n_1251), .B1(n_1267), .B2(n_1272), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_586), .A2(n_1259), .B1(n_1263), .B2(n_1272), .Y(n_1277) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_588), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_588), .A2(n_677), .B1(n_839), .B2(n_849), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_588), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1171) );
INVx4_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_589), .Y(n_697) );
INVx2_ASAP7_75t_L g757 ( .A(n_589), .Y(n_757) );
INVx2_ASAP7_75t_SL g951 ( .A(n_589), .Y(n_951) );
INVx2_ASAP7_75t_L g1085 ( .A(n_589), .Y(n_1085) );
INVx1_ASAP7_75t_L g1311 ( .A(n_589), .Y(n_1311) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_591), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g1275 ( .A1(n_591), .A2(n_595), .B1(n_1257), .B2(n_1262), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_591), .A2(n_595), .B1(n_1253), .B2(n_1268), .Y(n_1276) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g752 ( .A(n_592), .Y(n_752) );
INVx2_ASAP7_75t_L g1156 ( .A(n_592), .Y(n_1156) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx2_ASAP7_75t_L g681 ( .A(n_593), .Y(n_681) );
BUFx2_ASAP7_75t_L g687 ( .A(n_593), .Y(n_687) );
INVx1_ASAP7_75t_L g749 ( .A(n_593), .Y(n_749) );
BUFx3_ASAP7_75t_L g921 ( .A(n_593), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_594), .A2(n_609), .B1(n_623), .B2(n_626), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_596), .A2(n_610), .B1(n_629), .B2(n_631), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_599), .A2(n_748), .B1(n_957), .B2(n_958), .Y(n_956) );
OAI211xp5_ASAP7_75t_L g1042 ( .A1(n_599), .A2(n_1043), .B(n_1044), .C(n_1047), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_599), .A2(n_685), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_599), .A2(n_685), .B1(n_1296), .B2(n_1306), .Y(n_1312) );
INVx5_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
BUFx3_ASAP7_75t_L g763 ( .A(n_601), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_601), .B(n_1166), .Y(n_1165) );
BUFx2_ASAP7_75t_SL g1315 ( .A(n_601), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1660 ( .A(n_601), .B(n_1659), .Y(n_1660) );
OAI33xp33_ASAP7_75t_L g1269 ( .A1(n_603), .A2(n_1270), .A3(n_1271), .B1(n_1275), .B2(n_1276), .B3(n_1277), .Y(n_1269) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI33xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .A3(n_622), .B1(n_628), .B2(n_632), .B3(n_636), .Y(n_611) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g700 ( .A(n_613), .Y(n_700) );
BUFx8_ASAP7_75t_L g715 ( .A(n_613), .Y(n_715) );
BUFx4f_ASAP7_75t_L g1249 ( .A(n_613), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1624 ( .A(n_614), .Y(n_1624) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_618), .A2(n_703), .B1(n_1227), .B2(n_1228), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_619), .A2(n_717), .B1(n_718), .B2(n_721), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_619), .A2(n_1252), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_619), .A2(n_702), .B1(n_1300), .B2(n_1301), .Y(n_1299) );
OAI22xp33_ASAP7_75t_L g1302 ( .A1(n_619), .A2(n_850), .B1(n_1303), .B2(n_1304), .Y(n_1302) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g881 ( .A(n_620), .Y(n_881) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_621), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_621), .A2(n_678), .B1(n_690), .B2(n_702), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g1715 ( .A1(n_623), .A2(n_733), .B1(n_1716), .B2(n_1717), .C(n_1718), .Y(n_1715) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g706 ( .A(n_625), .Y(n_706) );
INVx3_ASAP7_75t_L g967 ( .A(n_625), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_626), .A2(n_1257), .B1(n_1258), .B2(n_1259), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_626), .A2(n_1261), .B1(n_1262), .B2(n_1263), .Y(n_1260) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g631 ( .A(n_627), .Y(n_631) );
INVx1_ASAP7_75t_L g707 ( .A(n_627), .Y(n_707) );
CKINVDCx8_ASAP7_75t_R g733 ( .A(n_627), .Y(n_733) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_631), .A2(n_682), .B1(n_698), .B2(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_631), .A2(n_706), .B1(n_799), .B2(n_800), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_631), .A2(n_709), .B1(n_846), .B2(n_847), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_631), .A2(n_1087), .B1(n_1093), .B2(n_1101), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1721 ( .A1(n_631), .A2(n_706), .B1(n_1722), .B2(n_1723), .C(n_1724), .Y(n_1721) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g1252 ( .A(n_634), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g1714 ( .A1(n_636), .A2(n_1248), .B1(n_1715), .B2(n_1721), .Y(n_1714) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_637), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g1066 ( .A(n_637), .B(n_1067), .C(n_1069), .Y(n_1066) );
INVx2_ASAP7_75t_L g1373 ( .A(n_637), .Y(n_1373) );
INVx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g939 ( .A(n_638), .Y(n_939) );
OAI33xp33_ASAP7_75t_L g962 ( .A1(n_638), .A2(n_715), .A3(n_963), .B1(n_965), .B2(n_968), .B3(n_970), .Y(n_962) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_787), .B1(n_884), .B2(n_885), .Y(n_641) );
INVx1_ASAP7_75t_L g884 ( .A(n_642), .Y(n_884) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_711), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_659), .C(n_673), .Y(n_644) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_651), .A3(n_655), .B(n_658), .Y(n_645) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_647), .A2(n_723), .B1(n_730), .B2(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g772 ( .A(n_654), .Y(n_772) );
INVx1_ASAP7_75t_L g1122 ( .A(n_654), .Y(n_1122) );
INVx1_ASAP7_75t_L g1117 ( .A(n_656), .Y(n_1117) );
OAI31xp33_ASAP7_75t_L g904 ( .A1(n_658), .A2(n_905), .A3(n_909), .B(n_910), .Y(n_904) );
OAI31xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .A3(n_670), .B(n_672), .Y(n_659) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI31xp33_ASAP7_75t_L g826 ( .A1(n_672), .A2(n_827), .A3(n_829), .B(n_832), .Y(n_826) );
OAI31xp33_ASAP7_75t_SL g872 ( .A1(n_672), .A2(n_873), .A3(n_876), .B(n_880), .Y(n_872) );
OAI31xp33_ASAP7_75t_L g1104 ( .A1(n_672), .A2(n_1105), .A3(n_1109), .B(n_1113), .Y(n_1104) );
NOR2xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_699), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_676), .A2(n_688), .B1(n_702), .B2(n_703), .Y(n_701) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B1(n_682), .B2(n_683), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_680), .A2(n_695), .B1(n_706), .B2(n_707), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_681), .A2(n_763), .B1(n_799), .B2(n_802), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_681), .A2(n_763), .B1(n_795), .B2(n_808), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_681), .A2(n_843), .B1(n_846), .B2(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g1202 ( .A(n_683), .B(n_1203), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_685), .A2(n_689), .B1(n_840), .B2(n_851), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_685), .A2(n_924), .B1(n_925), .B2(n_926), .Y(n_923) );
INVx4_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g954 ( .A(n_686), .Y(n_954) );
INVx2_ASAP7_75t_L g1314 ( .A(n_686), .Y(n_1314) );
INVx4_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI33xp33_ASAP7_75t_L g809 ( .A1(n_691), .A2(n_810), .A3(n_813), .B1(n_814), .B2(n_815), .B3(n_816), .Y(n_809) );
OAI33xp33_ASAP7_75t_L g853 ( .A1(n_691), .A2(n_854), .A3(n_856), .B1(n_857), .B2(n_858), .B3(n_859), .Y(n_853) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_696), .B2(n_698), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_694), .A2(n_696), .B1(n_928), .B2(n_929), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_694), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1310 ( .A1(n_694), .A2(n_1300), .B1(n_1303), .B2(n_1311), .Y(n_1310) );
INVx5_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx6_ASAP7_75t_L g1317 ( .A(n_697), .Y(n_1317) );
BUFx4f_ASAP7_75t_SL g794 ( .A(n_702), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_702), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_702), .A2(n_779), .B1(n_1082), .B2(n_1090), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_702), .A2(n_796), .B1(n_1083), .B2(n_1091), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_703), .Y(n_897) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_706), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_706), .A2(n_707), .B1(n_843), .B2(n_844), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_758), .C(n_774), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_743), .Y(n_713) );
OAI33xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .A3(n_722), .B1(n_729), .B2(n_734), .B3(n_735), .Y(n_714) );
OAI33xp33_ASAP7_75t_L g930 ( .A1(n_715), .A2(n_931), .A3(n_933), .B1(n_936), .B2(n_937), .B3(n_940), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_718), .A2(n_947), .B1(n_957), .B2(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g737 ( .A(n_720), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_721), .A2(n_742), .B1(n_751), .B2(n_753), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_726), .A2(n_918), .B1(n_928), .B2(n_934), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_726), .A2(n_955), .B1(n_961), .B2(n_969), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_726), .A2(n_1058), .B1(n_1059), .B2(n_1060), .C(n_1061), .Y(n_1057) );
OAI22xp33_ASAP7_75t_SL g1295 ( .A1(n_726), .A2(n_1296), .B1(n_1297), .B2(n_1298), .Y(n_1295) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_731), .A2(n_1306), .B1(n_1307), .B2(n_1308), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_733), .A2(n_953), .B1(n_960), .B2(n_966), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_733), .A2(n_1058), .B1(n_1088), .B2(n_1097), .Y(n_1103) );
OAI221xp5_ASAP7_75t_L g1362 ( .A1(n_733), .A2(n_1363), .B1(n_1364), .B2(n_1365), .C(n_1366), .Y(n_1362) );
OAI221xp5_ASAP7_75t_L g1369 ( .A1(n_733), .A2(n_966), .B1(n_1351), .B2(n_1370), .C(n_1371), .Y(n_1369) );
OAI33xp33_ASAP7_75t_L g1294 ( .A1(n_734), .A2(n_1248), .A3(n_1295), .B1(n_1299), .B2(n_1302), .B3(n_1305), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B1(n_739), .B2(n_742), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_736), .A2(n_914), .B1(n_924), .B2(n_932), .Y(n_931) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_736), .A2(n_916), .B1(n_926), .B2(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_740), .Y(n_852) );
INVx1_ASAP7_75t_L g964 ( .A(n_740), .Y(n_964) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g797 ( .A(n_741), .Y(n_797) );
OR2x6_ASAP7_75t_L g1636 ( .A(n_741), .B(n_1637), .Y(n_1636) );
OAI33xp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_746), .A3(n_747), .B1(n_750), .B2(n_754), .B3(n_756), .Y(n_743) );
OAI33xp33_ASAP7_75t_L g945 ( .A1(n_744), .A2(n_754), .A3(n_946), .B1(n_952), .B2(n_956), .B3(n_959), .Y(n_945) );
OAI21xp5_ASAP7_75t_L g1670 ( .A1(n_744), .A2(n_1671), .B(n_1676), .Y(n_1670) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx4_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI211xp5_ASAP7_75t_L g1211 ( .A1(n_753), .A2(n_1212), .B(n_1213), .C(n_1214), .Y(n_1211) );
OAI33xp33_ASAP7_75t_L g912 ( .A1(n_754), .A2(n_810), .A3(n_913), .B1(n_917), .B2(n_923), .B3(n_927), .Y(n_912) );
OAI33xp33_ASAP7_75t_L g1080 ( .A1(n_754), .A2(n_810), .A3(n_1081), .B1(n_1086), .B2(n_1089), .B3(n_1092), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g1318 ( .A(n_755), .Y(n_1318) );
AOI211xp5_ASAP7_75t_L g1664 ( .A1(n_755), .A2(n_1665), .B(n_1670), .C(n_1680), .Y(n_1664) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_757), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_757), .A2(n_1093), .B1(n_1094), .B2(n_1097), .Y(n_1092) );
OAI31xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .A3(n_770), .B(n_773), .Y(n_758) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI211xp5_ASAP7_75t_L g1735 ( .A1(n_763), .A2(n_1736), .B(n_1737), .C(n_1738), .Y(n_1735) );
OAI211xp5_ASAP7_75t_SL g1739 ( .A1(n_763), .A2(n_1722), .B(n_1740), .C(n_1741), .Y(n_1739) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_767), .B2(n_769), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_765), .A2(n_820), .B1(n_821), .B2(n_822), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_765), .A2(n_821), .B1(n_868), .B2(n_869), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_765), .A2(n_767), .B1(n_900), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_765), .A2(n_975), .B1(n_984), .B2(n_986), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_765), .A2(n_984), .B1(n_1323), .B2(n_1333), .Y(n_1332) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g821 ( .A(n_768), .Y(n_821) );
OAI31xp33_ASAP7_75t_L g979 ( .A1(n_773), .A2(n_980), .A3(n_981), .B(n_987), .Y(n_979) );
OAI31xp33_ASAP7_75t_L g1327 ( .A1(n_773), .A2(n_1328), .A3(n_1329), .B(n_1334), .Y(n_1327) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g877 ( .A(n_784), .Y(n_877) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g885 ( .A(n_787), .Y(n_885) );
XOR2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_833), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_817), .C(n_826), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_809), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_792) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_794), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_794), .A2(n_941), .B1(n_1212), .B2(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g841 ( .A(n_797), .Y(n_841) );
INVx1_ASAP7_75t_L g1255 ( .A(n_807), .Y(n_1255) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
XNOR2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
AND3x1_ASAP7_75t_L g835 ( .A(n_836), .B(n_860), .C(n_872), .Y(n_835) );
NOR2xp33_ASAP7_75t_SL g836 ( .A(n_837), .B(n_853), .Y(n_836) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_855), .A2(n_918), .B1(n_919), .B2(n_922), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_855), .A2(n_953), .B1(n_954), .B2(n_955), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_855), .A2(n_954), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
INVx1_ASAP7_75t_L g1331 ( .A(n_855), .Y(n_1331) );
OAI31xp33_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_862), .A3(n_870), .B(n_871), .Y(n_860) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g982 ( .A(n_864), .Y(n_982) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_866), .Y(n_1039) );
OAI31xp33_ASAP7_75t_SL g1114 ( .A1(n_871), .A2(n_1115), .A3(n_1118), .B(n_1121), .Y(n_1114) );
INVx2_ASAP7_75t_SL g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_1180), .B2(n_1181), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
XNOR2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_988), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
XNOR2x1_ASAP7_75t_L g891 ( .A(n_892), .B(n_942), .Y(n_891) );
NAND3xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_904), .C(n_911), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_930), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_915), .A2(n_1298), .B1(n_1308), .B2(n_1317), .Y(n_1316) );
OAI221xp5_ASAP7_75t_L g1671 ( .A1(n_919), .A2(n_1672), .B1(n_1673), .B2(n_1674), .C(n_1675), .Y(n_1671) );
INVx3_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
OAI211xp5_ASAP7_75t_SL g1346 ( .A1(n_925), .A2(n_1347), .B(n_1348), .C(n_1349), .Y(n_1346) );
OAI211xp5_ASAP7_75t_SL g1350 ( .A1(n_925), .A2(n_1351), .B(n_1352), .C(n_1354), .Y(n_1350) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_SL g1363 ( .A(n_935), .Y(n_1363) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_939), .Y(n_1265) );
NAND3xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_971), .C(n_979), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_962), .Y(n_944) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_948), .B1(n_950), .B2(n_951), .Y(n_946) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
OAI31xp33_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .A3(n_977), .B(n_978), .Y(n_971) );
OAI31xp33_ASAP7_75t_L g1319 ( .A1(n_978), .A2(n_1320), .A3(n_1321), .B(n_1325), .Y(n_1319) );
INVx2_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
XNOR2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_1075), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1073 ( .A(n_991), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_995), .C(n_1009), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_993), .A2(n_1051), .B1(n_1052), .B2(n_1053), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_997), .B1(n_1002), .B2(n_1003), .Y(n_995) );
INVxp67_ASAP7_75t_L g1188 ( .A(n_997), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_1001), .Y(n_997) );
INVx3_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_1000), .B(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1003), .Y(n_1189) );
NAND2x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1006), .Y(n_1003) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1663 ( .A(n_1007), .Y(n_1663) );
NOR3xp33_ASAP7_75t_SL g1009 ( .A(n_1010), .B(n_1020), .C(n_1056), .Y(n_1009) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1017), .B1(n_1018), .B2(n_1019), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_1016), .B(n_1032), .Y(n_1031) );
AOI222xp33_ASAP7_75t_L g1127 ( .A1(n_1017), .A2(n_1019), .B1(n_1128), .B2(n_1129), .C1(n_1131), .C2(n_1132), .Y(n_1127) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_1018), .A2(n_1034), .B1(n_1036), .B2(n_1037), .C(n_1038), .Y(n_1033) );
AOI31xp33_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1042), .A3(n_1050), .B(n_1054), .Y(n_1020) );
AOI21xp5_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1027), .B(n_1030), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1023 ( .A(n_1024), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1160 ( .A1(n_1025), .A2(n_1143), .B1(n_1147), .B2(n_1161), .C(n_1163), .Y(n_1160) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1033), .B(n_1040), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_1034), .A2(n_1194), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1034), .Y(n_1360) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1036), .Y(n_1359) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
A2O1A1Ixp33_ASAP7_75t_L g1164 ( .A1(n_1041), .A2(n_1132), .B(n_1152), .C(n_1165), .Y(n_1164) );
A2O1A1Ixp33_ASAP7_75t_L g1199 ( .A1(n_1041), .A2(n_1200), .B(n_1201), .C(n_1202), .Y(n_1199) );
A2O1A1Ixp33_ASAP7_75t_SL g1356 ( .A1(n_1041), .A2(n_1201), .B(n_1357), .C(n_1358), .Y(n_1356) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1051), .Y(n_1216) );
AOI21xp5_ASAP7_75t_L g1616 ( .A1(n_1054), .A2(n_1617), .B(n_1651), .Y(n_1616) );
BUFx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
BUFx2_ASAP7_75t_L g1627 ( .A(n_1064), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_1068), .A2(n_1357), .B1(n_1377), .B2(n_1378), .Y(n_1376) );
INVx3_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1071), .Y(n_1130) );
INVx8_ASAP7_75t_L g1135 ( .A(n_1071), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_1071), .Y(n_1367) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1071), .Y(n_1647) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1077), .B1(n_1123), .B2(n_1179), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_1077), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1104), .C(n_1114), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1098), .Y(n_1079) );
BUFx6f_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx3_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
BUFx6f_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx4_ASAP7_75t_L g1173 ( .A(n_1096), .Y(n_1173) );
INVx3_ASAP7_75t_L g1274 ( .A(n_1096), .Y(n_1274) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1124), .Y(n_1179) );
XNOR2x1_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1178), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1144), .Y(n_1125) );
NAND3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1133), .C(n_1142), .Y(n_1126) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NAND3xp33_ASAP7_75t_SL g1144 ( .A(n_1145), .B(n_1148), .C(n_1175), .Y(n_1144) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx3_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
BUFx6f_ASAP7_75t_L g1201 ( .A(n_1152), .Y(n_1201) );
OAI21xp33_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1160), .B(n_1164), .Y(n_1157) );
INVxp67_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OAI21xp5_ASAP7_75t_L g1343 ( .A1(n_1159), .A2(n_1344), .B(n_1345), .Y(n_1343) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1287), .B1(n_1288), .B2(n_1387), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
HB1xp67_ASAP7_75t_L g1387 ( .A(n_1183), .Y(n_1387) );
AO22x2_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1230), .B1(n_1231), .B2(n_1286), .Y(n_1183) );
INVx1_ASAP7_75t_SL g1286 ( .A(n_1184), .Y(n_1286) );
XNOR2x1_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .Y(n_1184) );
NOR2x1_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1190), .Y(n_1186) );
NAND3xp33_ASAP7_75t_SL g1190 ( .A(n_1191), .B(n_1197), .C(n_1219), .Y(n_1190) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
OAI21xp5_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1215), .B(n_1218), .Y(n_1197) );
NAND3xp33_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1206), .C(n_1211), .Y(n_1198) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NAND3xp33_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1246), .C(n_1278), .Y(n_1233) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1243), .B(n_1398), .Y(n_1397) );
AND2x4_ASAP7_75t_SL g1688 ( .A(n_1243), .B(n_1689), .Y(n_1688) );
NOR2xp33_ASAP7_75t_SL g1246 ( .A(n_1247), .B(n_1269), .Y(n_1246) );
OAI33xp33_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1250), .A3(n_1256), .B1(n_1260), .B2(n_1264), .B3(n_1266), .Y(n_1247) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_1248), .A2(n_1362), .B1(n_1369), .B2(n_1373), .Y(n_1361) );
BUFx3_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1250) );
INVx2_ASAP7_75t_SL g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
OAI33xp33_ASAP7_75t_L g1309 ( .A1(n_1270), .A2(n_1310), .A3(n_1312), .B1(n_1313), .B2(n_1316), .B3(n_1318), .Y(n_1309) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx2_ASAP7_75t_SL g1273 ( .A(n_1274), .Y(n_1273) );
OAI22xp33_ASAP7_75t_L g1667 ( .A1(n_1274), .A2(n_1317), .B1(n_1668), .B2(n_1669), .Y(n_1667) );
OAI31xp33_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1280), .A3(n_1283), .B(n_1284), .Y(n_1278) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1290), .B1(n_1335), .B2(n_1336), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1319), .C(n_1327), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1309), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_1301), .A2(n_1304), .B1(n_1314), .B2(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
XNOR2x1_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1374), .Y(n_1339) );
AOI21xp5_ASAP7_75t_L g1340 ( .A1(n_1341), .A2(n_1342), .B(n_1361), .Y(n_1340) );
NAND4xp25_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1346), .C(n_1350), .D(n_1356), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1645 ( .A1(n_1372), .A2(n_1646), .B1(n_1647), .B2(n_1648), .Y(n_1645) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1396), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1394), .Y(n_1391) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1392), .B(n_1395), .Y(n_1693) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1392), .Y(n_1751) );
HB1xp67_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
NOR2xp33_ASAP7_75t_L g1753 ( .A(n_1395), .B(n_1751), .Y(n_1753) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1610), .B1(n_1613), .B2(n_1686), .C(n_1690), .Y(n_1399) );
AOI21xp5_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1523), .B(n_1567), .Y(n_1400) );
OAI211xp5_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1417), .B(n_1463), .C(n_1509), .Y(n_1401) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_1402), .A2(n_1515), .B1(n_1593), .B2(n_1599), .Y(n_1592) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_1403), .Y(n_1402) );
CKINVDCx6p67_ASAP7_75t_R g1475 ( .A(n_1403), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1403), .B(n_1435), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1594 ( .A(n_1403), .B(n_1435), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1609 ( .A(n_1403), .B(n_1499), .Y(n_1609) );
OR2x6_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1411), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1496 ( .A(n_1404), .B(n_1411), .Y(n_1496) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1405), .Y(n_1506) );
AND2x6_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1407), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1406), .B(n_1410), .Y(n_1409) );
AND2x4_ASAP7_75t_L g1412 ( .A(n_1406), .B(n_1413), .Y(n_1412) );
AND2x6_ASAP7_75t_L g1415 ( .A(n_1406), .B(n_1416), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1406), .B(n_1410), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1406), .B(n_1410), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1408), .B(n_1414), .Y(n_1413) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1415), .Y(n_1612) );
HB1xp67_ASAP7_75t_L g1750 ( .A(n_1416), .Y(n_1750) );
O2A1O1Ixp33_ASAP7_75t_L g1417 ( .A1(n_1418), .A2(n_1433), .B(n_1438), .C(n_1452), .Y(n_1417) );
NOR2xp33_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1423), .Y(n_1418) );
INVx2_ASAP7_75t_L g1446 ( .A(n_1419), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1419), .B(n_1454), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1419), .B(n_1428), .Y(n_1460) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1419), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1419), .B(n_1491), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1533 ( .A(n_1419), .B(n_1495), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1419), .B(n_1448), .Y(n_1565) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1419), .B(n_1448), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1421), .Y(n_1419) );
INVxp67_ASAP7_75t_L g1508 ( .A(n_1422), .Y(n_1508) );
OR2x2_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1428), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1424), .B(n_1457), .Y(n_1462) );
AND3x1_ASAP7_75t_L g1479 ( .A(n_1424), .B(n_1440), .C(n_1445), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1424), .B(n_1440), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1424), .B(n_1428), .Y(n_1598) );
INVx2_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1425), .B(n_1440), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1425), .B(n_1457), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1425), .B(n_1428), .Y(n_1495) );
OR2x2_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1427), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1428), .B(n_1457), .Y(n_1456) );
OR2x2_ASAP7_75t_L g1481 ( .A(n_1428), .B(n_1440), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1428), .B(n_1486), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1428), .B(n_1440), .Y(n_1563) );
BUFx2_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
INVx2_ASAP7_75t_L g1445 ( .A(n_1429), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1429), .B(n_1439), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1429), .B(n_1462), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1429), .B(n_1470), .Y(n_1530) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1429), .B(n_1552), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1431), .Y(n_1429) );
O2A1O1Ixp33_ASAP7_75t_L g1438 ( .A1(n_1433), .A2(n_1439), .B(n_1443), .C(n_1447), .Y(n_1438) );
CKINVDCx14_ASAP7_75t_R g1433 ( .A(n_1434), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_1434), .A2(n_1514), .B1(n_1517), .B2(n_1520), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1534 ( .A(n_1434), .B(n_1502), .Y(n_1534) );
AOI211xp5_ASAP7_75t_L g1558 ( .A1(n_1434), .A2(n_1559), .B(n_1560), .C(n_1561), .Y(n_1558) );
AOI221xp5_ASAP7_75t_L g1568 ( .A1(n_1434), .A2(n_1479), .B1(n_1569), .B2(n_1571), .C(n_1572), .Y(n_1568) );
INVx3_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1435), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1465 ( .A(n_1435), .B(n_1448), .Y(n_1465) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_1435), .A2(n_1490), .B1(n_1493), .B2(n_1494), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1435), .B(n_1448), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1435), .B(n_1454), .Y(n_1500) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1435), .B(n_1475), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1435), .B(n_1565), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1435), .B(n_1475), .Y(n_1591) );
AND2x4_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1437), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1439), .B(n_1446), .Y(n_1513) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1439), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1439), .B(n_1460), .Y(n_1596) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1440), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1440), .B(n_1445), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1442), .Y(n_1440) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1444), .B(n_1462), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1446), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1445), .B(n_1470), .Y(n_1469) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_1445), .B(n_1513), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1445), .B(n_1462), .Y(n_1555) );
OR2x2_ASAP7_75t_L g1604 ( .A(n_1445), .B(n_1522), .Y(n_1604) );
NAND2xp5_ASAP7_75t_SL g1606 ( .A(n_1445), .B(n_1607), .Y(n_1606) );
NOR2xp33_ASAP7_75t_L g1484 ( .A(n_1446), .B(n_1485), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1519 ( .A(n_1446), .B(n_1481), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1446), .B(n_1474), .Y(n_1529) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1446), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1446), .B(n_1563), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1447), .B(n_1475), .Y(n_1482) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1447), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1451), .Y(n_1447) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1448), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1450), .Y(n_1448) );
OAI21xp33_ASAP7_75t_L g1452 ( .A1(n_1453), .A2(n_1455), .B(n_1458), .Y(n_1452) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1454), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1454), .B(n_1475), .Y(n_1487) );
OAI211xp5_ASAP7_75t_SL g1525 ( .A1(n_1455), .A2(n_1526), .B(n_1527), .C(n_1531), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g1550 ( .A(n_1455), .B(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
A2O1A1Ixp33_ASAP7_75t_L g1483 ( .A1(n_1456), .A2(n_1468), .B(n_1484), .C(n_1487), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g1509 ( .A1(n_1456), .A2(n_1510), .B1(n_1511), .B2(n_1514), .C(n_1516), .Y(n_1509) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1458), .Y(n_1559) );
OR2x2_ASAP7_75t_L g1586 ( .A(n_1458), .B(n_1474), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1461), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1462), .B(n_1468), .Y(n_1522) );
AOI211xp5_ASAP7_75t_L g1463 ( .A1(n_1464), .A2(n_1466), .B(n_1471), .C(n_1488), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1464), .B(n_1468), .Y(n_1510) );
OAI322xp33_ASAP7_75t_L g1537 ( .A1(n_1464), .A2(n_1481), .A3(n_1496), .B1(n_1513), .B2(n_1538), .C1(n_1541), .C2(n_1543), .Y(n_1537) );
AND2x2_ASAP7_75t_SL g1560 ( .A(n_1464), .B(n_1479), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1464), .B(n_1467), .Y(n_1570) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1469), .Y(n_1466) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_1467), .B(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1467), .Y(n_1542) );
AOI31xp33_ASAP7_75t_L g1549 ( .A1(n_1467), .A2(n_1545), .A3(n_1550), .B(n_1553), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1467), .B(n_1479), .Y(n_1590) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
NAND2xp5_ASAP7_75t_SL g1526 ( .A(n_1468), .B(n_1493), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1468), .B(n_1548), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1469), .B(n_1542), .Y(n_1541) );
OR2x2_ASAP7_75t_L g1607 ( .A(n_1470), .B(n_1486), .Y(n_1607) );
OAI211xp5_ASAP7_75t_L g1471 ( .A1(n_1472), .A2(n_1476), .B(n_1478), .C(n_1483), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1475), .Y(n_1473) );
INVx2_ASAP7_75t_L g1515 ( .A(n_1474), .Y(n_1515) );
A2O1A1Ixp33_ASAP7_75t_L g1587 ( .A1(n_1474), .A2(n_1588), .B(n_1590), .C(n_1591), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1535 ( .A(n_1475), .B(n_1536), .Y(n_1535) );
NOR2xp33_ASAP7_75t_SL g1539 ( .A(n_1475), .B(n_1540), .Y(n_1539) );
NOR2xp33_ASAP7_75t_L g1581 ( .A(n_1475), .B(n_1582), .Y(n_1581) );
O2A1O1Ixp33_ASAP7_75t_L g1572 ( .A1(n_1476), .A2(n_1573), .B(n_1574), .C(n_1575), .Y(n_1572) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
OAI21xp33_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1480), .B(n_1482), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1482), .B(n_1498), .Y(n_1566) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1487), .Y(n_1543) );
OAI221xp5_ASAP7_75t_L g1488 ( .A1(n_1489), .A2(n_1496), .B1(n_1497), .B2(n_1499), .C(n_1501), .Y(n_1488) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
AOI22xp5_ASAP7_75t_L g1577 ( .A1(n_1496), .A2(n_1578), .B1(n_1583), .B2(n_1585), .Y(n_1577) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
CKINVDCx6p67_ASAP7_75t_R g1499 ( .A(n_1500), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1500), .B(n_1557), .Y(n_1556) );
INVx3_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVx2_ASAP7_75t_SL g1502 ( .A(n_1503), .Y(n_1502) );
OAI21xp33_ASAP7_75t_L g1531 ( .A1(n_1503), .A2(n_1532), .B(n_1534), .Y(n_1531) );
INVx2_ASAP7_75t_SL g1536 ( .A(n_1503), .Y(n_1536) );
OAI22xp5_ASAP7_75t_SL g1504 ( .A1(n_1505), .A2(n_1506), .B1(n_1507), .B2(n_1508), .Y(n_1504) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1510), .Y(n_1579) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1514), .B(n_1519), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1514), .B(n_1559), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1514), .B(n_1601), .Y(n_1600) );
INVx2_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
NAND5xp2_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1544), .C(n_1549), .D(n_1558), .E(n_1566), .Y(n_1523) );
AOI21xp5_ASAP7_75t_L g1524 ( .A1(n_1525), .A2(n_1535), .B(n_1537), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1530), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
NAND3xp33_ASAP7_75t_L g1588 ( .A(n_1533), .B(n_1554), .C(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1547), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g1593 ( .A1(n_1546), .A2(n_1594), .B1(n_1595), .B2(n_1597), .Y(n_1593) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1548), .Y(n_1584) );
AOI21xp33_ASAP7_75t_L g1553 ( .A1(n_1552), .A2(n_1554), .B(n_1556), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1554), .B(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVxp67_ASAP7_75t_SL g1561 ( .A(n_1562), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1564), .Y(n_1562) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1563), .Y(n_1573) );
CKINVDCx14_ASAP7_75t_R g1574 ( .A(n_1565), .Y(n_1574) );
NAND5xp2_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1577), .C(n_1587), .D(n_1592), .E(n_1602), .Y(n_1567) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
NAND2xp5_ASAP7_75t_SL g1578 ( .A(n_1579), .B(n_1580), .Y(n_1578) );
INVxp67_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
CKINVDCx14_ASAP7_75t_R g1597 ( .A(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
OAI21xp5_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1605), .B(n_1608), .Y(n_1602) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVxp67_ASAP7_75t_SL g1605 ( .A(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
CKINVDCx20_ASAP7_75t_R g1610 ( .A(n_1611), .Y(n_1610) );
CKINVDCx20_ASAP7_75t_R g1611 ( .A(n_1612), .Y(n_1611) );
BUFx2_ASAP7_75t_SL g1613 ( .A(n_1614), .Y(n_1613) );
AOI21xp5_ASAP7_75t_L g1614 ( .A1(n_1615), .A2(n_1684), .B(n_1685), .Y(n_1614) );
AND3x1_ASAP7_75t_L g1615 ( .A(n_1616), .B(n_1652), .C(n_1664), .Y(n_1615) );
AOI31xp33_ASAP7_75t_L g1685 ( .A1(n_1616), .A2(n_1652), .A3(n_1664), .B(n_1684), .Y(n_1685) );
NAND3xp33_ASAP7_75t_SL g1617 ( .A(n_1618), .B(n_1630), .C(n_1638), .Y(n_1617) );
AOI22xp5_ASAP7_75t_L g1618 ( .A1(n_1619), .A2(n_1621), .B1(n_1625), .B2(n_1626), .Y(n_1618) );
INVx2_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
INVx3_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
AOI221xp5_ASAP7_75t_L g1630 ( .A1(n_1631), .A2(n_1632), .B1(n_1633), .B2(n_1634), .C(n_1635), .Y(n_1630) );
CKINVDCx5p33_ASAP7_75t_R g1635 ( .A(n_1636), .Y(n_1635) );
AOI22xp33_ASAP7_75t_L g1638 ( .A1(n_1639), .A2(n_1643), .B1(n_1649), .B2(n_1650), .Y(n_1638) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
HB1xp67_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1653), .B(n_1661), .Y(n_1652) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVxp67_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1663), .Y(n_1661) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
NAND2x2_ASAP7_75t_L g1681 ( .A(n_1678), .B(n_1682), .Y(n_1681) );
INVx2_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
INVx2_ASAP7_75t_SL g1682 ( .A(n_1683), .Y(n_1682) );
INVx2_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
BUFx3_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
BUFx3_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
BUFx3_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVxp33_ASAP7_75t_SL g1694 ( .A(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
HB1xp67_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1744 ( .A(n_1709), .B(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1710), .Y(n_1728) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
NOR2xp33_ASAP7_75t_L g1730 ( .A(n_1731), .B(n_1733), .Y(n_1730) );
INVx2_ASAP7_75t_SL g1747 ( .A(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
OAI21xp5_ASAP7_75t_L g1749 ( .A1(n_1750), .A2(n_1751), .B(n_1752), .Y(n_1749) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
endmodule