module fake_jpeg_28518_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx8_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_5),
.B(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_15),
.C(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_1),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_12),
.B1(n_25),
.B2(n_18),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_50),
.B(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_12),
.B1(n_25),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_43),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_17),
.B1(n_13),
.B2(n_4),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_27),
.A2(n_17),
.B1(n_13),
.B2(n_4),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_30),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_3),
.B1(n_7),
.B2(n_53),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_13),
.B1(n_3),
.B2(n_7),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_46),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_65),
.B1(n_45),
.B2(n_63),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_49),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_40),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_54),
.B1(n_66),
.B2(n_71),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_42),
.B(n_52),
.Y(n_95)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_67),
.B1(n_70),
.B2(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_83),
.C(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_65),
.B1(n_64),
.B2(n_44),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_69),
.B1(n_64),
.B2(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_86),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_82),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_82),
.B(n_86),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_92),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_94),
.C(n_93),
.Y(n_107)
);

AOI222xp33_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_95),
.B1(n_88),
.B2(n_87),
.C1(n_77),
.C2(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_108),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_91),
.C(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_104),
.B1(n_101),
.B2(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_85),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_100),
.B(n_87),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.C(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_52),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_112),
.C(n_52),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_118),
.B(n_42),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_42),
.Y(n_121)
);


endmodule