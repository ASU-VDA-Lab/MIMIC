module fake_jpeg_7561_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_29),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_23),
.B(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_67),
.B1(n_20),
.B2(n_21),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_18),
.B1(n_27),
.B2(n_47),
.Y(n_85)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_41),
.B1(n_37),
.B2(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_21),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_69),
.B(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_63),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_26),
.B1(n_18),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_97),
.B1(n_53),
.B2(n_48),
.Y(n_111)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_100),
.B1(n_49),
.B2(n_48),
.Y(n_109)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_45),
.A2(n_23),
.B(n_41),
.C(n_37),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_23),
.B(n_19),
.Y(n_102)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AO22x2_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_19),
.B1(n_23),
.B2(n_52),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_106),
.B(n_94),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_63),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_75),
.B(n_96),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_101),
.B1(n_78),
.B2(n_86),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_87),
.B1(n_80),
.B2(n_91),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_90),
.B1(n_99),
.B2(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_82),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_130),
.B1(n_134),
.B2(n_136),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_77),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_140),
.B(n_150),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_68),
.B1(n_71),
.B2(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_144),
.Y(n_155)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

XNOR2x2_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_95),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_116),
.B1(n_112),
.B2(n_113),
.C(n_120),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_154),
.B1(n_123),
.B2(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_98),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_152),
.Y(n_163)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_2),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_14),
.B(n_4),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_3),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_4),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_109),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_161),
.C(n_176),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_110),
.B(n_109),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_160),
.B(n_173),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_110),
.B(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_105),
.C(n_121),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_177),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_134),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_123),
.B(n_103),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_154),
.B1(n_166),
.B2(n_158),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_126),
.C(n_6),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_126),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_133),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_130),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_193),
.C(n_160),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_136),
.B1(n_143),
.B2(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_194),
.B1(n_163),
.B2(n_176),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_151),
.A3(n_143),
.B1(n_147),
.B2(n_150),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_196),
.B(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_141),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_148),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_167),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_192),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_5),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_187),
.B(n_157),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_174),
.B1(n_196),
.B2(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_157),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_170),
.C(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_170),
.C(n_163),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_208),
.C(n_193),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_169),
.C(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_195),
.B1(n_185),
.B2(n_186),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_212),
.B(n_197),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_199),
.B(n_8),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_184),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_223),
.C(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_206),
.B(n_178),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_201),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_172),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_172),
.B1(n_180),
.B2(n_8),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_6),
.C(n_7),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_219),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_204),
.B1(n_211),
.B2(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_225),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_221),
.C(n_217),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_238),
.B(n_231),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_230),
.C(n_8),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_223),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_6),
.C(n_9),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_226),
.B1(n_230),
.B2(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_228),
.B(n_216),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_234),
.B1(n_11),
.B2(n_12),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_SL g248 ( 
.A1(n_246),
.A2(n_9),
.B(n_11),
.Y(n_248)
);

AOI21x1_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_241),
.B(n_11),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_247),
.A2(n_248),
.B(n_9),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_245),
.C(n_13),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_13),
.Y(n_251)
);


endmodule