module fake_jpeg_9023_n_312 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_34),
.B1(n_35),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_51),
.B1(n_65),
.B2(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_55),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_34),
.B1(n_28),
.B2(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_59),
.B1(n_63),
.B2(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_34),
.B1(n_17),
.B2(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_58),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_24),
.B(n_20),
.C(n_30),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_62),
.B(n_66),
.C(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_18),
.B1(n_27),
.B2(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_27),
.B(n_43),
.C(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_44),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_29),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_23),
.B1(n_22),
.B2(n_36),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_23),
.B1(n_31),
.B2(n_36),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_100),
.B(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_3),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_83),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_5),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_5),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_90),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_45),
.B1(n_44),
.B2(n_42),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_48),
.B1(n_54),
.B2(n_53),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_31),
.B1(n_19),
.B2(n_8),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_52),
.B1(n_13),
.B2(n_14),
.Y(n_134)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_6),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_96),
.B(n_103),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_102),
.B(n_105),
.Y(n_111)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_7),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_97),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_7),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_101),
.C(n_106),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_48),
.Y(n_99)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_45),
.A3(n_44),
.B1(n_12),
.B2(n_13),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_46),
.B(n_44),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_8),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_11),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_11),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_50),
.B(n_62),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_88),
.B(n_97),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_123),
.B1(n_130),
.B2(n_132),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_76),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_126),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_76),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_137),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_69),
.B1(n_54),
.B2(n_71),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_134),
.B1(n_109),
.B2(n_106),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_50),
.B1(n_54),
.B2(n_52),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_52),
.B1(n_47),
.B2(n_14),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_90),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_167),
.B(n_137),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_142),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_150),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_145),
.B1(n_113),
.B2(n_131),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_82),
.B1(n_101),
.B2(n_75),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_74),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_148),
.B(n_149),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_79),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_74),
.C(n_105),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_161),
.C(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_92),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_109),
.B1(n_103),
.B2(n_82),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_131),
.B1(n_135),
.B2(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_73),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_170),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_108),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_126),
.B(n_84),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_80),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_85),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_85),
.B(n_94),
.C(n_98),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_85),
.A3(n_83),
.B1(n_93),
.B2(n_89),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_116),
.B(n_85),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_114),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_183),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_190),
.B(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_136),
.B1(n_120),
.B2(n_95),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_188),
.B1(n_202),
.B2(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_136),
.B1(n_120),
.B2(n_95),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_197),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_194),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_136),
.C(n_113),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_206),
.Y(n_230)
);

NAND2xp67_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_145),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_209),
.B1(n_146),
.B2(n_144),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_173),
.B(n_183),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_217),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_194),
.B(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_182),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_214),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_227),
.B1(n_167),
.B2(n_152),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_193),
.B1(n_140),
.B2(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_141),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_177),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_181),
.C(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_238),
.C(n_240),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_185),
.B1(n_202),
.B2(n_172),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_214),
.B1(n_209),
.B2(n_211),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_178),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_248),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_186),
.C(n_172),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_141),
.C(n_179),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_176),
.C(n_175),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_242),
.C(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_249),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_167),
.C(n_193),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_167),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_149),
.C(n_166),
.Y(n_248)
);

OA21x2_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_167),
.B(n_113),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_203),
.B1(n_218),
.B2(n_217),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_266),
.B1(n_213),
.B2(n_205),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_118),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_207),
.B(n_211),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_264),
.B(n_265),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_230),
.B(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_262),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_248),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_216),
.B1(n_215),
.B2(n_227),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_207),
.B(n_223),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_232),
.C(n_235),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_238),
.C(n_244),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_247),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_220),
.C(n_234),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_118),
.C(n_117),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_117),
.C(n_131),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_266),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_288),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_250),
.C(n_258),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_252),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_261),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_277),
.B(n_270),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.C(n_12),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_261),
.B1(n_284),
.B2(n_285),
.Y(n_294)
);

NOR2x1_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_15),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_269),
.B(n_99),
.C(n_14),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_299),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_303),
.B(n_304),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_296),
.B(n_292),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_15),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_297),
.C(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_299),
.B(n_86),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_307),
.B(n_86),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_86),
.Y(n_312)
);


endmodule