module fake_jpeg_19651_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_35),
.B(n_23),
.C(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_56),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_37),
.B1(n_20),
.B2(n_36),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_27),
.C(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_34),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_33),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_29),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_66),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_37),
.B1(n_21),
.B2(n_43),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_72),
.B1(n_92),
.B2(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_70),
.B(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_56),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_37),
.B(n_36),
.C(n_43),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_76),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_88),
.B1(n_30),
.B2(n_28),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_89),
.Y(n_125)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_94),
.B1(n_98),
.B2(n_53),
.Y(n_115)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_93),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_39),
.B1(n_38),
.B2(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_17),
.B1(n_24),
.B2(n_26),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_25),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_23),
.A3(n_35),
.B1(n_24),
.B2(n_26),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_30),
.B1(n_32),
.B2(n_28),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_27),
.B(n_33),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_53),
.B1(n_39),
.B2(n_38),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_117),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_88),
.Y(n_146)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_35),
.B1(n_50),
.B2(n_32),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_40),
.B1(n_28),
.B2(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_85),
.Y(n_144)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_65),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_126),
.B1(n_85),
.B2(n_79),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_92),
.CI(n_72),
.CON(n_140),
.SN(n_140)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_64),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_134),
.C(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_63),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_135),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_64),
.C(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_64),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_152),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_84),
.B(n_77),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_140),
.B(n_144),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_100),
.C(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_95),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_146),
.B1(n_157),
.B2(n_110),
.Y(n_168)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_27),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_155),
.B(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

AO21x2_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_90),
.B(n_80),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_156),
.B1(n_146),
.B2(n_153),
.Y(n_166)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_0),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_91),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_97),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_27),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_103),
.A2(n_86),
.B1(n_80),
.B2(n_66),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_106),
.A2(n_76),
.B(n_75),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_73),
.B(n_34),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_116),
.B(n_123),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_108),
.B1(n_105),
.B2(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_166),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_110),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_163),
.B(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_108),
.B1(n_122),
.B2(n_68),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_176),
.B1(n_178),
.B2(n_139),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_180),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_78),
.B1(n_116),
.B2(n_111),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_111),
.B(n_1),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_2),
.B(n_3),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_34),
.B1(n_18),
.B2(n_2),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_18),
.Y(n_180)
);

INVx6_ASAP7_75t_SL g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_135),
.B(n_18),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_140),
.B1(n_145),
.B2(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_148),
.B(n_1),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_188),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_132),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_196),
.C(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_186),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_150),
.B1(n_140),
.B2(n_159),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_200),
.B(n_177),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_209),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_3),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_16),
.C(n_5),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_15),
.C(n_5),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_4),
.C(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_199),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_162),
.B(n_4),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_214),
.A2(n_160),
.B1(n_185),
.B2(n_180),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_222),
.B1(n_225),
.B2(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_226),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_174),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_205),
.Y(n_250)
);

NAND2x1_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_162),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_183),
.B(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_230),
.B(n_232),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_169),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_198),
.B1(n_201),
.B2(n_204),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_219),
.B1(n_220),
.B2(n_229),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_191),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_241),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_196),
.C(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_246),
.C(n_247),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_217),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_179),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_179),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_209),
.C(n_226),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_192),
.C(n_172),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_228),
.B(n_251),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_221),
.A2(n_161),
.B1(n_167),
.B2(n_178),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_214),
.C(n_215),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_261),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_233),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_257),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_221),
.B(n_172),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_247),
.B(n_203),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_232),
.B(n_234),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_231),
.B(n_206),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_249),
.B(n_244),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_165),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_216),
.C(n_168),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_241),
.C(n_242),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_264),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_274),
.B1(n_257),
.B2(n_10),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_270),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_240),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_272),
.Y(n_277)
);

OAI322xp33_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_250),
.A3(n_237),
.B1(n_183),
.B2(n_230),
.C1(n_176),
.C2(n_181),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_6),
.C(n_8),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_263),
.C(n_254),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_6),
.B(n_9),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_281),
.A3(n_282),
.B1(n_9),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_262),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_267),
.B1(n_259),
.B2(n_11),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_267),
.B(n_259),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_277),
.B(n_12),
.Y(n_289)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_286),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_12),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_14),
.C(n_287),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_292),
.A2(n_287),
.B(n_285),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_291),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_293),
.Y(n_298)
);


endmodule