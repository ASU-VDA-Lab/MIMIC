module fake_jpeg_14885_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_50),
.Y(n_64)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_1),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_51),
.Y(n_58)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_41),
.B1(n_44),
.B2(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_2),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_38),
.B1(n_42),
.B2(n_40),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_4),
.Y(n_71)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_78),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_61),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_16),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_37),
.B1(n_18),
.B2(n_7),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_11),
.C(n_12),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_15),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.C(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_79),
.B1(n_76),
.B2(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_98),
.A3(n_91),
.B1(n_92),
.B2(n_34),
.C1(n_35),
.C2(n_31),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_32),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_92),
.B1(n_99),
.B2(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_99),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_96),
.B(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_84),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_97),
.Y(n_109)
);


endmodule