module real_jpeg_25531_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx6_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_0),
.Y(n_118)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_0),
.B(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_28),
.B1(n_33),
.B2(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_28),
.B1(n_33),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_71),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_10),
.A2(n_28),
.B1(n_63),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_12),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_93),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_93),
.Y(n_154)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_14),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_16),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_16),
.B(n_73),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_16),
.B(n_56),
.C(n_58),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_105),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_16),
.B(n_67),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_16),
.A2(n_55),
.B1(n_56),
.B2(n_105),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_16),
.B(n_39),
.C(n_89),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_16),
.A2(n_38),
.B(n_198),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_95),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_23),
.B(n_52),
.C(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_24),
.B(n_36),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.A3(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_26),
.B(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_43),
.B1(n_46),
.B2(n_49),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_37),
.A2(n_209),
.B1(n_211),
.B2(n_213),
.Y(n_208)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_38),
.A2(n_47),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_38),
.A2(n_83),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_38),
.A2(n_44),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_38),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_38),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_39),
.A2(n_40),
.B1(n_89),
.B2(n_90),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_40),
.B(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_42),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_48),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_68),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_64),
.Y(n_52)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_53),
.A2(n_64),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_54),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_54),
.A2(n_135),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_56),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_56),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_67),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_102),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B(n_74),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_104),
.B(n_107),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_80),
.B(n_95),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_86),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_86),
.A2(n_186),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_87),
.A2(n_122),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_92),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_91),
.A2(n_98),
.B(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_91),
.B(n_105),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_103),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_105),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_125),
.B2(n_126),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_243),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_156),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_142),
.B(n_156),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_148),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_143),
.A2(n_144),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_147),
.B(n_148),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_237),
.B(n_242),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_187),
.B(n_236),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_176),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_176),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_169),
.C(n_173),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_169),
.A2(n_173),
.B1(n_174),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_183),
.C(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_230),
.B(n_235),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_206),
.B(n_229),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_200),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_216),
.B(n_228),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_214),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_212),
.B(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_221),
.B(n_227),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);


endmodule