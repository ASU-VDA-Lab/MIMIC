module fake_jpeg_6264_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_9),
.B(n_4),
.Y(n_10)
);

BUFx4f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx9p33_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_37),
.Y(n_48)
);

A2O1A1O1Ixp25_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_14),
.B(n_16),
.C(n_5),
.D(n_2),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_7),
.B1(n_8),
.B2(n_4),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_20),
.B(n_5),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_28),
.B(n_23),
.C(n_16),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_43),
.B(n_34),
.C(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_37),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_39),
.B1(n_34),
.B2(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_56),
.B(n_44),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_30),
.C(n_31),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_46),
.C(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_43),
.C(n_42),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_42),
.C(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_51),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_64),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.A3(n_65),
.B1(n_64),
.B2(n_50),
.C1(n_33),
.C2(n_38),
.Y(n_70)
);

OAI21x1_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_62),
.B(n_44),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_50),
.Y(n_71)
);


endmodule