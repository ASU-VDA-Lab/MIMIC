module fake_netlist_6_3718_n_308 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_51, n_44, n_308);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_51;
input n_44;

output n_308;

wire n_52;
wire n_91;
wire n_256;
wire n_209;
wire n_63;
wire n_223;
wire n_278;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_68;
wire n_304;
wire n_212;
wire n_144;
wire n_125;
wire n_168;
wire n_297;
wire n_77;
wire n_106;
wire n_160;
wire n_131;
wire n_188;
wire n_186;
wire n_245;
wire n_78;
wire n_84;
wire n_142;
wire n_143;
wire n_180;
wire n_62;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_214;
wire n_67;
wire n_246;
wire n_289;
wire n_59;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_108;
wire n_280;
wire n_287;
wire n_65;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_71;
wire n_74;
wire n_229;
wire n_305;
wire n_72;
wire n_173;
wire n_250;
wire n_111;
wire n_183;
wire n_79;
wire n_56;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_73;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_70;
wire n_234;
wire n_82;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_58;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_80;
wire n_196;
wire n_107;
wire n_89;
wire n_103;
wire n_272;
wire n_185;
wire n_69;
wire n_293;
wire n_53;
wire n_232;
wire n_163;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_265;
wire n_260;
wire n_279;
wire n_252;
wire n_228;
wire n_166;
wire n_184;
wire n_216;
wire n_83;
wire n_152;
wire n_92;
wire n_105;
wire n_227;
wire n_132;
wire n_102;
wire n_204;
wire n_261;
wire n_66;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_150;
wire n_264;
wire n_263;
wire n_61;
wire n_237;
wire n_244;
wire n_76;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_231;
wire n_240;
wire n_139;
wire n_134;
wire n_273;
wire n_95;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_88;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_149;
wire n_90;
wire n_54;
wire n_87;
wire n_195;
wire n_285;
wire n_85;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_75;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_110;
wire n_81;
wire n_55;
wire n_267;
wire n_64;
wire n_288;
wire n_135;
wire n_165;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_60;
wire n_170;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_29),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVxp33_ASAP7_75t_SL g67 ( 
.A(n_6),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_15),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_0),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_1),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_5),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_7),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_SL g110 ( 
.A(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_58),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_83),
.Y(n_121)
);

OAI221xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_82),
.B1(n_60),
.B2(n_80),
.C(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_81),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_69),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_72),
.B1(n_68),
.B2(n_9),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_9),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_10),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_12),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_16),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_17),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_19),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_87),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_103),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_103),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_84),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_98),
.B1(n_102),
.B2(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_89),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g148 ( 
.A(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_86),
.B1(n_100),
.B2(n_92),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_150),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_141),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_115),
.B(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_141),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_150),
.B1(n_134),
.B2(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_113),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_114),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_142),
.Y(n_163)
);

O2A1O1Ixp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_123),
.B(n_130),
.C(n_121),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_122),
.B1(n_144),
.B2(n_145),
.C(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_127),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_132),
.B1(n_110),
.B2(n_131),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_133),
.B(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_21),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_22),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_23),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_110),
.C(n_25),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_154),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_24),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_26),
.B(n_28),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_30),
.B(n_32),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_33),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_34),
.B(n_35),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_161),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_162),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_191),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_159),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_155),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_155),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_157),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_161),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_205),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_165),
.B1(n_161),
.B2(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_188),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_161),
.B1(n_160),
.B2(n_188),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_157),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_193),
.B1(n_180),
.B2(n_176),
.Y(n_226)
);

INVx5_ASAP7_75t_SL g227 ( 
.A(n_208),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_195),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_203),
.C(n_174),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_210),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_206),
.Y(n_237)
);

AOI221xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_200),
.B1(n_228),
.B2(n_223),
.C(n_169),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_216),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_220),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_174),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_227),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_197),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_221),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_248),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_251),
.C(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_257),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_256),
.B(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_268),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_269),
.C(n_270),
.Y(n_279)
);

NOR2x1p5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_266),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_276),
.B1(n_275),
.B2(n_263),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_265),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_260),
.Y(n_283)
);

AO22x2_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_279),
.B1(n_283),
.B2(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

NAND5xp2_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_254),
.C(n_247),
.D(n_170),
.E(n_172),
.Y(n_289)
);

OAI322xp33_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_254),
.A3(n_247),
.B1(n_179),
.B2(n_181),
.C1(n_208),
.C2(n_186),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_221),
.B1(n_187),
.B2(n_192),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_183),
.B(n_192),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_192),
.Y(n_293)
);

OAI221xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_288),
.B1(n_173),
.B2(n_192),
.C(n_199),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_36),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

NAND4xp25_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_186),
.C(n_221),
.D(n_39),
.Y(n_298)
);

AOI32xp33_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_213),
.A3(n_212),
.B1(n_185),
.B2(n_184),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_185),
.C(n_176),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_184),
.B(n_212),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_40),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_302),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

AOI221xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_304),
.B1(n_307),
.B2(n_305),
.C(n_299),
.Y(n_308)
);


endmodule