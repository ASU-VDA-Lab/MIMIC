module fake_jpeg_32128_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_1),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_60),
.Y(n_67)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_52),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_86),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_50),
.C(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_5),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_64),
.B(n_62),
.C(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_55),
.B1(n_21),
.B2(n_22),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_3),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_23),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_106),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_20),
.B1(n_41),
.B2(n_39),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_18),
.B(n_38),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_103),
.B(n_28),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_17),
.B(n_37),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_6),
.B(n_7),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_13),
.C(n_14),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_16),
.B1(n_27),
.B2(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_117),
.B1(n_98),
.B2(n_96),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_116),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_32),
.C(n_34),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_35),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_123),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_118),
.C(n_117),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B1(n_123),
.B2(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_110),
.B1(n_93),
.B2(n_107),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_36),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_42),
.C(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_101),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule