module fake_jpeg_10847_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2x1p5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_20),
.B1(n_10),
.B2(n_16),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_42),
.B1(n_23),
.B2(n_26),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_19),
.B(n_21),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g38 ( 
.A(n_22),
.B(n_19),
.CON(n_38),
.SN(n_38)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_10),
.B1(n_20),
.B2(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_53),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_51),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_27),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_15),
.B1(n_2),
.B2(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_57),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_36),
.B(n_34),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_63),
.C(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_69),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_55),
.B(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_37),
.B1(n_40),
.B2(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_73),
.B1(n_59),
.B2(n_66),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_37),
.C(n_40),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_41),
.B1(n_45),
.B2(n_9),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_41),
.C(n_7),
.Y(n_74)
);

XOR2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_72),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_80),
.Y(n_84)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_65),
.C(n_61),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_79),
.C(n_76),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g86 ( 
.A(n_84),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_88),
.C(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_8),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_85),
.C(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_78),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_89),
.Y(n_93)
);


endmodule