module fake_jpeg_4946_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_30),
.Y(n_61)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_29),
.C(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_41),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_26),
.B(n_39),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_52),
.B(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_57),
.B1(n_66),
.B2(n_62),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_41),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_23),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_20),
.B(n_19),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_23),
.C(n_16),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_67),
.B1(n_44),
.B2(n_58),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_20),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_70),
.B1(n_82),
.B2(n_71),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_112),
.B(n_24),
.Y(n_130)
);

AO21x2_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_46),
.B(n_59),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_79),
.B(n_59),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_81),
.B1(n_78),
.B2(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_100),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_34),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_23),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_34),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_107),
.CI(n_20),
.CON(n_135),
.SN(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_20),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_51),
.B1(n_47),
.B2(n_46),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_115),
.B1(n_133),
.B2(n_138),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_85),
.B1(n_71),
.B2(n_43),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_119),
.B1(n_125),
.B2(n_126),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_107),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_112),
.B(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_73),
.B1(n_88),
.B2(n_89),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_79),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_101),
.C(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_102),
.Y(n_143)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_73),
.B1(n_89),
.B2(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_137),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_91),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_96),
.B1(n_100),
.B2(n_92),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_147),
.B1(n_150),
.B2(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_96),
.B1(n_110),
.B2(n_97),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_102),
.B(n_109),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_96),
.B1(n_102),
.B2(n_111),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_124),
.C(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_96),
.B(n_93),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_17),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_103),
.B1(n_86),
.B2(n_76),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_127),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_118),
.B1(n_117),
.B2(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_108),
.B1(n_103),
.B2(n_76),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_118),
.A2(n_76),
.B1(n_104),
.B2(n_33),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_173),
.B1(n_189),
.B2(n_150),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_177),
.C(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_117),
.B1(n_119),
.B2(n_135),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_179),
.B1(n_32),
.B2(n_9),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_138),
.B1(n_136),
.B2(n_131),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_116),
.B1(n_47),
.B2(n_19),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_182),
.B1(n_165),
.B2(n_161),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_121),
.C(n_24),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_178),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_33),
.B1(n_20),
.B2(n_30),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_142),
.C(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_147),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_32),
.C(n_28),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_158),
.C(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_30),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_146),
.A2(n_21),
.B1(n_32),
.B2(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_197),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_201),
.B(n_206),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_163),
.B(n_155),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_200),
.B(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_151),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_144),
.B(n_143),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_177),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_209),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_139),
.C(n_157),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_208),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_157),
.B1(n_21),
.B2(n_28),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_32),
.C(n_2),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_32),
.B1(n_2),
.B2(n_1),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_210),
.A2(n_182),
.B1(n_176),
.B2(n_174),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_219),
.C(n_196),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_221),
.B1(n_226),
.B2(n_198),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_218),
.B(n_200),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_175),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_166),
.B1(n_171),
.B2(n_169),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_170),
.B1(n_173),
.B2(n_1),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_228),
.A2(n_229),
.B(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_219),
.C(n_192),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_238),
.C(n_213),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_240),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_209),
.B1(n_210),
.B2(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_2),
.C(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_222),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

NAND5xp2_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_9),
.C(n_3),
.D(n_4),
.E(n_6),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_239),
.A2(n_216),
.B1(n_218),
.B2(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_2),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_250),
.C(n_251),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_236),
.C(n_238),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_220),
.C(n_214),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_234),
.B1(n_230),
.B2(n_8),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_7),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_7),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_8),
.C(n_10),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_8),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_245),
.Y(n_260)
);

AOI31xp33_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_254),
.A3(n_241),
.B(n_257),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_246),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_243),
.B1(n_246),
.B2(n_12),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_264),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_271),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_262),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_11),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_13),
.B(n_14),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_11),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_275),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_277),
.B1(n_14),
.B2(n_15),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_13),
.C(n_15),
.Y(n_281)
);


endmodule