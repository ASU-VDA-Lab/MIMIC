module fake_netlist_6_2339_n_806 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_806);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_806;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_772;
wire n_656;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_102),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_45),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_90),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_18),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_23),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_80),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_79),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_38),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_31),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_95),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_129),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_94),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_18),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_17),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_60),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_17),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_14),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_136),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_53),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_75),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_29),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_47),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_52),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_0),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_12),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_40),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_86),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_103),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_26),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_0),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_1),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_154),
.B(n_27),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_157),
.B(n_1),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_2),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_2),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_3),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_4),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_28),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_162),
.B(n_30),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_163),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_4),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_164),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_169),
.B(n_171),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_173),
.B(n_5),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_175),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_158),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_158),
.B(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_176),
.B(n_6),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_219),
.B1(n_191),
.B2(n_216),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_159),
.B1(n_172),
.B2(n_177),
.Y(n_263)
);

OR2x6_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_195),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_201),
.B1(n_212),
.B2(n_205),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_215),
.A2(n_213),
.B1(n_212),
.B2(n_205),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_217),
.A2(n_160),
.B1(n_184),
.B2(n_202),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_246),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_184),
.B1(n_203),
.B2(n_198),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_204),
.B1(n_194),
.B2(n_192),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_259),
.B1(n_251),
.B2(n_255),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_SL g273 ( 
.A(n_232),
.B(n_178),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_185),
.B1(n_181),
.B2(n_180),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_216),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_188),
.B1(n_8),
.B2(n_9),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_33),
.Y(n_279)
);

OR2x6_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_11),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_216),
.B(n_245),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

OR2x6_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_19),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_222),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_R g293 ( 
.A1(n_238),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_293)
);

AO22x2_ASAP7_75t_L g294 ( 
.A1(n_227),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_35),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_236),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

AO22x2_ASAP7_75t_L g298 ( 
.A1(n_227),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g299 ( 
.A1(n_261),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_248),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_300)
);

OR2x6_ASAP7_75t_L g301 ( 
.A(n_231),
.B(n_56),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_260),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_233),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_230),
.B(n_61),
.Y(n_304)
);

AO22x2_ASAP7_75t_L g305 ( 
.A1(n_243),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_224),
.A2(n_249),
.B1(n_254),
.B2(n_230),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

OR2x6_ASAP7_75t_L g309 ( 
.A(n_231),
.B(n_65),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_230),
.B(n_66),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_263),
.B(n_245),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_269),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

INVx4_ASAP7_75t_SL g325 ( 
.A(n_301),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_247),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_265),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_252),
.Y(n_331)
);

INVx4_ASAP7_75t_SL g332 ( 
.A(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_266),
.B(n_247),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_252),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_264),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_271),
.B(n_243),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_270),
.B(n_252),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_272),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_245),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_312),
.B(n_247),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_267),
.B(n_252),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_273),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_252),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_275),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_274),
.B(n_233),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_286),
.B(n_243),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

XNOR2x2_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_220),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_289),
.B(n_257),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_264),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_302),
.A2(n_299),
.B(n_226),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_277),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_280),
.B(n_257),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_276),
.B(n_257),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_287),
.B(n_257),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_280),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_278),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_283),
.A2(n_226),
.B(n_223),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_306),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_263),
.B(n_67),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_306),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_283),
.B(n_257),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_365),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_68),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_229),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_229),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_373),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

OR2x6_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_229),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_331),
.B(n_229),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_234),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_352),
.B(n_234),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_234),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_343),
.B(n_226),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_316),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

INVx3_ASAP7_75t_SL g407 ( 
.A(n_317),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_234),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_346),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_360),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_318),
.B(n_234),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_319),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_221),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_361),
.B(n_221),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_321),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_223),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_376),
.B(n_69),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_335),
.B(n_378),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_321),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_338),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_362),
.B(n_223),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_325),
.B(n_70),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_329),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_347),
.B(n_223),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_351),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_223),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_323),
.B(n_71),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_321),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_359),
.B(n_218),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_338),
.B(n_218),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_369),
.B(n_218),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_325),
.B(n_218),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_325),
.B(n_218),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_332),
.B(n_355),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_366),
.B(n_72),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_314),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_332),
.B(n_73),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_332),
.B(n_367),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_74),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_323),
.B(n_356),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_368),
.A2(n_77),
.B(n_78),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_407),
.B(n_344),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_356),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_368),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_372),
.Y(n_456)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_450),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_383),
.B(n_358),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_333),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_377),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_403),
.B(n_349),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_391),
.B(n_370),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_391),
.B(n_370),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_426),
.B(n_353),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_393),
.A2(n_81),
.B(n_82),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_389),
.B(n_83),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_327),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_327),
.Y(n_476)
);

NAND2x1_ASAP7_75t_SL g477 ( 
.A(n_447),
.B(n_336),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

OR2x6_ASAP7_75t_SL g479 ( 
.A(n_442),
.B(n_363),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_384),
.B(n_84),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

BUFx4f_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_403),
.B(n_85),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_87),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_414),
.Y(n_489)
);

AND2x2_ASAP7_75t_SL g490 ( 
.A(n_448),
.B(n_401),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_408),
.B(n_392),
.Y(n_492)
);

BUFx6f_ASAP7_75t_SL g493 ( 
.A(n_420),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_408),
.B(n_88),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_393),
.A2(n_152),
.B(n_91),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_449),
.B(n_89),
.Y(n_496)
);

BUFx2_ASAP7_75t_SL g497 ( 
.A(n_447),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_384),
.B(n_92),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_421),
.B(n_93),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_392),
.B(n_96),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_398),
.B(n_97),
.Y(n_502)
);

OR2x6_ASAP7_75t_L g503 ( 
.A(n_384),
.B(n_99),
.Y(n_503)
);

OR2x6_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_100),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_101),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_388),
.B(n_104),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_381),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_474),
.Y(n_509)
);

INVx6_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_455),
.A2(n_433),
.B1(n_387),
.B2(n_424),
.Y(n_512)
);

CKINVDCx8_ASAP7_75t_R g513 ( 
.A(n_470),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_467),
.Y(n_514)
);

BUFx12f_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_480),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_480),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_478),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_454),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_486),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_458),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_492),
.A2(n_451),
.B1(n_387),
.B2(n_416),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_488),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

BUFx2_ASAP7_75t_SL g527 ( 
.A(n_491),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_484),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_489),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_483),
.B(n_389),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_484),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_483),
.B(n_389),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

BUFx12f_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

BUFx2_ASAP7_75t_SL g536 ( 
.A(n_491),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_415),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_457),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_457),
.B(n_387),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_508),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

INVx8_ASAP7_75t_L g543 ( 
.A(n_493),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_466),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_456),
.B(n_431),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_460),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_487),
.Y(n_549)
);

BUFx2_ASAP7_75t_SL g550 ( 
.A(n_493),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_487),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_485),
.A2(n_451),
.B1(n_416),
.B2(n_415),
.Y(n_553)
);

BUFx12f_ASAP7_75t_L g554 ( 
.A(n_473),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

BUFx8_ASAP7_75t_L g556 ( 
.A(n_523),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_516),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_537),
.A2(n_462),
.B1(n_486),
.B2(n_496),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_510),
.A2(n_452),
.B1(n_463),
.B2(n_461),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_528),
.Y(n_560)
);

BUFx2_ASAP7_75t_SL g561 ( 
.A(n_516),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

OAI22x1_ASAP7_75t_L g563 ( 
.A1(n_512),
.A2(n_475),
.B1(n_546),
.B2(n_461),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_453),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_463),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_453),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_518),
.B(n_468),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_552),
.B(n_506),
.Y(n_570)
);

INVx6_ASAP7_75t_L g571 ( 
.A(n_543),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_510),
.A2(n_473),
.B1(n_476),
.B2(n_470),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_518),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_553),
.A2(n_462),
.B1(n_496),
.B2(n_504),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_524),
.A2(n_464),
.B1(n_493),
.B2(n_497),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_520),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_553),
.A2(n_524),
.B1(n_504),
.B2(n_490),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_529),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_520),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_543),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_517),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_526),
.Y(n_586)
);

CKINVDCx11_ASAP7_75t_R g587 ( 
.A(n_523),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_522),
.A2(n_504),
.B1(n_490),
.B2(n_503),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_522),
.A2(n_504),
.B1(n_481),
.B2(n_503),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_534),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_539),
.B(n_468),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_552),
.B(n_507),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_539),
.B(n_469),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_522),
.A2(n_481),
.B1(n_503),
.B2(n_482),
.Y(n_596)
);

CKINVDCx11_ASAP7_75t_R g597 ( 
.A(n_535),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_578),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_575),
.A2(n_539),
.B1(n_479),
.B2(n_473),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_565),
.B(n_476),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_555),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_578),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_582),
.Y(n_603)
);

CKINVDCx14_ASAP7_75t_R g604 ( 
.A(n_587),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_562),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_564),
.A2(n_479),
.B1(n_482),
.B2(n_539),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_591),
.A2(n_513),
.B1(n_510),
.B2(n_503),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_566),
.B(n_469),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_563),
.A2(n_476),
.B1(n_470),
.B2(n_554),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_569),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_567),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_579),
.A2(n_470),
.B1(n_388),
.B2(n_417),
.Y(n_612)
);

NOR2x1_ASAP7_75t_R g613 ( 
.A(n_587),
.B(n_535),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_579),
.A2(n_470),
.B1(n_417),
.B2(n_388),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_577),
.A2(n_509),
.B1(n_515),
.B2(n_536),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_575),
.A2(n_513),
.B1(n_527),
.B2(n_507),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_594),
.A2(n_509),
.B1(n_515),
.B2(n_481),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_592),
.B(n_399),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_559),
.A2(n_417),
.B1(n_481),
.B2(n_505),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_574),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_399),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_592),
.B(n_534),
.Y(n_622)
);

BUFx12f_ASAP7_75t_L g623 ( 
.A(n_597),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_584),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_580),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_586),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_501),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_549),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_572),
.A2(n_420),
.B1(n_507),
.B2(n_500),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_558),
.A2(n_552),
.B1(n_410),
.B2(n_389),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_560),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_558),
.A2(n_420),
.B1(n_500),
.B2(n_406),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_589),
.A2(n_410),
.B1(n_404),
.B2(n_533),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_589),
.A2(n_410),
.B1(n_404),
.B2(n_533),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_581),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_588),
.A2(n_405),
.B1(n_406),
.B2(n_550),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_588),
.A2(n_596),
.B1(n_405),
.B2(n_446),
.Y(n_637)
);

OAI21xp33_ASAP7_75t_L g638 ( 
.A1(n_596),
.A2(n_477),
.B(n_382),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_561),
.B(n_557),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_571),
.A2(n_410),
.B1(n_404),
.B2(n_541),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_570),
.B(n_549),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_571),
.A2(n_472),
.B1(n_502),
.B2(n_494),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_576),
.A2(n_498),
.B1(n_502),
.B2(n_499),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_571),
.A2(n_404),
.B1(n_410),
.B2(n_541),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_568),
.Y(n_645)
);

CKINVDCx11_ASAP7_75t_R g646 ( 
.A(n_597),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_570),
.B(n_551),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_629),
.A2(n_573),
.B1(n_557),
.B2(n_576),
.Y(n_648)
);

OAI222xp33_ASAP7_75t_L g649 ( 
.A1(n_599),
.A2(n_472),
.B1(n_531),
.B2(n_427),
.C1(n_397),
.C2(n_400),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_603),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_606),
.A2(n_573),
.B1(n_542),
.B2(n_595),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_638),
.A2(n_542),
.B1(n_400),
.B2(n_395),
.Y(n_652)
);

AOI222xp33_ASAP7_75t_L g653 ( 
.A1(n_600),
.A2(n_556),
.B1(n_427),
.B2(n_422),
.C1(n_395),
.C2(n_396),
.Y(n_653)
);

AOI222xp33_ASAP7_75t_L g654 ( 
.A1(n_632),
.A2(n_556),
.B1(n_396),
.B2(n_398),
.C1(n_531),
.C2(n_413),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_619),
.A2(n_595),
.B1(n_583),
.B2(n_542),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_612),
.A2(n_595),
.B1(n_583),
.B2(n_542),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_583),
.Y(n_657)
);

OAI222xp33_ASAP7_75t_L g658 ( 
.A1(n_615),
.A2(n_397),
.B1(n_560),
.B2(n_438),
.C1(n_437),
.C2(n_444),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_614),
.A2(n_609),
.B1(n_636),
.B2(n_617),
.Y(n_659)
);

AOI222xp33_ASAP7_75t_L g660 ( 
.A1(n_616),
.A2(n_413),
.B1(n_419),
.B2(n_441),
.C1(n_431),
.C2(n_444),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_637),
.A2(n_610),
.B1(n_643),
.B2(n_639),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_618),
.A2(n_444),
.B1(n_538),
.B2(n_410),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_618),
.A2(n_538),
.B1(n_404),
.B2(n_541),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_622),
.B(n_568),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_607),
.A2(n_538),
.B1(n_441),
.B2(n_439),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_621),
.A2(n_538),
.B1(n_404),
.B2(n_394),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_642),
.A2(n_402),
.B(n_438),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_627),
.A2(n_397),
.B1(n_528),
.B2(n_530),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_622),
.B(n_551),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_621),
.A2(n_394),
.B1(n_495),
.B2(n_471),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_604),
.A2(n_495),
.B1(n_471),
.B2(n_397),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_601),
.B(n_585),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_605),
.A2(n_397),
.B1(n_532),
.B2(n_530),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_611),
.B(n_585),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_620),
.A2(n_532),
.B1(n_530),
.B2(n_528),
.Y(n_675)
);

OAI222xp33_ASAP7_75t_L g676 ( 
.A1(n_604),
.A2(n_437),
.B1(n_394),
.B2(n_402),
.C1(n_435),
.C2(n_419),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_SL g677 ( 
.A(n_625),
.B(n_432),
.C(n_436),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_623),
.A2(n_435),
.B1(n_386),
.B2(n_428),
.Y(n_678)
);

OAI222xp33_ASAP7_75t_L g679 ( 
.A1(n_630),
.A2(n_435),
.B1(n_521),
.B2(n_519),
.C1(n_511),
.C2(n_386),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_635),
.B(n_585),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_633),
.A2(n_528),
.B1(n_532),
.B2(n_530),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_623),
.A2(n_435),
.B1(n_428),
.B2(n_429),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_646),
.A2(n_428),
.B1(n_429),
.B2(n_532),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_635),
.B(n_585),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_646),
.A2(n_603),
.B1(n_624),
.B2(n_626),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_650),
.B(n_626),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_659),
.A2(n_634),
.B1(n_647),
.B2(n_641),
.Y(n_687)
);

NOR2x1_ASAP7_75t_SL g688 ( 
.A(n_677),
.B(n_644),
.Y(n_688)
);

OAI221xp5_ASAP7_75t_SL g689 ( 
.A1(n_685),
.A2(n_613),
.B1(n_624),
.B2(n_641),
.C(n_647),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_664),
.B(n_602),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_661),
.B(n_631),
.C(n_640),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_685),
.B(n_598),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_654),
.A2(n_631),
.B1(n_645),
.B2(n_628),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_657),
.B(n_631),
.Y(n_694)
);

NAND4xp25_ASAP7_75t_L g695 ( 
.A(n_653),
.B(n_628),
.C(n_602),
.D(n_598),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_658),
.B(n_648),
.C(n_651),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_568),
.Y(n_697)
);

OA211x2_ASAP7_75t_L g698 ( 
.A1(n_652),
.A2(n_667),
.B(n_683),
.C(n_670),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_672),
.B(n_568),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_665),
.A2(n_521),
.B1(n_519),
.B2(n_511),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_674),
.B(n_106),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_680),
.B(n_107),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_684),
.B(n_671),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_676),
.B(n_521),
.C(n_519),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_660),
.B(n_109),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_655),
.A2(n_429),
.B1(n_432),
.B2(n_511),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_SL g707 ( 
.A1(n_683),
.A2(n_436),
.B1(n_430),
.B2(n_425),
.C(n_440),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_668),
.B(n_434),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_663),
.B(n_434),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_656),
.B(n_434),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_662),
.B(n_517),
.Y(n_711)
);

OAI221xp5_ASAP7_75t_SL g712 ( 
.A1(n_678),
.A2(n_430),
.B1(n_425),
.B2(n_440),
.C(n_117),
.Y(n_712)
);

NAND4xp25_ASAP7_75t_SL g713 ( 
.A(n_682),
.B(n_112),
.C(n_113),
.D(n_115),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_703),
.B(n_675),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_686),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_686),
.Y(n_716)
);

XNOR2xp5_ASAP7_75t_L g717 ( 
.A(n_690),
.B(n_682),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_703),
.B(n_673),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_690),
.B(n_666),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_689),
.B(n_649),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_692),
.B(n_681),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_694),
.B(n_678),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_699),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_118),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_696),
.B(n_517),
.C(n_418),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_715),
.B(n_688),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_714),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_716),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

NAND4xp75_ASAP7_75t_L g731 ( 
.A(n_720),
.B(n_698),
.C(n_705),
.D(n_702),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_714),
.Y(n_732)
);

NAND4xp75_ASAP7_75t_L g733 ( 
.A(n_720),
.B(n_698),
.C(n_705),
.D(n_702),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_718),
.B(n_697),
.Y(n_734)
);

OAI22x1_ASAP7_75t_L g735 ( 
.A1(n_732),
.A2(n_717),
.B1(n_718),
.B2(n_725),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_730),
.B(n_719),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_727),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_726),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_732),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_730),
.Y(n_740)
);

AO22x1_ASAP7_75t_L g741 ( 
.A1(n_740),
.A2(n_726),
.B1(n_728),
.B2(n_727),
.Y(n_741)
);

XOR2x2_ASAP7_75t_L g742 ( 
.A(n_736),
.B(n_733),
.Y(n_742)
);

AOI22x1_ASAP7_75t_L g743 ( 
.A1(n_735),
.A2(n_731),
.B1(n_729),
.B2(n_724),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_740),
.B(n_734),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_739),
.Y(n_745)
);

OAI322xp33_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_744),
.A3(n_738),
.B1(n_745),
.B2(n_737),
.C1(n_734),
.C2(n_742),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_741),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_745),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_749),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_746),
.B(n_738),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_750),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_L g753 ( 
.A1(n_751),
.A2(n_747),
.B1(n_748),
.B2(n_712),
.C(n_695),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_751),
.A2(n_724),
.B(n_707),
.C(n_691),
.Y(n_754)
);

OA22x2_ASAP7_75t_L g755 ( 
.A1(n_752),
.A2(n_722),
.B1(n_719),
.B2(n_706),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_754),
.B(n_701),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_753),
.A2(n_713),
.B1(n_693),
.B2(n_704),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_752),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_752),
.Y(n_759)
);

NOR4xp25_ASAP7_75t_L g760 ( 
.A(n_753),
.B(n_708),
.C(n_710),
.D(n_709),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_758),
.Y(n_761)
);

AO22x2_ASAP7_75t_L g762 ( 
.A1(n_759),
.A2(n_688),
.B1(n_711),
.B2(n_700),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_755),
.B(n_423),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_757),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_756),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_760),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_758),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_765),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_761),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_767),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_764),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_763),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_766),
.B(n_119),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_762),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_769),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_769),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_768),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_773),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_771),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_774),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_770),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_772),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_777),
.A2(n_762),
.B1(n_418),
.B2(n_423),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_778),
.A2(n_418),
.B1(n_423),
.B2(n_412),
.Y(n_784)
);

OAI22x1_ASAP7_75t_L g785 ( 
.A1(n_776),
.A2(n_418),
.B1(n_123),
.B2(n_124),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_776),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_775),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_780),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_SL g789 ( 
.A1(n_779),
.A2(n_423),
.B1(n_412),
.B2(n_126),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_782),
.A2(n_423),
.B1(n_412),
.B2(n_679),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_781),
.A2(n_423),
.B1(n_412),
.B2(n_128),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_786),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_787),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_788),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_784),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_785),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_789),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_790),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_797),
.A2(n_783),
.B1(n_791),
.B2(n_412),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_792),
.A2(n_412),
.B1(n_125),
.B2(n_130),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_796),
.A2(n_121),
.B1(n_131),
.B2(n_133),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_801),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_802),
.A2(n_794),
.B1(n_793),
.B2(n_798),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_803),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_804),
.A2(n_794),
.B1(n_799),
.B2(n_795),
.Y(n_805)
);

AOI211xp5_ASAP7_75t_L g806 ( 
.A1(n_805),
.A2(n_800),
.B(n_135),
.C(n_137),
.Y(n_806)
);


endmodule