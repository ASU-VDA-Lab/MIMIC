module fake_jpeg_2210_n_536 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_536);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_60),
.B(n_75),
.Y(n_143)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_61),
.Y(n_209)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_12),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_22),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_69),
.A2(n_102),
.B1(n_75),
.B2(n_109),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_12),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_76),
.B(n_102),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_81),
.Y(n_181)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_87),
.Y(n_151)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_90),
.Y(n_201)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_43),
.B(n_12),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_36),
.B(n_18),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_36),
.B(n_9),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_110),
.B(n_15),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_39),
.B(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_119),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_28),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_117),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_38),
.B(n_0),
.CON(n_121),
.SN(n_121)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_121),
.B(n_123),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_26),
.B(n_9),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_137),
.A2(n_162),
.B1(n_202),
.B2(n_203),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_82),
.A2(n_48),
.B1(n_52),
.B2(n_51),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_138),
.A2(n_142),
.B1(n_158),
.B2(n_160),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_42),
.B1(n_39),
.B2(n_46),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_149),
.B(n_200),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_48),
.B1(n_51),
.B2(n_26),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_88),
.A2(n_51),
.B1(n_40),
.B2(n_26),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_69),
.A2(n_51),
.B1(n_40),
.B2(n_26),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_123),
.B(n_45),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_77),
.B(n_45),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_193),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_92),
.A2(n_40),
.B1(n_119),
.B2(n_116),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_206),
.B1(n_6),
.B2(n_16),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_79),
.B(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_117),
.B(n_40),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_13),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_203),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_83),
.B(n_13),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_85),
.A2(n_54),
.B1(n_38),
.B2(n_3),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_98),
.A2(n_38),
.B1(n_1),
.B2(n_0),
.Y(n_207)
);

AO22x1_ASAP7_75t_SL g222 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_222)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_210),
.Y(n_290)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_164),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_112),
.B1(n_8),
.B2(n_3),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_212),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_215),
.B(n_226),
.Y(n_328)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_0),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_218),
.Y(n_306)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_125),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_221),
.B(n_241),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_222),
.A2(n_134),
.B(n_181),
.Y(n_297)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_225),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_227),
.Y(n_327)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_229),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_6),
.B1(n_16),
.B2(n_3),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_231),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_124),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_234),
.Y(n_316)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_235),
.Y(n_308)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_153),
.A2(n_14),
.B1(n_16),
.B2(n_5),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_240),
.B1(n_242),
.B2(n_256),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_124),
.Y(n_238)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_157),
.A2(n_5),
.B1(n_6),
.B2(n_14),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_139),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_143),
.A2(n_5),
.B1(n_15),
.B2(n_17),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_184),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_152),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_255),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_143),
.A2(n_5),
.B1(n_15),
.B2(n_0),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_248),
.A2(n_268),
.B1(n_271),
.B2(n_274),
.Y(n_312)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_164),
.Y(n_249)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

BUFx16f_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_252),
.Y(n_303)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_1),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_184),
.A2(n_1),
.B1(n_207),
.B2(n_141),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_158),
.A2(n_206),
.B1(n_207),
.B2(n_160),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_222),
.B1(n_255),
.B2(n_259),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_159),
.A2(n_151),
.B1(n_126),
.B2(n_150),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_259),
.A2(n_254),
.B1(n_265),
.B2(n_277),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_140),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_192),
.Y(n_262)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_166),
.Y(n_263)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_155),
.B(n_165),
.C(n_170),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_218),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g267 ( 
.A(n_152),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_272),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_147),
.A2(n_156),
.B1(n_195),
.B2(n_163),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_128),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_173),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_273),
.Y(n_309)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_128),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_188),
.B(n_136),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_190),
.A2(n_196),
.B1(n_138),
.B2(n_204),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_129),
.B(n_197),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_276),
.Y(n_321)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_174),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_187),
.B(n_151),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_130),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_280),
.A2(n_247),
.B1(n_267),
.B2(n_251),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_191),
.B1(n_130),
.B2(n_132),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_284),
.A2(n_318),
.B1(n_280),
.B2(n_271),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_214),
.B(n_191),
.C(n_132),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_288),
.B(n_299),
.C(n_314),
.Y(n_344)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_250),
.A2(n_146),
.A3(n_135),
.B1(n_144),
.B2(n_127),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_291),
.B(n_311),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_134),
.B(n_181),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_296),
.A2(n_322),
.B(n_325),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_297),
.A2(n_331),
.B1(n_238),
.B2(n_269),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_305),
.Y(n_334)
);

AOI32xp33_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_242),
.A3(n_257),
.B1(n_256),
.B2(n_218),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_244),
.B(n_266),
.C(n_239),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_315),
.A2(n_225),
.B1(n_229),
.B2(n_264),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_222),
.A2(n_255),
.B1(n_219),
.B2(n_216),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_224),
.B(n_227),
.C(n_220),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_319),
.B(n_305),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_261),
.A2(n_236),
.B(n_252),
.Y(n_322)
);

XOR2x2_ASAP7_75t_L g324 ( 
.A(n_213),
.B(n_223),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_276),
.C(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_313),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_338),
.A2(n_356),
.B1(n_359),
.B2(n_368),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_339),
.A2(n_369),
.B1(n_355),
.B2(n_346),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_340),
.A2(n_343),
.B1(n_369),
.B2(n_363),
.Y(n_400)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_296),
.A2(n_230),
.B1(n_253),
.B2(n_228),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_357),
.B1(n_367),
.B2(n_372),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_283),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_346),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_288),
.B(n_243),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_233),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_349),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_232),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_350),
.Y(n_386)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_352),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_310),
.A2(n_210),
.B1(n_278),
.B2(n_263),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_353),
.A2(n_364),
.B1(n_293),
.B2(n_313),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_287),
.A2(n_252),
.B(n_249),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_354),
.A2(n_367),
.B(n_345),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_309),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_360),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_315),
.A2(n_211),
.B1(n_234),
.B2(n_314),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_282),
.A2(n_297),
.B1(n_318),
.B2(n_306),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_328),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_363),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_297),
.A2(n_332),
.B1(n_299),
.B2(n_285),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_361),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_305),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_362),
.A2(n_366),
.B(n_354),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_289),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_298),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_371),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_302),
.B(n_305),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_287),
.A2(n_300),
.B1(n_285),
.B2(n_302),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_332),
.A2(n_325),
.B1(n_312),
.B2(n_300),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_281),
.B(n_320),
.C(n_303),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_308),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_321),
.B(n_319),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_304),
.A2(n_281),
.B1(n_326),
.B2(n_289),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_371),
.A2(n_322),
.B(n_329),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_373),
.A2(n_378),
.B(n_391),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_342),
.B1(n_336),
.B2(n_364),
.Y(n_415)
);

A2O1A1O1Ixp25_ASAP7_75t_L g378 ( 
.A1(n_344),
.A2(n_327),
.B(n_286),
.C(n_292),
.D(n_290),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_357),
.A2(n_330),
.B1(n_329),
.B2(n_323),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_387),
.A2(n_400),
.B1(n_339),
.B2(n_370),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_356),
.A2(n_323),
.B1(n_327),
.B2(n_292),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_389),
.A2(n_390),
.B1(n_372),
.B2(n_335),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_338),
.B1(n_334),
.B2(n_340),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_368),
.A2(n_290),
.B1(n_293),
.B2(n_308),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_344),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_394),
.B(n_341),
.C(n_365),
.Y(n_422)
);

AO22x1_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_366),
.B1(n_334),
.B2(n_337),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_395),
.A2(n_403),
.B(n_404),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_348),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_399),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_366),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_352),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_347),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_345),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_409),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_406),
.A2(n_389),
.B1(n_387),
.B2(n_402),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_407),
.B(n_421),
.Y(n_443)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_333),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_411),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_412),
.A2(n_389),
.B1(n_377),
.B2(n_393),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_384),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_413),
.Y(n_456)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_414),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_422),
.B(n_373),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_347),
.C(n_349),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_425),
.C(n_427),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g418 ( 
.A(n_385),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_431),
.Y(n_452)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_375),
.A2(n_342),
.B1(n_350),
.B2(n_364),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_424),
.A2(n_426),
.B1(n_412),
.B2(n_391),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_351),
.C(n_350),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_375),
.A2(n_390),
.B1(n_400),
.B2(n_377),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_380),
.C(n_379),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_385),
.B(n_379),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_398),
.C(n_383),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_403),
.A2(n_404),
.B(n_399),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_432),
.B(n_394),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_380),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_373),
.A2(n_393),
.B(n_395),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_388),
.Y(n_434)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_434),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_438),
.A2(n_440),
.B1(n_447),
.B2(n_424),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_405),
.B(n_388),
.Y(n_439)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_439),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_441),
.A2(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_432),
.A2(n_394),
.B(n_402),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_449),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_426),
.A2(n_391),
.B1(n_394),
.B2(n_386),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_407),
.B(n_378),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_450),
.B(n_429),
.Y(n_459)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_420),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_378),
.B1(n_376),
.B2(n_386),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_419),
.A2(n_383),
.B1(n_397),
.B2(n_421),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_427),
.C(n_416),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_474),
.C(n_450),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_460),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_443),
.B(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_425),
.Y(n_461)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_457),
.B1(n_434),
.B2(n_444),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_473),
.Y(n_483)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_467),
.C(n_471),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_452),
.B(n_428),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_406),
.Y(n_469)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_469),
.Y(n_480)
);

AOI21xp33_ASAP7_75t_L g471 ( 
.A1(n_433),
.A2(n_420),
.B(n_417),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_454),
.A2(n_438),
.B1(n_455),
.B2(n_447),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_472),
.A2(n_441),
.B1(n_440),
.B2(n_439),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_443),
.B(n_417),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_423),
.C(n_408),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_433),
.B(n_410),
.Y(n_476)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_476),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_477),
.A2(n_470),
.B1(n_462),
.B2(n_468),
.Y(n_493)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_487),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_453),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_489),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_486),
.A2(n_472),
.B1(n_470),
.B2(n_469),
.Y(n_492)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_463),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_437),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_442),
.C(n_451),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_491),
.C(n_462),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_444),
.C(n_448),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_493),
.B1(n_486),
.B2(n_481),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_483),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_461),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_478),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_460),
.C(n_473),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_499),
.C(n_479),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_498),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_459),
.C(n_475),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_477),
.A2(n_468),
.B1(n_449),
.B2(n_422),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_422),
.Y(n_507)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_502),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_483),
.B(n_422),
.Y(n_503)
);

NOR2x1_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_480),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_500),
.Y(n_516)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_495),
.B1(n_479),
.B2(n_496),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_509),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_484),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_508),
.B(n_511),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_499),
.B(n_482),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_498),
.B(n_494),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_516),
.Y(n_524)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_510),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_513),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_506),
.A2(n_501),
.B1(n_437),
.B2(n_435),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_513),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_510),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_522),
.A2(n_525),
.B(n_526),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_523),
.A2(n_521),
.B(n_520),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_518),
.A2(n_509),
.B(n_504),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_529),
.B(n_512),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_524),
.A2(n_516),
.B(n_507),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_531),
.B(n_435),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_522),
.C(n_503),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_445),
.Y(n_533)
);

AO21x1_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_414),
.B(n_445),
.Y(n_534)
);

OAI221xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_446),
.B1(n_448),
.B2(n_422),
.C(n_397),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_446),
.Y(n_536)
);


endmodule