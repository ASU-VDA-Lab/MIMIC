module fake_aes_192_n_21 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
INVx1_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_1), .B(n_8), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_0), .B(n_5), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
AND2x6_ASAP7_75t_SL g14 ( .A(n_12), .B(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_13), .B(n_2), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
AOI211xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_10), .B(n_14), .C(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_19), .B(n_9), .Y(n_20) );
NAND3xp33_ASAP7_75t_L g21 ( .A(n_20), .B(n_6), .C(n_7), .Y(n_21) );
endmodule