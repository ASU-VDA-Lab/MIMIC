module fake_jpeg_2429_n_382 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_61),
.Y(n_118)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_9),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_26),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_63),
.B(n_83),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g155 ( 
.A(n_64),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_15),
.B(n_14),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_0),
.C(n_1),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_72),
.Y(n_166)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_11),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_82),
.B(n_84),
.Y(n_157)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_35),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx2_ASAP7_75t_SL g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_10),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_92),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_94),
.Y(n_121)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_102),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g170 ( 
.A(n_97),
.B(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_100),
.Y(n_154)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_108),
.Y(n_132)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_104),
.B(n_105),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_35),
.B(n_10),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_107),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_38),
.B(n_0),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_110),
.B1(n_48),
.B2(n_17),
.Y(n_114)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_48),
.B1(n_36),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_112),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_43),
.B1(n_41),
.B2(n_44),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_73),
.A2(n_43),
.B1(n_37),
.B2(n_33),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_19),
.B1(n_42),
.B2(n_25),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_136),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_66),
.A2(n_27),
.B1(n_44),
.B2(n_20),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_64),
.A2(n_42),
.B1(n_25),
.B2(n_22),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_56),
.A2(n_29),
.B1(n_17),
.B2(n_2),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_137),
.A2(n_148),
.B1(n_150),
.B2(n_153),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_144),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_58),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g205 ( 
.A1(n_141),
.A2(n_145),
.B1(n_152),
.B2(n_163),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_29),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_29),
.C(n_4),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_59),
.A2(n_1),
.B1(n_6),
.B2(n_65),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_64),
.A2(n_109),
.B1(n_57),
.B2(n_74),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_71),
.A2(n_106),
.B1(n_86),
.B2(n_110),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_102),
.A2(n_91),
.B1(n_89),
.B2(n_94),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_89),
.A2(n_94),
.B1(n_99),
.B2(n_86),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_156),
.A2(n_168),
.B1(n_173),
.B2(n_114),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_83),
.B(n_99),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_84),
.B(n_63),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_157),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_92),
.A2(n_93),
.B1(n_65),
.B2(n_59),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_73),
.A2(n_52),
.B1(n_53),
.B2(n_51),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_73),
.A2(n_52),
.B1(n_53),
.B2(n_51),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_92),
.A2(n_93),
.B1(n_65),
.B2(n_59),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_163),
.B1(n_112),
.B2(n_137),
.Y(n_224)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_179),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_180),
.B(n_189),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_114),
.B1(n_129),
.B2(n_131),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_181),
.A2(n_193),
.B1(n_194),
.B2(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_203),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_166),
.B1(n_119),
.B2(n_133),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_111),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_188),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_134),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_152),
.A2(n_149),
.B1(n_174),
.B2(n_117),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_118),
.B(n_135),
.CI(n_162),
.CON(n_191),
.SN(n_191)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_191),
.B(n_206),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_117),
.A2(n_147),
.B1(n_167),
.B2(n_177),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_192),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_173),
.B1(n_125),
.B2(n_126),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_163),
.A2(n_141),
.B1(n_175),
.B2(n_150),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_143),
.B1(n_141),
.B2(n_154),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_198),
.A2(n_208),
.B(n_214),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_121),
.B(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_139),
.B(n_121),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_211),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_143),
.A2(n_127),
.B1(n_165),
.B2(n_153),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_113),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

AND2x4_ASAP7_75t_SL g214 ( 
.A(n_124),
.B(n_151),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_156),
.A2(n_130),
.B1(n_124),
.B2(n_151),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_220),
.B1(n_224),
.B2(n_228),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_155),
.A2(n_171),
.B(n_138),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_218),
.C(n_215),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_164),
.Y(n_218)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_155),
.A2(n_115),
.B1(n_138),
.B2(n_159),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_132),
.A2(n_114),
.B1(n_129),
.B2(n_131),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_140),
.B(n_132),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_230),
.B1(n_214),
.B2(n_199),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_143),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_132),
.A2(n_140),
.B1(n_112),
.B2(n_148),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_186),
.Y(n_244)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_133),
.B(n_162),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_240),
.A2(n_264),
.B1(n_197),
.B2(n_196),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_244),
.B(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_187),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_205),
.B1(n_228),
.B2(n_226),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_205),
.A2(n_183),
.B1(n_210),
.B2(n_184),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_205),
.A2(n_183),
.B1(n_213),
.B2(n_201),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_178),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_265),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_209),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_231),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_214),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_202),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_242),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_204),
.B(n_229),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_261),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_217),
.B(n_232),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_258),
.B(n_235),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_239),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_277),
.Y(n_306)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_218),
.B1(n_222),
.B2(n_211),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_279),
.A2(n_294),
.B1(n_269),
.B2(n_255),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

XOR2x1_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_191),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_301),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_237),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_283),
.B(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_245),
.B(n_207),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_285),
.B(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_291),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_195),
.C(n_203),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_296),
.C(n_297),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_218),
.B1(n_221),
.B2(n_212),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_292),
.B1(n_235),
.B2(n_276),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_200),
.B1(n_191),
.B2(n_219),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_297),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_266),
.B1(n_256),
.B2(n_249),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_251),
.B(n_238),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_251),
.B(n_261),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_243),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_275),
.A2(n_234),
.B(n_249),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_317),
.B(n_285),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_R g309 ( 
.A1(n_282),
.A2(n_264),
.B(n_257),
.C(n_234),
.Y(n_309)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_295),
.A3(n_257),
.B1(n_283),
.B2(n_287),
.C(n_277),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_240),
.B1(n_254),
.B2(n_235),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_284),
.B1(n_290),
.B2(n_292),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_318),
.B1(n_288),
.B2(n_280),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_315),
.A2(n_263),
.B(n_243),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_289),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_241),
.B(n_255),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_273),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_320),
.A2(n_323),
.B1(n_333),
.B2(n_311),
.Y(n_339)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_325),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_329),
.B1(n_314),
.B2(n_318),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_279),
.B1(n_293),
.B2(n_273),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_296),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_299),
.C(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_331),
.Y(n_345)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_310),
.A3(n_309),
.B1(n_308),
.B2(n_303),
.C(n_302),
.Y(n_335)
);

O2A1O1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_281),
.B(n_278),
.C(n_298),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_330),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_312),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_247),
.B(n_271),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_332),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_295),
.B1(n_274),
.B2(n_248),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_312),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_328),
.C(n_327),
.Y(n_355)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_334),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_340),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_322),
.A2(n_304),
.B1(n_311),
.B2(n_313),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_346),
.B(n_339),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_347),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_324),
.B(n_332),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_349),
.A2(n_324),
.B(n_330),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_326),
.C(n_316),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_342),
.C(n_304),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_326),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_353),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_327),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_355),
.A2(n_356),
.B1(n_302),
.B2(n_331),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_364),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_360),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_352),
.A2(n_340),
.B1(n_341),
.B2(n_347),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_352),
.A2(n_335),
.B(n_336),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_361),
.A2(n_349),
.B(n_341),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_353),
.B(n_310),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_362),
.B(n_302),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_336),
.B(n_335),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_370),
.B(n_363),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_367),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_358),
.B(n_357),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_350),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_367),
.C(n_351),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_371),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_374),
.B(n_325),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_342),
.C(n_348),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_376),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_354),
.C(n_348),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_354),
.B(n_338),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_R g381 ( 
.A(n_380),
.B(n_379),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_344),
.Y(n_382)
);


endmodule