module fake_jpeg_19112_n_228 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_24),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_49),
.B1(n_39),
.B2(n_24),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_30),
.C(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_38),
.B(n_34),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_63),
.B(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_73),
.B1(n_58),
.B2(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_47),
.B1(n_37),
.B2(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_42),
.B1(n_32),
.B2(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_89),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_79),
.B1(n_42),
.B2(n_27),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_56),
.B1(n_44),
.B2(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_53),
.C(n_47),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_51),
.B1(n_37),
.B2(n_65),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_35),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_25),
.B(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_31),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_31),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_11),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_69),
.B(n_64),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_96),
.B(n_103),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_64),
.B(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_89),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_42),
.B1(n_37),
.B2(n_65),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_106),
.B1(n_107),
.B2(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_20),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_42),
.B1(n_60),
.B2(n_74),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_28),
.B(n_18),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_17),
.B(n_18),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_48),
.B(n_12),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_66),
.B(n_2),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_60),
.B1(n_70),
.B2(n_40),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_60),
.B1(n_40),
.B2(n_27),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_112),
.B1(n_116),
.B2(n_131),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_126),
.B1(n_128),
.B2(n_22),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_77),
.B1(n_92),
.B2(n_100),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_86),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_130),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_75),
.B1(n_90),
.B2(n_80),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_82),
.B(n_84),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_12),
.B(n_16),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_36),
.C(n_29),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_124),
.C(n_132),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_96),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_29),
.C(n_46),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_18),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_19),
.B1(n_22),
.B2(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_129),
.B1(n_17),
.B2(n_20),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_40),
.B1(n_46),
.B2(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_101),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_23),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_105),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_137),
.Y(n_167)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_135),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_106),
.B1(n_98),
.B2(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_148),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_23),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_10),
.C(n_16),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_16),
.B(n_13),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_17),
.B(n_20),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_22),
.B1(n_19),
.B2(n_12),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_29),
.C(n_22),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_23),
.C(n_15),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_132),
.B1(n_128),
.B2(n_109),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_114),
.B1(n_117),
.B2(n_116),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_124),
.B1(n_118),
.B2(n_121),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_131),
.CI(n_23),
.CON(n_162),
.SN(n_162)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_29),
.C(n_19),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_169),
.C(n_138),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_134),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

OAI321xp33_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_143),
.A3(n_149),
.B1(n_146),
.B2(n_148),
.C(n_136),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_183),
.B1(n_161),
.B2(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_180),
.B(n_23),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_144),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_182),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_158),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_155),
.B1(n_159),
.B2(n_154),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_193),
.B1(n_189),
.B2(n_187),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_160),
.B1(n_159),
.B2(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_141),
.B1(n_162),
.B2(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_150),
.B1(n_162),
.B2(n_13),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_179),
.B1(n_182),
.B2(n_181),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_175),
.B(n_180),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_196),
.B(n_203),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_201),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_13),
.B(n_10),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_1),
.B(n_2),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_15),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_1),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_194),
.B1(n_190),
.B2(n_3),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_211),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_1),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_199),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_4),
.B(n_5),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_6),
.B(n_7),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_5),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_6),
.Y(n_218)
);

OAI321xp33_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_168),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_212),
.B1(n_213),
.B2(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_220),
.C(n_8),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_8),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_9),
.Y(n_228)
);


endmodule