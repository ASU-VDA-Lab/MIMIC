module real_aes_3720_n_5 (n_4, n_0, n_3, n_2, n_1, n_5);
input n_4;
input n_0;
input n_3;
input n_2;
input n_1;
output n_5;
wire n_16;
wire n_13;
wire n_15;
wire n_7;
wire n_9;
wire n_6;
wire n_12;
wire n_8;
wire n_14;
wire n_10;
wire n_11;
NAND3xp33_ASAP7_75t_SL g6 ( .A(n_0), .B(n_7), .C(n_9), .Y(n_6) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx2_ASAP7_75t_SL g14 ( .A(n_3), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
AOI31xp33_ASAP7_75t_L g5 ( .A1(n_6), .A2(n_12), .A3(n_15), .B(n_16), .Y(n_5) );
INVx1_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
BUFx2_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_12), .B(n_15), .Y(n_16) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
endmodule