module fake_jpeg_19597_n_300 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_24),
.B1(n_28),
.B2(n_14),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_24),
.B1(n_28),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_92)
);

OR2x4_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_40),
.B(n_36),
.C(n_35),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_62),
.A2(n_65),
.B1(n_69),
.B2(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_33),
.B1(n_43),
.B2(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_43),
.B1(n_33),
.B2(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_43),
.B1(n_33),
.B2(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_30),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_78),
.B1(n_26),
.B2(n_17),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_23),
.B(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_94),
.B1(n_96),
.B2(n_102),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_28),
.B1(n_21),
.B2(n_29),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_86),
.B1(n_88),
.B2(n_100),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_35),
.C(n_36),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_84),
.Y(n_117)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_93),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_28),
.B1(n_21),
.B2(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_16),
.B1(n_34),
.B2(n_44),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_41),
.B1(n_42),
.B2(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_32),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_29),
.B1(n_17),
.B2(n_25),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_42),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_29),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_15),
.B1(n_14),
.B2(n_18),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_22),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_102),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_107),
.B(n_110),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_101),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_125),
.B1(n_80),
.B2(n_83),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_127),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_31),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_14),
.B1(n_15),
.B2(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_31),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_31),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_136),
.C(n_79),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_25),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_22),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_15),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_78),
.A3(n_64),
.B1(n_68),
.B2(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_65),
.Y(n_144)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_74),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_152),
.Y(n_172)
);

OR2x2_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_62),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_144),
.B(n_153),
.Y(n_171)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_145),
.Y(n_193)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_146),
.B(n_161),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_136),
.Y(n_168)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_90),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_157),
.B1(n_160),
.B2(n_126),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_66),
.C(n_89),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_158),
.C(n_165),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_87),
.B1(n_77),
.B2(n_84),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_100),
.B1(n_88),
.B2(n_22),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_125),
.B1(n_138),
.B2(n_121),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_61),
.B1(n_89),
.B2(n_25),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_89),
.C(n_67),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_16),
.A3(n_31),
.B1(n_13),
.B2(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_163),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_16),
.B1(n_11),
.B2(n_2),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_105),
.B(n_11),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_0),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_166),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_91),
.C(n_44),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_0),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_177),
.C(n_194),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_131),
.B(n_107),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_187),
.B1(n_108),
.B2(n_148),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_107),
.C(n_132),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_145),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_121),
.B(n_119),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_182),
.B(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_109),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_109),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_130),
.B(n_119),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_143),
.B1(n_16),
.B2(n_156),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_111),
.B1(n_123),
.B2(n_134),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_183),
.B1(n_170),
.B2(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_111),
.B1(n_135),
.B2(n_108),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_111),
.B1(n_108),
.B2(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_104),
.B(n_128),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_124),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_140),
.A2(n_128),
.B(n_129),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_104),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_194),
.C(n_168),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_176),
.C(n_167),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_173),
.B1(n_184),
.B2(n_180),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_200),
.B1(n_206),
.B2(n_212),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_158),
.B1(n_165),
.B2(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_214),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_169),
.B(n_152),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_220),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_208),
.B(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_129),
.B(n_1),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_188),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_156),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_181),
.A2(n_16),
.B1(n_44),
.B2(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_219),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_16),
.B1(n_1),
.B2(n_3),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_172),
.A3(n_195),
.B1(n_177),
.B2(n_171),
.C1(n_188),
.C2(n_190),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_198),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_216),
.B1(n_219),
.B2(n_214),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_213),
.C(n_206),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_176),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_246),
.C(n_252),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_199),
.B1(n_201),
.B2(n_197),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_244),
.B1(n_239),
.B2(n_227),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_201),
.B1(n_217),
.B2(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_213),
.C(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_250),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_210),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_253),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_209),
.C(n_202),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_220),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_225),
.B(n_239),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_267),
.B(n_269),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_264),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_227),
.B1(n_232),
.B2(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_228),
.B1(n_221),
.B2(n_230),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_221),
.B1(n_185),
.B2(n_167),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_255),
.C(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_248),
.C(n_249),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_275),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_253),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_268),
.C(n_267),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_286),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_278),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_270),
.B(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_285),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_271),
.C(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_0),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g288 ( 
.A1(n_285),
.A2(n_257),
.B(n_185),
.C(n_4),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_282),
.B1(n_3),
.B2(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_288),
.A3(n_290),
.B1(n_289),
.B2(n_7),
.C(n_3),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_5),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_296),
.B(n_6),
.C(n_9),
.D(n_10),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_298),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_5),
.Y(n_300)
);


endmodule