module fake_netlist_5_2199_n_1147 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1147);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1147;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_983;
wire n_725;
wire n_823;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_443;
wire n_293;
wire n_372;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_1048;
wire n_946;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_1032;
wire n_981;
wire n_929;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_1104;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_449;
wire n_325;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_1020;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_897;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_517;
wire n_482;
wire n_342;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_1014;
wire n_917;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_1091;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_647;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_952;
wire n_870;
wire n_809;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_985;
wire n_904;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_131),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_114),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_64),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_42),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_36),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_75),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_141),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_38),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_77),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_83),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_37),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_89),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_74),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_96),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_82),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_98),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_81),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_171),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_80),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_55),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_161),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_108),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_130),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_158),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_176),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_107),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_66),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_137),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_163),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_172),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_23),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_120),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_139),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_32),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_128),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_58),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_22),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_67),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_2),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_27),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_100),
.Y(n_264)
);

BUFx8_ASAP7_75t_SL g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_94),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_62),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_47),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_198),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_0),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_122),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_218),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_206),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_252),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_206),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_211),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_260),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_211),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_215),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_240),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_251),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_245),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_245),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_272),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_262),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_212),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_225),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_204),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_292),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_235),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_244),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_282),
.A2(n_234),
.B(n_207),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_253),
.Y(n_333)
);

OAI22x1_ASAP7_75t_SL g334 ( 
.A1(n_319),
.A2(n_212),
.B1(n_210),
.B2(n_208),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_282),
.A2(n_289),
.B(n_286),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_213),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g345 ( 
.A1(n_321),
.A2(n_225),
.B(n_216),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_295),
.B(n_214),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_301),
.A2(n_237),
.B1(n_259),
.B2(n_257),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_278),
.B(n_0),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_290),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_221),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_222),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_224),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_303),
.A2(n_266),
.B1(n_256),
.B2(n_254),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_306),
.A2(n_236),
.B1(n_247),
.B2(n_246),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_304),
.B(n_226),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_304),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_310),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_283),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_285),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_338),
.Y(n_385)
);

AO21x2_ASAP7_75t_L g386 ( 
.A1(n_345),
.A2(n_225),
.B(n_228),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_329),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_277),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

AOI21x1_ASAP7_75t_L g391 ( 
.A1(n_353),
.A2(n_225),
.B(n_229),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_355),
.A2(n_225),
.B(n_230),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_329),
.B(n_232),
.Y(n_397)
);

AO22x2_ASAP7_75t_L g398 ( 
.A1(n_376),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_277),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_314),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_335),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_357),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_378),
.B(n_374),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_320),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_329),
.B(n_233),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_238),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

INVx8_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_351),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_378),
.B(n_374),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_239),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_284),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_379),
.B(n_39),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_378),
.B(n_242),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_378),
.B(n_243),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_378),
.B(n_249),
.Y(n_433)
);

OAI22xp33_ASAP7_75t_L g434 ( 
.A1(n_350),
.A2(n_370),
.B1(n_375),
.B2(n_343),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

OAI22xp33_ASAP7_75t_L g436 ( 
.A1(n_375),
.A2(n_312),
.B1(n_311),
.B2(n_307),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_374),
.B(n_296),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_374),
.B(n_298),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_359),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_349),
.B(n_40),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_374),
.B(n_1),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_369),
.B(n_3),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_360),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g452 ( 
.A1(n_345),
.A2(n_43),
.B(n_41),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_371),
.B(n_4),
.Y(n_454)
);

INVx4_ASAP7_75t_SL g455 ( 
.A(n_428),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_385),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_401),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_399),
.B(n_375),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_385),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_404),
.B(n_349),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_438),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_403),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_389),
.B(n_326),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_422),
.B(n_348),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_425),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_400),
.B(n_373),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_380),
.B(n_351),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_395),
.B(n_373),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_404),
.B(n_349),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_417),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_419),
.Y(n_479)
);

INVx3_ASAP7_75t_R g480 ( 
.A(n_423),
.Y(n_480)
);

XOR2x2_ASAP7_75t_L g481 ( 
.A(n_408),
.B(n_333),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_383),
.B(n_362),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_341),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_383),
.B(n_365),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_407),
.B(n_372),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_431),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_371),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_420),
.B(n_372),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_449),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_432),
.B(n_334),
.Y(n_493)
);

XNOR2x2_ASAP7_75t_L g494 ( 
.A(n_398),
.B(n_339),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_362),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_444),
.B(n_369),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_427),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_427),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_444),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_382),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_397),
.B(n_340),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_409),
.B(n_339),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_381),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_390),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_362),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_390),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_454),
.B(n_364),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_450),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_390),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_364),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_398),
.B(n_340),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_395),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_402),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_405),
.B(n_364),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_454),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_428),
.Y(n_519)
);

BUFx5_ASAP7_75t_L g520 ( 
.A(n_428),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_405),
.B(n_369),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

INVx4_ASAP7_75t_SL g523 ( 
.A(n_428),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_428),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_435),
.B(n_369),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_396),
.B(n_340),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_439),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_441),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_442),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_396),
.B(n_354),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_467),
.B(n_388),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_520),
.B(n_388),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_459),
.B(n_388),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_485),
.B(n_388),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_468),
.B(n_415),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_472),
.B(n_415),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_415),
.Y(n_548)
);

AND2x6_ASAP7_75t_SL g549 ( 
.A(n_484),
.B(n_496),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_415),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_463),
.A2(n_428),
.B1(n_386),
.B2(n_451),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_499),
.Y(n_553)
);

O2A1O1Ixp5_ASAP7_75t_L g554 ( 
.A1(n_486),
.A2(n_391),
.B(n_394),
.C(n_451),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_477),
.A2(n_398),
.B1(n_416),
.B2(n_445),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_482),
.B(n_411),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_500),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_502),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_527),
.B(n_411),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_491),
.B(n_414),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_471),
.B(n_354),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_497),
.A2(n_453),
.B(n_426),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_414),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_465),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_466),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_489),
.A2(n_492),
.B1(n_457),
.B2(n_519),
.Y(n_567)
);

INVx8_ASAP7_75t_L g568 ( 
.A(n_489),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_489),
.A2(n_386),
.B1(n_445),
.B2(n_416),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_509),
.B(n_386),
.Y(n_570)
);

O2A1O1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_510),
.A2(n_346),
.B(n_342),
.C(n_344),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_539),
.B(n_458),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_460),
.B(n_421),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_507),
.B(n_421),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_520),
.B(n_519),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_473),
.B(n_429),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_455),
.B(n_398),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_504),
.B(n_429),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_512),
.B(n_384),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_489),
.A2(n_384),
.B1(n_392),
.B2(n_387),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_474),
.B(n_387),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_520),
.B(n_393),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_488),
.A2(n_452),
.B1(n_342),
.B2(n_346),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_503),
.A2(n_392),
.B1(n_413),
.B2(n_410),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_520),
.B(n_393),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_524),
.A2(n_361),
.B1(n_344),
.B2(n_356),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_470),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_514),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_519),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_534),
.Y(n_593)
);

AND2x6_ASAP7_75t_SL g594 ( 
.A(n_462),
.B(n_356),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_520),
.B(n_393),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_479),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_494),
.A2(n_487),
.B1(n_495),
.B2(n_483),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_474),
.B(n_410),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_464),
.A2(n_413),
.B1(n_453),
.B2(n_426),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_538),
.B(n_393),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_455),
.B(n_336),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_538),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_525),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_501),
.B(n_426),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_506),
.B(n_393),
.Y(n_605)
);

A2O1A1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_528),
.A2(n_361),
.B(n_325),
.C(n_368),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_529),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_530),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_508),
.B(n_426),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_513),
.B(n_426),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_549),
.B(n_456),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_573),
.B(n_511),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_591),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_564),
.B(n_556),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_545),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_544),
.A2(n_540),
.B(n_537),
.C(n_536),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_591),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_610),
.A2(n_481),
.B1(n_493),
.B2(n_515),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_562),
.B(n_368),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_590),
.B(n_523),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_545),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_602),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_602),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_577),
.B(n_541),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_601),
.B(n_578),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_570),
.A2(n_452),
.B1(n_533),
.B2(n_532),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_592),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_570),
.B(n_516),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_568),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_523),
.Y(n_634)
);

BUFx4f_ASAP7_75t_L g635 ( 
.A(n_572),
.Y(n_635)
);

OAI21xp33_ASAP7_75t_L g636 ( 
.A1(n_597),
.A2(n_535),
.B(n_531),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_607),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_592),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_568),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_572),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_593),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_604),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_R g643 ( 
.A(n_601),
.B(n_522),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_607),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_594),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_546),
.B(n_505),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_547),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_553),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_557),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_599),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_558),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_558),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_589),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_579),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_589),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_578),
.B(n_336),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_596),
.B(n_475),
.Y(n_658)
);

BUFx8_ASAP7_75t_L g659 ( 
.A(n_603),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_583),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_548),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_574),
.B(n_490),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_593),
.Y(n_665)
);

AOI21xp33_ASAP7_75t_L g666 ( 
.A1(n_571),
.A2(n_452),
.B(n_336),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_608),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_559),
.B(n_526),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_560),
.B(n_526),
.Y(n_669)
);

BUFx8_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_566),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_576),
.B(n_526),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_575),
.B(n_526),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_576),
.B(n_325),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_606),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_675),
.A2(n_563),
.B(n_554),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_635),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_631),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_635),
.Y(n_679)
);

AO31x2_ASAP7_75t_L g680 ( 
.A1(n_618),
.A2(n_555),
.A3(n_606),
.B(n_551),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_615),
.B(n_588),
.Y(n_681)
);

AOI21xp33_ASAP7_75t_L g682 ( 
.A1(n_651),
.A2(n_585),
.B(n_561),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_615),
.B(n_567),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_658),
.A2(n_542),
.B(n_609),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_628),
.B(n_598),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_628),
.B(n_580),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_651),
.A2(n_569),
.B1(n_552),
.B2(n_568),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_658),
.A2(n_542),
.B(n_673),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_673),
.A2(n_581),
.B(n_600),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_633),
.Y(n_690)
);

BUFx2_ASAP7_75t_SL g691 ( 
.A(n_617),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_626),
.B(n_633),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_632),
.A2(n_605),
.B(n_582),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_640),
.Y(n_694)
);

OA21x2_ASAP7_75t_L g695 ( 
.A1(n_630),
.A2(n_394),
.B(n_391),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_632),
.A2(n_587),
.B(n_584),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_659),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_621),
.B(n_363),
.C(n_360),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_648),
.A2(n_587),
.B(n_584),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_623),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_648),
.A2(n_595),
.B(n_453),
.Y(n_701)
);

BUFx4_ASAP7_75t_SL g702 ( 
.A(n_645),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_637),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_660),
.B(n_595),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_659),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_647),
.A2(n_453),
.B(n_430),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_670),
.Y(n_708)
);

AOI21xp33_ASAP7_75t_L g709 ( 
.A1(n_643),
.A2(n_611),
.B(n_620),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_669),
.A2(n_480),
.B(n_453),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_622),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_669),
.A2(n_430),
.B(n_46),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_618),
.A2(n_430),
.B(n_363),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_611),
.B(n_363),
.C(n_360),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_647),
.A2(n_430),
.B(n_363),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_660),
.B(n_363),
.Y(n_716)
);

NAND2x1_ASAP7_75t_L g717 ( 
.A(n_619),
.B(n_430),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_613),
.A2(n_630),
.B(n_666),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_613),
.A2(n_48),
.B(n_44),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_638),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_720)
);

NOR2x1_ASAP7_75t_L g721 ( 
.A(n_642),
.B(n_49),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_666),
.A2(n_52),
.B(n_51),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_636),
.A2(n_57),
.B(n_53),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_670),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_667),
.A2(n_634),
.B(n_655),
.C(n_627),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_622),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_657),
.B(n_6),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_671),
.B(n_7),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_646),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_663),
.A2(n_60),
.B(n_59),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_672),
.A2(n_63),
.B(n_61),
.Y(n_731)
);

AO21x1_ASAP7_75t_L g732 ( 
.A1(n_643),
.A2(n_7),
.B(n_8),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_644),
.B(n_653),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_634),
.B(n_65),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_616),
.A2(n_69),
.B(n_68),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_672),
.A2(n_72),
.B(n_70),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_668),
.B(n_203),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_629),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_689),
.A2(n_625),
.B(n_624),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_703),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_725),
.A2(n_650),
.B1(n_654),
.B2(n_656),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_709),
.A2(n_652),
.B(n_661),
.C(n_674),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_694),
.B(n_664),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_702),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_712),
.A2(n_641),
.B(n_665),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_679),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_718),
.A2(n_626),
.B(n_674),
.Y(n_747)
);

AOI21x1_ASAP7_75t_SL g748 ( 
.A1(n_686),
.A2(n_681),
.B(n_683),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_722),
.A2(n_732),
.A3(n_699),
.B(n_701),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_682),
.A2(n_626),
.B(n_641),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_682),
.A2(n_685),
.B(n_704),
.Y(n_751)
);

AOI211x1_ASAP7_75t_L g752 ( 
.A1(n_720),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_720),
.A2(n_668),
.B(n_619),
.C(n_629),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_706),
.B(n_629),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_SL g756 ( 
.A1(n_687),
.A2(n_639),
.B(n_633),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_716),
.A2(n_626),
.B(n_633),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_728),
.A2(n_629),
.B(n_662),
.C(n_12),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_734),
.A2(n_738),
.B1(n_737),
.B2(n_726),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_677),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_691),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_723),
.A2(n_639),
.B(n_614),
.C(n_612),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_733),
.Y(n_763)
);

OA22x2_ASAP7_75t_L g764 ( 
.A1(n_734),
.A2(n_629),
.B1(n_10),
.B2(n_12),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_729),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_714),
.A2(n_662),
.B(n_612),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_687),
.A2(n_639),
.B(n_662),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_676),
.A2(n_662),
.B(n_639),
.Y(n_768)
);

O2A1O1Ixp5_ASAP7_75t_SL g769 ( 
.A1(n_713),
.A2(n_662),
.B(n_13),
.C(n_14),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_711),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_713),
.A2(n_612),
.B(n_614),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_727),
.B(n_614),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_711),
.B(n_612),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_700),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_714),
.A2(n_9),
.B(n_13),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_698),
.A2(n_202),
.B(n_136),
.Y(n_776)
);

AOI21xp33_ASAP7_75t_L g777 ( 
.A1(n_698),
.A2(n_14),
.B(n_15),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_737),
.Y(n_778)
);

AOI221xp5_ASAP7_75t_SL g779 ( 
.A1(n_719),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_779)
);

AO31x2_ASAP7_75t_L g780 ( 
.A1(n_715),
.A2(n_16),
.A3(n_17),
.B(n_18),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_721),
.B(n_73),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_711),
.B(n_19),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_690),
.B(n_730),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_697),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_731),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_690),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_708),
.B(n_76),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_705),
.B(n_78),
.Y(n_789)
);

O2A1O1Ixp5_ASAP7_75t_L g790 ( 
.A1(n_736),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_724),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_692),
.B(n_79),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_710),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_707),
.A2(n_201),
.B(n_147),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_684),
.A2(n_146),
.B(n_197),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_693),
.A2(n_688),
.B(n_735),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_680),
.B(n_24),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_692),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_798)
);

AO31x2_ASAP7_75t_L g799 ( 
.A1(n_680),
.A2(n_28),
.A3(n_29),
.B(n_30),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_717),
.B(n_84),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_695),
.A2(n_152),
.B(n_196),
.Y(n_801)
);

AOI21x1_ASAP7_75t_L g802 ( 
.A1(n_695),
.A2(n_151),
.B(n_195),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_686),
.A2(n_29),
.B(n_30),
.Y(n_803)
);

NOR2x1_ASAP7_75t_R g804 ( 
.A(n_679),
.B(n_199),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_685),
.B(n_31),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_718),
.A2(n_153),
.B(n_194),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_677),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_767),
.B(n_85),
.Y(n_808)
);

BUFx4f_ASAP7_75t_SL g809 ( 
.A(n_746),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_803),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_764),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_761),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_775),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_755),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_778),
.A2(n_781),
.B1(n_791),
.B2(n_754),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_805),
.A2(n_37),
.B1(n_86),
.B2(n_87),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_763),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_765),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_799),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_782),
.B(n_88),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_781),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_781),
.A2(n_95),
.B1(n_97),
.B2(n_99),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_772),
.Y(n_824)
);

BUFx8_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_743),
.Y(n_826)
);

INVx6_ASAP7_75t_L g827 ( 
.A(n_788),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_781),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_799),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_799),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_751),
.B(n_797),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_740),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_774),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_747),
.A2(n_105),
.B(n_106),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_807),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_780),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_770),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_785),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_777),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_787),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_SL g842 ( 
.A1(n_789),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_800),
.Y(n_843)
);

BUFx12f_ASAP7_75t_L g844 ( 
.A(n_788),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_773),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_759),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_752),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_847)
);

BUFx8_ASAP7_75t_L g848 ( 
.A(n_804),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_739),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_780),
.Y(n_850)
);

CKINVDCx11_ASAP7_75t_R g851 ( 
.A(n_800),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_786),
.A2(n_798),
.B1(n_756),
.B2(n_742),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_806),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_853)
);

CKINVDCx11_ASAP7_75t_R g854 ( 
.A(n_793),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_784),
.Y(n_855)
);

CKINVDCx6p67_ASAP7_75t_R g856 ( 
.A(n_748),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_SL g857 ( 
.A1(n_792),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_779),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_776),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_750),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_SL g861 ( 
.A1(n_758),
.A2(n_148),
.B(n_154),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_741),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_768),
.B(n_160),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_783),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_745),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_771),
.B(n_162),
.Y(n_866)
);

BUFx5_ASAP7_75t_L g867 ( 
.A(n_795),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_864),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_815),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_820),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_855),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_829),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_855),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_819),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_824),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_831),
.B(n_749),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_830),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_855),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_849),
.A2(n_796),
.B(n_802),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_824),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_836),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_865),
.B(n_749),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_837),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_831),
.B(n_850),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_841),
.B(n_833),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_854),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_818),
.B(n_826),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_867),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_813),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_867),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_832),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_863),
.Y(n_892)
);

BUFx2_ASAP7_75t_SL g893 ( 
.A(n_843),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_863),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_834),
.A2(n_766),
.B(n_801),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_867),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_867),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_843),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_867),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_856),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_808),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_866),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_845),
.B(n_749),
.Y(n_903)
);

AO21x1_ASAP7_75t_L g904 ( 
.A1(n_852),
.A2(n_753),
.B(n_794),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_808),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_866),
.Y(n_906)
);

BUFx5_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_SL g908 ( 
.A1(n_852),
.A2(n_790),
.B1(n_757),
.B2(n_769),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_816),
.B(n_821),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_827),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_834),
.A2(n_762),
.B(n_165),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_838),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_847),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_876),
.B(n_835),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_868),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_884),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_868),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_901),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_881),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_881),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_911),
.A2(n_861),
.B(n_817),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_887),
.B(n_861),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_883),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

AO21x2_ASAP7_75t_L g925 ( 
.A1(n_899),
.A2(n_879),
.B(n_890),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_876),
.B(n_884),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_887),
.B(n_875),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_870),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_870),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_890),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_872),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_908),
.A2(n_817),
.B(n_811),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_872),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_884),
.B(n_835),
.Y(n_934)
);

NOR2x1_ASAP7_75t_SL g935 ( 
.A(n_893),
.B(n_844),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_869),
.Y(n_936)
);

AO21x1_ASAP7_75t_SL g937 ( 
.A1(n_913),
.A2(n_814),
.B(n_828),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_869),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_877),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_890),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_885),
.Y(n_941)
);

AO21x2_ASAP7_75t_L g942 ( 
.A1(n_899),
.A2(n_847),
.B(n_812),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_877),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_874),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_884),
.B(n_835),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_874),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_880),
.B(n_827),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_919),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_926),
.B(n_888),
.Y(n_949)
);

BUFx2_ASAP7_75t_SL g950 ( 
.A(n_918),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_919),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_926),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_927),
.B(n_903),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_920),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_941),
.B(n_888),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_920),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_930),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_941),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_916),
.B(n_882),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_923),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_918),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_923),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_924),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_941),
.B(n_896),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_924),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_936),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_916),
.B(n_896),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_936),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_918),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_945),
.B(n_885),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_928),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_951),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_952),
.B(n_914),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_951),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_949),
.B(n_914),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_949),
.B(n_958),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_951),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_968),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_958),
.B(n_945),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_953),
.B(n_922),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_948),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_969),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_959),
.B(n_938),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_960),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_955),
.B(n_934),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_960),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_960),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_948),
.Y(n_988)
);

AND2x4_ASAP7_75t_SL g989 ( 
.A(n_976),
.B(n_898),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_988),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_973),
.B(n_955),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_973),
.B(n_970),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_980),
.B(n_966),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_982),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_982),
.B(n_935),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_985),
.B(n_889),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_976),
.B(n_964),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_983),
.B(n_934),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_988),
.Y(n_999)
);

AND2x4_ASAP7_75t_SL g1000 ( 
.A(n_979),
.B(n_898),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_985),
.B(n_967),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_993),
.B(n_983),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_990),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_992),
.B(n_975),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_SL g1005 ( 
.A(n_996),
.B(n_921),
.C(n_932),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_990),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_997),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_999),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_994),
.B(n_975),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_995),
.B(n_979),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1005),
.B(n_994),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_1010),
.B(n_995),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_SL g1013 ( 
.A(n_1010),
.B(n_900),
.Y(n_1013)
);

OAI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_1009),
.A2(n_900),
.B1(n_886),
.B2(n_947),
.C(n_910),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1004),
.B(n_991),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1007),
.B(n_1001),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1007),
.A2(n_995),
.B1(n_989),
.B2(n_1000),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1011),
.B(n_1015),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1016),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1012),
.B(n_989),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1017),
.B(n_1000),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_1014),
.B(n_1013),
.Y(n_1022)
);

NAND2x1_ASAP7_75t_L g1023 ( 
.A(n_1012),
.B(n_1006),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_1012),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1012),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1016),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1011),
.B(n_1002),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_1024),
.B(n_810),
.Y(n_1028)
);

AOI32xp33_ASAP7_75t_L g1029 ( 
.A1(n_1022),
.A2(n_1003),
.A3(n_1008),
.B1(n_886),
.B2(n_997),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_1023),
.Y(n_1030)
);

AOI211xp5_ASAP7_75t_L g1031 ( 
.A1(n_1018),
.A2(n_1003),
.B(n_886),
.C(n_904),
.Y(n_1031)
);

NAND4xp25_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_910),
.C(n_842),
.D(n_909),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1025),
.B(n_998),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1027),
.A2(n_978),
.B1(n_959),
.B2(n_950),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1019),
.B(n_981),
.Y(n_1035)
);

AOI32xp33_ASAP7_75t_L g1036 ( 
.A1(n_1021),
.A2(n_909),
.A3(n_969),
.B1(n_913),
.B2(n_842),
.Y(n_1036)
);

OAI31xp33_ASAP7_75t_L g1037 ( 
.A1(n_1030),
.A2(n_1019),
.A3(n_1026),
.B(n_1020),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1033),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_1028),
.B(n_809),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1035),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1032),
.B(n_839),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_1029),
.B(n_961),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1031),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1036),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1043),
.A2(n_969),
.B1(n_961),
.B2(n_987),
.Y(n_1046)
);

AOI221xp5_ASAP7_75t_L g1047 ( 
.A1(n_1044),
.A2(n_904),
.B1(n_859),
.B2(n_961),
.C(n_942),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_1037),
.A2(n_961),
.B1(n_942),
.B2(n_822),
.C(n_823),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1038),
.Y(n_1049)
);

AOI211xp5_ASAP7_75t_L g1050 ( 
.A1(n_1045),
.A2(n_961),
.B(n_905),
.C(n_906),
.Y(n_1050)
);

AOI332xp33_ASAP7_75t_L g1051 ( 
.A1(n_1040),
.A2(n_1045),
.A3(n_1042),
.B1(n_1041),
.B2(n_1039),
.B3(n_987),
.C1(n_977),
.C2(n_984),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_1037),
.A2(n_825),
.B(n_848),
.Y(n_1052)
);

AOI221xp5_ASAP7_75t_L g1053 ( 
.A1(n_1044),
.A2(n_961),
.B1(n_942),
.B2(n_977),
.C(n_950),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_1049),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1046),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1050),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_1052),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1051),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1053),
.B(n_935),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1047),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1049),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_1049),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1049),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_1063),
.B(n_825),
.C(n_857),
.Y(n_1065)
);

NAND4xp25_ASAP7_75t_L g1066 ( 
.A(n_1057),
.B(n_846),
.C(n_898),
.D(n_860),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1058),
.A2(n_851),
.B1(n_907),
.B2(n_848),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_L g1068 ( 
.A(n_1063),
.B(n_853),
.C(n_840),
.Y(n_1068)
);

AOI211xp5_ASAP7_75t_L g1069 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_1060),
.C(n_1062),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1063),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_1061),
.B(n_898),
.C(n_906),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_1054),
.B(n_905),
.C(n_902),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_1064),
.B(n_892),
.C(n_907),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_L g1074 ( 
.A(n_1064),
.B(n_907),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_1059),
.B(n_902),
.C(n_894),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_SL g1076 ( 
.A(n_1069),
.B(n_862),
.C(n_892),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1070),
.B(n_972),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_1074),
.B(n_972),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1067),
.B(n_974),
.Y(n_1079)
);

NAND4xp25_ASAP7_75t_SL g1080 ( 
.A(n_1075),
.B(n_986),
.C(n_984),
.D(n_974),
.Y(n_1080)
);

NAND4xp25_ASAP7_75t_L g1081 ( 
.A(n_1071),
.B(n_894),
.C(n_912),
.D(n_878),
.Y(n_1081)
);

NAND4xp25_ASAP7_75t_SL g1082 ( 
.A(n_1065),
.B(n_986),
.C(n_912),
.D(n_967),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_1073),
.B(n_838),
.C(n_918),
.Y(n_1083)
);

OAI211xp5_ASAP7_75t_SL g1084 ( 
.A1(n_1078),
.A2(n_1068),
.B(n_1072),
.C(n_1066),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1081),
.A2(n_893),
.B1(n_918),
.B2(n_963),
.C(n_962),
.Y(n_1085)
);

NOR4xp25_ASAP7_75t_SL g1086 ( 
.A(n_1076),
.B(n_971),
.C(n_965),
.D(n_963),
.Y(n_1086)
);

AOI211xp5_ASAP7_75t_L g1087 ( 
.A1(n_1082),
.A2(n_901),
.B(n_838),
.C(n_894),
.Y(n_1087)
);

AOI211xp5_ASAP7_75t_L g1088 ( 
.A1(n_1077),
.A2(n_901),
.B(n_894),
.C(n_954),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1079),
.B(n_907),
.Y(n_1089)
);

OAI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1083),
.A2(n_971),
.B(n_965),
.C(n_954),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1080),
.B(n_907),
.Y(n_1091)
);

XNOR2xp5_ASAP7_75t_L g1092 ( 
.A(n_1076),
.B(n_164),
.Y(n_1092)
);

INVxp33_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1089),
.A2(n_957),
.B1(n_901),
.B2(n_962),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1084),
.B(n_907),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_R g1096 ( 
.A(n_1091),
.B(n_166),
.Y(n_1096)
);

NAND4xp75_ASAP7_75t_L g1097 ( 
.A(n_1085),
.B(n_1086),
.C(n_1087),
.D(n_1088),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1090),
.B(n_956),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1084),
.B(n_167),
.C(n_168),
.Y(n_1099)
);

AOI322xp5_ASAP7_75t_L g1100 ( 
.A1(n_1085),
.A2(n_957),
.A3(n_964),
.B1(n_937),
.B2(n_956),
.C1(n_901),
.C2(n_871),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1092),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1089),
.B(n_957),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1095),
.B(n_907),
.Y(n_1103)
);

XNOR2x1_ASAP7_75t_L g1104 ( 
.A(n_1101),
.B(n_169),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1099),
.B(n_957),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1093),
.B(n_907),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1102),
.B(n_901),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1098),
.B(n_907),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_1097),
.B(n_873),
.C(n_174),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1096),
.B(n_937),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1102),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_1100),
.B(n_878),
.Y(n_1112)
);

NAND4xp25_ASAP7_75t_L g1113 ( 
.A(n_1094),
.B(n_871),
.C(n_873),
.D(n_891),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1095),
.A2(n_940),
.B1(n_930),
.B2(n_917),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_1101),
.B(n_873),
.C(n_175),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_1104),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1110),
.B(n_915),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1109),
.A2(n_873),
.B1(n_930),
.B2(n_940),
.Y(n_1118)
);

NOR4xp25_ASAP7_75t_L g1119 ( 
.A(n_1111),
.B(n_915),
.C(n_917),
.D(n_931),
.Y(n_1119)
);

OA22x2_ASAP7_75t_L g1120 ( 
.A1(n_1105),
.A2(n_930),
.B1(n_940),
.B2(n_943),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1108),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_1106),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1103),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_1115),
.B(n_944),
.C(n_891),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1116),
.A2(n_1112),
.B1(n_1107),
.B2(n_1114),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1122),
.A2(n_1113),
.B1(n_940),
.B2(n_925),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1121),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1123),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1118),
.A2(n_925),
.B1(n_928),
.B2(n_943),
.Y(n_1129)
);

AO22x2_ASAP7_75t_L g1130 ( 
.A1(n_1117),
.A2(n_931),
.B1(n_939),
.B2(n_933),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1120),
.Y(n_1131)
);

AOI311xp33_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_1119),
.A3(n_1124),
.B(n_939),
.C(n_933),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1127),
.A2(n_929),
.B1(n_944),
.B2(n_179),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1131),
.A2(n_895),
.B(n_897),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1133),
.B(n_1128),
.Y(n_1135)
);

OR3x1_ASAP7_75t_L g1136 ( 
.A(n_1135),
.B(n_1132),
.C(n_1126),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_SL g1137 ( 
.A(n_1136),
.B(n_1134),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_1129),
.B1(n_1130),
.B2(n_925),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1137),
.A2(n_929),
.B1(n_885),
.B2(n_897),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1137),
.A2(n_946),
.B1(n_938),
.B2(n_885),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_1140),
.B(n_170),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1138),
.A2(n_178),
.B(n_180),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1139),
.B(n_181),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_1143),
.B(n_1141),
.Y(n_1144)
);

AO21x2_ASAP7_75t_L g1145 ( 
.A1(n_1142),
.A2(n_183),
.B(n_184),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1145),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_1146)
);

AOI211xp5_ASAP7_75t_L g1147 ( 
.A1(n_1146),
.A2(n_1144),
.B(n_190),
.C(n_191),
.Y(n_1147)
);


endmodule