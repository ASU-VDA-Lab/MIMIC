module fake_jpeg_3424_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_5),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_42),
.B(n_58),
.Y(n_91)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_44),
.A2(n_72),
.B(n_69),
.Y(n_112)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_65),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_64),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_33),
.B(n_2),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_71),
.Y(n_98)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_76),
.Y(n_104)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_79),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_36),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_81),
.B(n_96),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_27),
.B1(n_21),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_84),
.A2(n_97),
.B1(n_34),
.B2(n_41),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_27),
.B1(n_21),
.B2(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_15),
.B1(n_107),
.B2(n_93),
.Y(n_135)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_53),
.B(n_39),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_110),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_38),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_43),
.B(n_19),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_35),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_35),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_20),
.B1(n_19),
.B2(n_8),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_122),
.B1(n_8),
.B2(n_10),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_46),
.B(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_120),
.B(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_52),
.B(n_2),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_83),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_3),
.Y(n_123)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_132),
.B1(n_143),
.B2(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_10),
.C(n_11),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_163),
.C(n_148),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_11),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_14),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_144),
.Y(n_167)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_93),
.B1(n_108),
.B2(n_85),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_80),
.B1(n_124),
.B2(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_86),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_119),
.B(n_122),
.C(n_111),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_162),
.B(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_153),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_115),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_157),
.Y(n_175)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_82),
.A2(n_117),
.B1(n_109),
.B2(n_118),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_158),
.B1(n_157),
.B2(n_134),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_82),
.B1(n_117),
.B2(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_115),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_125),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_87),
.A2(n_84),
.B1(n_89),
.B2(n_120),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_162),
.B1(n_143),
.B2(n_132),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_24),
.B1(n_28),
.B2(n_54),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_156),
.B(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_140),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_164),
.B1(n_183),
.B2(n_179),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_174),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_161),
.C(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_165),
.B1(n_178),
.B2(n_185),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_131),
.B(n_127),
.C(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_152),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_138),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_133),
.B(n_149),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_138),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_194),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_128),
.B(n_126),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_193),
.A2(n_211),
.B(n_209),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_158),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_199),
.C(n_204),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_206),
.B(n_207),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_155),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_155),
.B1(n_171),
.B2(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_208),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_173),
.B1(n_184),
.B2(n_167),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_192),
.Y(n_217)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_169),
.B(n_177),
.C(n_180),
.D(n_198),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_219),
.B(n_193),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_180),
.C(n_177),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_195),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_177),
.B1(n_197),
.B2(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_200),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_194),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_205),
.B(n_203),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_203),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_202),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_225),
.B(n_229),
.Y(n_230)
);

BUFx12f_ASAP7_75t_SL g226 ( 
.A(n_218),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_214),
.B(n_213),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_222),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_220),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_216),
.C(n_212),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_212),
.C(n_194),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_234),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_237),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_238),
.B(n_239),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_231),
.B(n_230),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_230),
.Y(n_243)
);


endmodule