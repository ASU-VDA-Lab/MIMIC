module fake_jpeg_13156_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_12),
.B(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_1),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_77),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_50),
.B1(n_47),
.B2(n_53),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_73),
.B1(n_45),
.B2(n_3),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_52),
.B1(n_49),
.B2(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_41),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_1),
.Y(n_88)
);

NOR2xp67_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_5),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_103),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_21),
.C(n_9),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.C(n_106),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_23),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_30),
.C(n_14),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_6),
.B(n_15),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_16),
.B(n_17),
.Y(n_111)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_115),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_18),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_29),
.B(n_31),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_97),
.C(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_107),
.B1(n_101),
.B2(n_110),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_115),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_120),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_123),
.B(n_96),
.Y(n_127)
);

AOI21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_119),
.B(n_107),
.Y(n_128)
);

NAND4xp25_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_101),
.C(n_117),
.D(n_34),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_33),
.Y(n_130)
);


endmodule