module fake_jpeg_13787_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_57),
.B1(n_65),
.B2(n_34),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_19),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g105 ( 
.A(n_56),
.B(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_19),
.B1(n_24),
.B2(n_28),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_71),
.B1(n_20),
.B2(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_38),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_30),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_24),
.B1(n_22),
.B2(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_36),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_31),
.B1(n_20),
.B2(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_87),
.B1(n_94),
.B2(n_61),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_78),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_29),
.B1(n_60),
.B2(n_54),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_85),
.B(n_97),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_46),
.B1(n_40),
.B2(n_39),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_44),
.B(n_49),
.C(n_46),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_54),
.B1(n_60),
.B2(n_74),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_37),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_27),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_22),
.B1(n_35),
.B2(n_29),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_105),
.B(n_25),
.Y(n_110)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_29),
.B1(n_34),
.B2(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_25),
.Y(n_121)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_127),
.B1(n_103),
.B2(n_100),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_117),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_32),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_61),
.B1(n_74),
.B2(n_60),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_129),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_126),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_87),
.B1(n_75),
.B2(n_84),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_58),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_140),
.Y(n_170)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_86),
.B1(n_88),
.B2(n_92),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_153),
.B1(n_166),
.B2(n_108),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_147),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_124),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_159),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_105),
.B(n_81),
.C(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_165),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_161),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_105),
.B(n_93),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_121),
.B(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_96),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_89),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_154),
.B(n_115),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_105),
.C(n_93),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_162),
.C(n_126),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_93),
.B(n_80),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_91),
.B(n_115),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_133),
.C(n_111),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_33),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_111),
.B(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_91),
.B1(n_104),
.B2(n_90),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_121),
.B(n_135),
.C(n_120),
.D(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_168),
.B(n_180),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_142),
.B(n_143),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_176),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_160),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_106),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_181),
.B(n_184),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_146),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_161),
.B1(n_138),
.B2(n_141),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_120),
.B(n_104),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_183),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_119),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_119),
.B1(n_117),
.B2(n_104),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_190),
.B1(n_196),
.B2(n_166),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_195),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_117),
.B1(n_113),
.B2(n_122),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_106),
.B(n_83),
.C(n_134),
.D(n_101),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_192),
.B(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_134),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_151),
.A2(n_82),
.B1(n_134),
.B2(n_58),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_147),
.B(n_36),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_82),
.B1(n_25),
.B2(n_26),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_26),
.B1(n_58),
.B2(n_53),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_204),
.B1(n_225),
.B2(n_228),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_167),
.B1(n_164),
.B2(n_186),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_173),
.B(n_170),
.C(n_201),
.D(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_164),
.B(n_165),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_164),
.B(n_167),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_212),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_148),
.Y(n_217)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_226),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_224),
.A2(n_199),
.B1(n_185),
.B2(n_198),
.Y(n_256)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_53),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_95),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_178),
.A2(n_95),
.B1(n_66),
.B2(n_55),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_196),
.B1(n_199),
.B2(n_187),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_66),
.B1(n_9),
.B2(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_192),
.Y(n_248)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_243),
.B1(n_248),
.B2(n_252),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_209),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_171),
.B1(n_179),
.B2(n_180),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_256),
.B1(n_204),
.B2(n_203),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_171),
.Y(n_243)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_214),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_66),
.B(n_8),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_193),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_217),
.C(n_218),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_208),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_185),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_229),
.B(n_197),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_198),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_205),
.B(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_276),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_264),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_221),
.B1(n_224),
.B2(n_211),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_215),
.C(n_212),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_266),
.C(n_269),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_210),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_210),
.C(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_231),
.B1(n_168),
.B2(n_230),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_199),
.C(n_177),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_177),
.B1(n_188),
.B2(n_66),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_66),
.C(n_9),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_275),
.C(n_276),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_234),
.A2(n_16),
.B(n_15),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_243),
.B(n_15),
.CI(n_13),
.CON(n_277),
.SN(n_277)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_11),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_273),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_288),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_238),
.C(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_284),
.B(n_286),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_236),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_267),
.A2(n_238),
.B1(n_248),
.B2(n_232),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_292),
.B1(n_295),
.B2(n_256),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_254),
.C(n_251),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_294),
.Y(n_299)
);

NAND4xp25_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_233),
.C(n_245),
.D(n_250),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_261),
.B(n_271),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_297),
.A2(n_306),
.B(n_12),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_249),
.B(n_260),
.C(n_245),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_302),
.B(n_293),
.Y(n_312)
);

A2O1A1O1Ixp25_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_249),
.B(n_269),
.C(n_259),
.D(n_264),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_279),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_308),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_274),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_277),
.B(n_270),
.C(n_235),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_277),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_1),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_13),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_294),
.B1(n_285),
.B2(n_293),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_318),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_3),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_12),
.B1(n_9),
.B2(n_2),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_320),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_317),
.B(n_321),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_0),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_299),
.A2(n_1),
.B(n_3),
.Y(n_321)
);

INVx11_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_322),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_302),
.C(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_323),
.B(n_325),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_3),
.B(n_4),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_329),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_4),
.B(n_5),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_310),
.B1(n_320),
.B2(n_5),
.Y(n_333)
);

AOI31xp67_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_5),
.A3(n_6),
.B(n_319),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_5),
.B(n_6),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_6),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_330),
.B(n_324),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_328),
.B(n_326),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_332),
.C(n_338),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_331),
.B(n_334),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_6),
.Y(n_343)
);


endmodule