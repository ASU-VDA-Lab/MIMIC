module fake_netlist_5_1607_n_2560 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2560);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2560;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2193;
wire n_2052;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_1587;
wire n_680;
wire n_1473;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2195;
wire n_2529;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2545;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_2339;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_2519;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2282;
wire n_2002;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_2494;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_257),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_204),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_567),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_225),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_181),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_482),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_106),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_57),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_206),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_15),
.Y(n_595)
);

CKINVDCx14_ASAP7_75t_R g596 ( 
.A(n_531),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_411),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_285),
.Y(n_598)
);

BUFx5_ASAP7_75t_L g599 ( 
.A(n_107),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_501),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_338),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_191),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_303),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_119),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_171),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_104),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_62),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_155),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_379),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_406),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_314),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_269),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_223),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_502),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_121),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_180),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_50),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_54),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_174),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_98),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_506),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_513),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_178),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_177),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_125),
.Y(n_626)
);

CKINVDCx16_ASAP7_75t_R g627 ( 
.A(n_73),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_48),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_246),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_444),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_303),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_282),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_178),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_560),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_566),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_453),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_122),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_524),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_240),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_541),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_122),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_359),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_40),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_55),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_204),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_129),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_320),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_448),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_225),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_164),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_254),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_83),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_313),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_42),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_98),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_400),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_171),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_22),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_441),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_284),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_477),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_103),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_459),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_182),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_76),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_344),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_529),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_199),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_184),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_422),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_387),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_492),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_304),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_110),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_266),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_488),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_68),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_443),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_25),
.Y(n_680)
);

INVxp33_ASAP7_75t_L g681 ( 
.A(n_447),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_87),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_164),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_54),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_497),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_577),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_192),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_407),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_364),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_9),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_224),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_468),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_130),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_175),
.Y(n_694)
);

BUFx10_ASAP7_75t_L g695 ( 
.A(n_559),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_411),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_520),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_572),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_219),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_383),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_221),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_110),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_210),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_19),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_460),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_479),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_80),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_449),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_189),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_563),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_489),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_292),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_456),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_231),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_445),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_14),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_569),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_191),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_124),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_369),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_233),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_151),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_24),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_565),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_542),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_536),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_237),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_179),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_129),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_450),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_410),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_253),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_442),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_183),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_333),
.Y(n_735)
);

CKINVDCx16_ASAP7_75t_R g736 ( 
.A(n_447),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_522),
.Y(n_737)
);

CKINVDCx16_ASAP7_75t_R g738 ( 
.A(n_268),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_176),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_284),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_215),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_190),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_527),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_278),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_450),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_117),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_332),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_77),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_78),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_277),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_507),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_422),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_259),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_97),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_410),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_414),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_508),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_86),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_367),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_366),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_296),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_198),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_106),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_40),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_77),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_220),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_317),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_34),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_51),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_331),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_15),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_394),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_499),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_34),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_240),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_65),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_9),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_287),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_316),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_291),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_370),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_46),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_446),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_222),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_294),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_84),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_393),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_571),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_94),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_272),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_67),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_420),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_345),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_104),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_405),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_333),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_229),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_695),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_599),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_627),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_599),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_637),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_599),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_599),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_599),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_599),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_736),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_685),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_599),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_602),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_648),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_648),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_738),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_706),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_590),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_590),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_706),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_604),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_590),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_590),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_748),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_601),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_781),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_601),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_759),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_601),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_601),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_744),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_744),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_744),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_706),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_671),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_585),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_681),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_671),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_773),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_587),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_719),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_723),
.Y(n_839)
);

BUFx2_ASAP7_75t_SL g840 ( 
.A(n_725),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_723),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_746),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_746),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_602),
.Y(n_844)
);

INVxp33_ASAP7_75t_SL g845 ( 
.A(n_595),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_617),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_769),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_744),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_589),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_617),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_706),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_763),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_596),
.Y(n_853)
);

CKINVDCx14_ASAP7_75t_R g854 ( 
.A(n_619),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_763),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_763),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_725),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_592),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_763),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_597),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_603),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_606),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_607),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_611),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_613),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_615),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_664),
.Y(n_867)
);

INVxp33_ASAP7_75t_L g868 ( 
.A(n_620),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_623),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_631),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_586),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_593),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_643),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_595),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_644),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_650),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_712),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_656),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_621),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_657),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_674),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_680),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_689),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_639),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_594),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_706),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_704),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_639),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_652),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_652),
.Y(n_890)
);

INVxp33_ASAP7_75t_L g891 ( 
.A(n_714),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_591),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_718),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_722),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_815),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_815),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_848),
.B(n_664),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_892),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_811),
.B(n_661),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_812),
.B(n_832),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_816),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_852),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_892),
.Y(n_903)
);

AND2x6_ASAP7_75t_L g904 ( 
.A(n_892),
.B(n_591),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_892),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_801),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_836),
.B(n_654),
.Y(n_907)
);

INVx6_ASAP7_75t_L g908 ( 
.A(n_867),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_801),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_814),
.Y(n_910)
);

NOR2x1_ASAP7_75t_L g911 ( 
.A(n_798),
.B(n_654),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_814),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_871),
.B(n_692),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_816),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_879),
.B(n_808),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_819),
.Y(n_916)
);

AND2x6_ASAP7_75t_L g917 ( 
.A(n_817),
.B(n_591),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_874),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_817),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_831),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_831),
.B(n_591),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_853),
.B(n_600),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_799),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_819),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_835),
.B(n_661),
.Y(n_925)
);

NOR2x1_ASAP7_75t_L g926 ( 
.A(n_798),
.B(n_692),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_803),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_820),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_867),
.B(n_622),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_800),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_851),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_820),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_800),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_822),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_822),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_824),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_851),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_824),
.B(n_624),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_826),
.Y(n_939)
);

BUFx12f_ASAP7_75t_L g940 ( 
.A(n_802),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_855),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_856),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_826),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_827),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_827),
.B(n_638),
.Y(n_945)
);

BUFx8_ASAP7_75t_SL g946 ( 
.A(n_810),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_886),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_840),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_828),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_828),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_833),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_840),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_804),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_829),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_829),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_913),
.B(n_830),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_900),
.B(n_913),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_898),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_908),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_906),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_938),
.B(n_805),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_923),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_917),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_918),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_900),
.B(n_834),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_923),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_906),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_923),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_906),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_927),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_927),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_933),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_927),
.Y(n_973)
);

NOR2x1_ASAP7_75t_L g974 ( 
.A(n_911),
.B(n_724),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_938),
.B(n_806),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_906),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_953),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_913),
.B(n_830),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_896),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_946),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_953),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_953),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_909),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_912),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_948),
.B(n_877),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_896),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_901),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_913),
.B(n_859),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_912),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_909),
.B(n_809),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_951),
.A2(n_823),
.B1(n_630),
.B2(n_715),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_909),
.B(n_837),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_909),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_898),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_912),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_912),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_930),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_920),
.B(n_837),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_920),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_920),
.B(n_849),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_901),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_938),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_902),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_902),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_938),
.B(n_751),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_902),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_914),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_941),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_914),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_897),
.B(n_858),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_934),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_934),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_941),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_924),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_910),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_941),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_948),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_898),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_924),
.Y(n_1019)
);

BUFx8_ASAP7_75t_L g1020 ( 
.A(n_940),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_924),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_899),
.B(n_838),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_942),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_930),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_910),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_915),
.B(n_858),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_898),
.Y(n_1027)
);

INVx6_ASAP7_75t_L g1028 ( 
.A(n_945),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_942),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_942),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_924),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_895),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_895),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_916),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_916),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_899),
.B(n_839),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_932),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_922),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_951),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_952),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_1002),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1028),
.A2(n_952),
.B1(n_907),
.B2(n_908),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_984),
.B(n_989),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_1002),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_984),
.B(n_908),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_960),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1032),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_960),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1033),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_957),
.B(n_925),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_957),
.B(n_925),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_1002),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_1028),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_965),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_960),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_1028),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_965),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_967),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1003),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_967),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1026),
.B(n_813),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1038),
.B(n_802),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_967),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_969),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_980),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_1020),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1033),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_1024),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_1022),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_974),
.B(n_911),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1024),
.B(n_857),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_969),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_1010),
.B(n_872),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_969),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_976),
.Y(n_1076)
);

INVx8_ASAP7_75t_L g1077 ( 
.A(n_1005),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_976),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_976),
.Y(n_1079)
);

INVxp33_ASAP7_75t_L g1080 ( 
.A(n_997),
.Y(n_1080)
);

NOR2x1p5_ASAP7_75t_L g1081 ( 
.A(n_1017),
.B(n_940),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_985),
.B(n_885),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_983),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1004),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1004),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_983),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1006),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_964),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_989),
.B(n_908),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_983),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_992),
.B(n_807),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_993),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_993),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_1039),
.B(n_618),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_998),
.B(n_807),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_1028),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_961),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1022),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1036),
.B(n_818),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_993),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1006),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_1036),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1008),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_996),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1034),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1034),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_996),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1035),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1000),
.B(n_821),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_961),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_961),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_999),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_999),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_995),
.B(n_945),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_974),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_999),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1001),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1035),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_SL g1120 ( 
.A(n_959),
.B(n_618),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1001),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1037),
.Y(n_1122)
);

INVxp33_ASAP7_75t_L g1123 ( 
.A(n_972),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_959),
.B(n_825),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1008),
.B(n_945),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1013),
.B(n_926),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1013),
.B(n_926),
.Y(n_1127)
);

NOR2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1020),
.B(n_825),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1040),
.B(n_929),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1001),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_979),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1031),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_961),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1037),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_962),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_956),
.B(n_854),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_979),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_986),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_1040),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_963),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1016),
.B(n_924),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_986),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_987),
.Y(n_1143)
);

INVx6_ASAP7_75t_L g1144 ( 
.A(n_963),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_962),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_987),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_975),
.Y(n_1147)
);

CKINVDCx6p67_ASAP7_75t_R g1148 ( 
.A(n_1020),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1007),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_966),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_966),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1016),
.B(n_928),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_968),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1007),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_968),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1023),
.B(n_928),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_975),
.B(n_845),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1009),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_970),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1023),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1029),
.B(n_810),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1030),
.B(n_928),
.Y(n_1163)
);

AND3x2_ASAP7_75t_L g1164 ( 
.A(n_1030),
.B(n_609),
.C(n_660),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1005),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1009),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1011),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_988),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_991),
.B(n_841),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1135),
.Y(n_1170)
);

INVxp33_ASAP7_75t_SL g1171 ( 
.A(n_1066),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1063),
.B(n_1058),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1080),
.B(n_844),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1135),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1099),
.B(n_844),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1055),
.B(n_978),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1145),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1145),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1151),
.Y(n_1179)
);

XNOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1066),
.B(n_846),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1151),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1099),
.B(n_846),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1055),
.B(n_842),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1042),
.B(n_963),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1069),
.B(n_1020),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1148),
.B(n_630),
.Y(n_1186)
);

XOR2xp5_ASAP7_75t_L g1187 ( 
.A(n_1067),
.B(n_850),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1152),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1051),
.B(n_850),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1152),
.Y(n_1190)
);

AND2x6_ASAP7_75t_L g1191 ( 
.A(n_1165),
.B(n_970),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1154),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1051),
.B(n_843),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1156),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_L g1195 ( 
.A(n_1116),
.B(n_1059),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1069),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1070),
.B(n_1098),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_R g1198 ( 
.A(n_1072),
.B(n_614),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1123),
.B(n_715),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1088),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1139),
.B(n_735),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1156),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1160),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1059),
.B(n_963),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1160),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1052),
.B(n_1070),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1041),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1048),
.Y(n_1208)
);

NAND2xp33_ASAP7_75t_R g1209 ( 
.A(n_1072),
.B(n_588),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1048),
.Y(n_1210)
);

XOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1067),
.B(n_1062),
.Y(n_1211)
);

AND2x6_ASAP7_75t_L g1212 ( 
.A(n_1165),
.B(n_971),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1059),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1050),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1061),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1052),
.B(n_1098),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1068),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1068),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1097),
.B(n_973),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1102),
.B(n_847),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1168),
.B(n_1105),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1105),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_1081),
.B(n_669),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1106),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1106),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1164),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1162),
.B(n_990),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1109),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1109),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1074),
.B(n_973),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1119),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1129),
.B(n_977),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1115),
.A2(n_981),
.B(n_977),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1122),
.Y(n_1234)
);

XOR2xp5_ASAP7_75t_L g1235 ( 
.A(n_1091),
.B(n_1095),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1122),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1134),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1134),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1149),
.B(n_981),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1136),
.B(n_868),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1161),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1169),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1136),
.B(n_891),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1161),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1064),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1082),
.B(n_982),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1148),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1064),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1169),
.B(n_608),
.Y(n_1249)
);

INVxp33_ASAP7_75t_L g1250 ( 
.A(n_1124),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1060),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1090),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1084),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1085),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1087),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1101),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1120),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1128),
.B(n_669),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1149),
.B(n_1042),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1103),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1131),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1094),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_1094),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1120),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1168),
.B(n_712),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1045),
.B(n_982),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1097),
.B(n_634),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1110),
.B(n_625),
.Y(n_1268)
);

XOR2xp5_ASAP7_75t_L g1269 ( 
.A(n_1043),
.B(n_635),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1137),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1137),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1167),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1090),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1167),
.Y(n_1274)
);

INVx4_ASAP7_75t_SL g1275 ( 
.A(n_1071),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1097),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1138),
.Y(n_1277)
);

BUFx5_ASAP7_75t_L g1278 ( 
.A(n_1147),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1158),
.B(n_653),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1045),
.B(n_676),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1047),
.B(n_1005),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1047),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1053),
.B(n_694),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1049),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1049),
.Y(n_1285)
);

XOR2xp5_ASAP7_75t_L g1286 ( 
.A(n_1097),
.B(n_1111),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1126),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1138),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1053),
.B(n_702),
.Y(n_1289)
);

XOR2xp5_ASAP7_75t_L g1290 ( 
.A(n_1097),
.B(n_636),
.Y(n_1290)
);

INVx4_ASAP7_75t_SL g1291 ( 
.A(n_1071),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1166),
.Y(n_1292)
);

XOR2xp5_ASAP7_75t_L g1293 ( 
.A(n_1111),
.B(n_640),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

INVxp33_ASAP7_75t_SL g1296 ( 
.A(n_1127),
.Y(n_1296)
);

XOR2xp5_ASAP7_75t_L g1297 ( 
.A(n_1111),
.B(n_662),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1143),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1056),
.B(n_1005),
.Y(n_1299)
);

XNOR2xp5_ASAP7_75t_L g1300 ( 
.A(n_1046),
.B(n_668),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1146),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1146),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1150),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1111),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1111),
.Y(n_1305)
);

INVxp33_ASAP7_75t_L g1306 ( 
.A(n_1089),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1155),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1155),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1159),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1159),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1071),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1118),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1118),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1121),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1121),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1130),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1130),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1054),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_1065),
.B(n_1014),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1073),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1073),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1075),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1076),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1044),
.A2(n_1012),
.B(n_1011),
.Y(n_1325)
);

XOR2xp5_ASAP7_75t_L g1326 ( 
.A(n_1112),
.B(n_673),
.Y(n_1326)
);

AND2x6_ASAP7_75t_L g1327 ( 
.A(n_1165),
.B(n_1031),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1076),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1078),
.Y(n_1329)
);

NAND2xp33_ASAP7_75t_R g1330 ( 
.A(n_1125),
.B(n_677),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1078),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1054),
.B(n_1031),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1079),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1079),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1083),
.B(n_1019),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1054),
.Y(n_1336)
);

XOR2xp5_ASAP7_75t_L g1337 ( 
.A(n_1112),
.B(n_686),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1083),
.B(n_782),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1086),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1086),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1092),
.Y(n_1341)
);

XNOR2xp5_ASAP7_75t_L g1342 ( 
.A(n_1141),
.B(n_697),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_SL g1343 ( 
.A(n_1077),
.B(n_695),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1112),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1092),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1112),
.B(n_860),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1093),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1093),
.B(n_861),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1196),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1296),
.B(n_1112),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1172),
.B(n_1133),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1200),
.B(n_1133),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1282),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1206),
.B(n_1100),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1284),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1200),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1285),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1227),
.A2(n_1071),
.B1(n_1133),
.B2(n_1057),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1201),
.B(n_1133),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1321),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1171),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1216),
.B(n_1104),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1338),
.B(n_1107),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1240),
.B(n_862),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1170),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1207),
.B(n_1107),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1174),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1177),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1322),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1197),
.B(n_1147),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1323),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1199),
.B(n_1108),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1330),
.A2(n_1071),
.B1(n_1057),
.B2(n_1054),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1178),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1179),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1283),
.B(n_1108),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1257),
.B(n_1113),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1181),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1247),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1287),
.B(n_1113),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1221),
.B(n_1114),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1188),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1190),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1304),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1193),
.B(n_1114),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1176),
.B(n_1117),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1257),
.B(n_1096),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1269),
.A2(n_1268),
.B1(n_1346),
.B2(n_1242),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1189),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1173),
.B(n_1096),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1192),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1208),
.B(n_1132),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1210),
.B(n_1096),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1249),
.A2(n_610),
.B1(n_612),
.B2(n_605),
.C(n_598),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1220),
.B(n_1157),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1324),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1328),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1246),
.A2(n_1077),
.B(n_1163),
.C(n_1153),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1259),
.B(n_1165),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1175),
.B(n_1182),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1243),
.B(n_863),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1300),
.B(n_698),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1329),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1214),
.B(n_1077),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1280),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1331),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1304),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1217),
.B(n_1019),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1226),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1289),
.Y(n_1410)
);

NOR2xp67_ASAP7_75t_L g1411 ( 
.A(n_1342),
.B(n_710),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1218),
.B(n_1021),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1194),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1222),
.B(n_1021),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1279),
.B(n_1265),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1250),
.B(n_626),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1202),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1286),
.A2(n_1319),
.B1(n_1336),
.B2(n_1235),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_SL g1419 ( 
.A(n_1186),
.B(n_695),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1241),
.A2(n_788),
.B1(n_706),
.B2(n_726),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1203),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1244),
.A2(n_726),
.B1(n_705),
.B2(n_713),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1263),
.B(n_864),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1205),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1230),
.A2(n_711),
.B1(n_737),
.B2(n_717),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1333),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1334),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1224),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1232),
.A2(n_761),
.B(n_760),
.C(n_731),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1305),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1262),
.A2(n_786),
.B1(n_612),
.B2(n_605),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1225),
.B(n_932),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1228),
.A2(n_761),
.B(n_760),
.C(n_734),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1229),
.B(n_955),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1231),
.B(n_955),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_L g1436 ( 
.A(n_1305),
.B(n_743),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1234),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1185),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1198),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1186),
.A2(n_610),
.B1(n_616),
.B2(n_598),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1236),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1237),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1238),
.B(n_1339),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1312),
.A2(n_1251),
.B1(n_1254),
.B2(n_1253),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1180),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1183),
.B(n_865),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1290),
.B(n_866),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1340),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1348),
.B(n_869),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1255),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1306),
.B(n_628),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1256),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1341),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1344),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1345),
.B(n_1140),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1260),
.B(n_870),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1185),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1347),
.B(n_1140),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1313),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1314),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1276),
.B(n_757),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1315),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1252),
.B(n_1144),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1233),
.A2(n_741),
.B(n_745),
.C(n_730),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1312),
.B(n_1266),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1316),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1239),
.B(n_705),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1261),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1266),
.A2(n_726),
.B1(n_705),
.B2(n_678),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1185),
.B(n_1144),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1318),
.B(n_1309),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1209),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1213),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1264),
.B(n_629),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1293),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1270),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1297),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1271),
.B(n_886),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1211),
.A2(n_707),
.B1(n_708),
.B2(n_699),
.C(n_616),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1195),
.A2(n_678),
.B1(n_683),
.B2(n_660),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1267),
.A2(n_875),
.B1(n_876),
.B2(n_873),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1191),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1272),
.B(n_632),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1343),
.A2(n_880),
.B1(n_881),
.B2(n_878),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1274),
.B(n_633),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1326),
.B(n_1337),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1219),
.A2(n_753),
.B(n_754),
.C(n_750),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1277),
.B(n_641),
.Y(n_1489)
);

BUFx8_ASAP7_75t_L g1490 ( 
.A(n_1191),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_L g1491 ( 
.A(n_1278),
.B(n_904),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1288),
.B(n_642),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1215),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1187),
.B(n_645),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1191),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1245),
.A2(n_691),
.B1(n_703),
.B2(n_683),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1278),
.B(n_882),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1248),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1292),
.B(n_646),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1294),
.A2(n_708),
.B1(n_709),
.B2(n_707),
.C(n_699),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1273),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1295),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1298),
.B(n_647),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1191),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1301),
.B(n_709),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1302),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1303),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1307),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1308),
.B(n_917),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1310),
.B(n_917),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1258),
.B(n_883),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1311),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1335),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1223),
.B(n_691),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1258),
.B(n_649),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1320),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1281),
.A2(n_893),
.B1(n_894),
.B2(n_887),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1299),
.A2(n_921),
.B1(n_917),
.B2(n_655),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1275),
.B(n_651),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1320),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1258),
.B(n_1223),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1223),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1325),
.B(n_921),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1275),
.B(n_921),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1332),
.B(n_884),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1407),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1415),
.B(n_1291),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1372),
.B(n_1291),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1359),
.B(n_1212),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1450),
.Y(n_1530)
);

BUFx2_ASAP7_75t_SL g1531 ( 
.A(n_1356),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1446),
.B(n_1212),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1398),
.A2(n_1204),
.B(n_1184),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1361),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1360),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1400),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1410),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1395),
.B(n_1212),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1369),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1405),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1439),
.B(n_658),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1452),
.Y(n_1542)
);

NOR2x2_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1471),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1349),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1473),
.B(n_659),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1371),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1364),
.B(n_1327),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1365),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1401),
.B(n_1327),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1523),
.A2(n_905),
.B(n_903),
.Y(n_1550)
);

BUFx12f_ASAP7_75t_L g1551 ( 
.A(n_1522),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1385),
.A2(n_919),
.B(n_910),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1381),
.A2(n_919),
.B(n_910),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1390),
.B(n_758),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1423),
.B(n_884),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1386),
.B(n_767),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1358),
.A2(n_1404),
.B(n_1491),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1392),
.A2(n_919),
.B(n_910),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1388),
.A2(n_770),
.B1(n_772),
.B2(n_768),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1392),
.A2(n_937),
.B(n_931),
.Y(n_1560)
);

OAI321xp33_ASAP7_75t_L g1561 ( 
.A1(n_1440),
.A2(n_774),
.A3(n_777),
.B1(n_784),
.B2(n_780),
.C(n_776),
.Y(n_1561)
);

NAND2xp33_ASAP7_75t_L g1562 ( 
.A(n_1483),
.B(n_1495),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1497),
.A2(n_937),
.B(n_931),
.Y(n_1563)
);

O2A1O1Ixp5_ASAP7_75t_L g1564 ( 
.A1(n_1351),
.A2(n_733),
.B(n_762),
.C(n_703),
.Y(n_1564)
);

BUFx12f_ASAP7_75t_L g1565 ( 
.A(n_1514),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1363),
.B(n_785),
.Y(n_1566)
);

INVx11_ASAP7_75t_L g1567 ( 
.A(n_1490),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1419),
.B(n_779),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1407),
.Y(n_1569)
);

INVx11_ASAP7_75t_L g1570 ( 
.A(n_1490),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1523),
.A2(n_905),
.B(n_903),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1483),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1354),
.B(n_787),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1354),
.B(n_793),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1362),
.B(n_796),
.Y(n_1575)
);

BUFx12f_ASAP7_75t_L g1576 ( 
.A(n_1514),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1362),
.B(n_663),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1513),
.B(n_665),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1367),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1487),
.A2(n_667),
.B1(n_670),
.B2(n_666),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1376),
.A2(n_937),
.B(n_931),
.Y(n_1581)
);

NOR2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1379),
.B(n_779),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1483),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1447),
.B(n_783),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1407),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1389),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1368),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1438),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1374),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1454),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1375),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1411),
.B(n_783),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1475),
.B(n_888),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1494),
.A2(n_675),
.B1(n_679),
.B2(n_672),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1463),
.A2(n_1377),
.B(n_1366),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1409),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1418),
.B(n_888),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1445),
.B(n_682),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1485),
.A2(n_795),
.B(n_789),
.C(n_790),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1503),
.B(n_684),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1449),
.B(n_687),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1476),
.B(n_786),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1465),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1396),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1480),
.A2(n_1468),
.B(n_1429),
.C(n_1394),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1416),
.B(n_789),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1382),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1402),
.B(n_790),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1383),
.B(n_688),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1391),
.B(n_690),
.Y(n_1611)
);

AOI22x1_ASAP7_75t_L g1612 ( 
.A1(n_1516),
.A2(n_792),
.B1(n_794),
.B2(n_791),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1457),
.Y(n_1613)
);

NOR2xp67_ASAP7_75t_L g1614 ( 
.A(n_1478),
.B(n_452),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1525),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1454),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1464),
.A2(n_1387),
.B(n_1451),
.C(n_1517),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1397),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1495),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1413),
.B(n_693),
.Y(n_1620)
);

INVx11_ASAP7_75t_L g1621 ( 
.A(n_1454),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1417),
.B(n_696),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1403),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1421),
.B(n_700),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1424),
.B(n_701),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1428),
.B(n_716),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1444),
.A2(n_1479),
.B(n_1373),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1433),
.A2(n_1350),
.B(n_1444),
.C(n_1484),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1486),
.A2(n_890),
.B(n_889),
.C(n_903),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1437),
.B(n_720),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1441),
.B(n_1442),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_L g1632 ( 
.A(n_1495),
.B(n_791),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1380),
.B(n_721),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1406),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1505),
.B(n_792),
.Y(n_1635)
);

AO21x1_ASAP7_75t_L g1636 ( 
.A1(n_1393),
.A2(n_890),
.B(n_889),
.Y(n_1636)
);

NOR2xp67_ASAP7_75t_L g1637 ( 
.A(n_1489),
.B(n_454),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1456),
.B(n_794),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1426),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1492),
.B(n_1499),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1455),
.A2(n_1458),
.B(n_1399),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1352),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1427),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1469),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1471),
.B(n_455),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1511),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1443),
.B(n_727),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1472),
.A2(n_947),
.B(n_1015),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1472),
.A2(n_947),
.B(n_1025),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1431),
.B(n_728),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1521),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1515),
.B(n_797),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1425),
.B(n_1370),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1432),
.B(n_1434),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1470),
.B(n_729),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1432),
.B(n_732),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1479),
.A2(n_921),
.B(n_904),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1461),
.A2(n_947),
.B(n_1025),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1471),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1434),
.B(n_739),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1488),
.A2(n_797),
.B(n_742),
.C(n_747),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1430),
.B(n_457),
.Y(n_1662)
);

NOR2xp67_ASAP7_75t_L g1663 ( 
.A(n_1519),
.B(n_458),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1504),
.Y(n_1664)
);

INVx11_ASAP7_75t_L g1665 ( 
.A(n_1384),
.Y(n_1665)
);

AND2x6_ASAP7_75t_L g1666 ( 
.A(n_1504),
.B(n_928),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1508),
.B(n_740),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1500),
.B(n_749),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_L g1669 ( 
.A(n_1474),
.B(n_461),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1435),
.B(n_752),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1504),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1422),
.B(n_755),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1384),
.Y(n_1673)
);

AO21x1_ASAP7_75t_L g1674 ( 
.A1(n_1520),
.A2(n_2),
.B(n_1),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_SL g1675 ( 
.A(n_1481),
.B(n_756),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1414),
.A2(n_921),
.B(n_904),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1448),
.B(n_462),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1477),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1435),
.A2(n_921),
.B(n_904),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1436),
.A2(n_1412),
.B(n_1408),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1453),
.Y(n_1681)
);

A2O1A1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1502),
.A2(n_765),
.B(n_766),
.C(n_764),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1506),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_SL g1684 ( 
.A1(n_1459),
.A2(n_465),
.B(n_463),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1507),
.B(n_771),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1536),
.B(n_1482),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1654),
.A2(n_1512),
.B(n_1462),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1595),
.A2(n_1466),
.B(n_1460),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1603),
.B(n_1467),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1493),
.Y(n_1690)
);

A2O1A1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1605),
.A2(n_1617),
.B(n_1628),
.C(n_1653),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1557),
.A2(n_1510),
.B(n_1509),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1606),
.A2(n_1481),
.B(n_1355),
.C(n_1357),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1631),
.Y(n_1694)
);

AO22x1_ASAP7_75t_L g1695 ( 
.A1(n_1650),
.A2(n_778),
.B1(n_775),
.B2(n_1353),
.Y(n_1695)
);

INVx5_ASAP7_75t_L g1696 ( 
.A(n_1526),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1533),
.A2(n_1510),
.B(n_1509),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1680),
.A2(n_1524),
.B(n_1518),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1530),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1627),
.A2(n_1524),
.B(n_1501),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1627),
.A2(n_1498),
.B(n_1420),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1615),
.B(n_1496),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1640),
.A2(n_994),
.B(n_958),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1641),
.A2(n_994),
.B(n_958),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1615),
.B(n_0),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1598),
.B(n_466),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1593),
.B(n_2),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1655),
.A2(n_1668),
.B1(n_1675),
.B2(n_1600),
.Y(n_1708)
);

AO21x1_ASAP7_75t_L g1709 ( 
.A1(n_1554),
.A2(n_3),
.B(n_4),
.Y(n_1709)
);

AOI33xp33_ASAP7_75t_L g1710 ( 
.A1(n_1559),
.A2(n_7),
.A3(n_10),
.B1(n_5),
.B2(n_6),
.B3(n_8),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1535),
.Y(n_1711)
);

AND2x2_ASAP7_75t_SL g1712 ( 
.A(n_1645),
.B(n_5),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1659),
.Y(n_1713)
);

O2A1O1Ixp33_ASAP7_75t_SL g1714 ( 
.A1(n_1528),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1537),
.B(n_467),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1607),
.B(n_10),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1537),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1539),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1646),
.B(n_469),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1568),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_1720)
);

AO21x1_ASAP7_75t_L g1721 ( 
.A1(n_1529),
.A2(n_11),
.B(n_12),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1538),
.A2(n_1027),
.B(n_1018),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1545),
.B(n_470),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1532),
.A2(n_1027),
.B(n_1018),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1652),
.A2(n_16),
.B(n_13),
.C(n_14),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1542),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1534),
.B(n_904),
.Y(n_1727)
);

INVx3_ASAP7_75t_SL g1728 ( 
.A(n_1543),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1548),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1555),
.B(n_16),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1579),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_SL g1732 ( 
.A(n_1544),
.B(n_904),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1597),
.B(n_17),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1540),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1541),
.B(n_471),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1584),
.B(n_472),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1527),
.B(n_1635),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1547),
.B(n_1549),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1672),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1587),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1602),
.A2(n_935),
.B1(n_939),
.B2(n_936),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1531),
.B(n_935),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1550),
.A2(n_1027),
.B(n_1018),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1656),
.B(n_18),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1596),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1565),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1660),
.A2(n_904),
.B(n_20),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1586),
.B(n_473),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1589),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_SL g1750 ( 
.A(n_1551),
.B(n_939),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_SL g1751 ( 
.A1(n_1561),
.A2(n_24),
.B(n_21),
.C(n_23),
.Y(n_1751)
);

NOR2xp67_ASAP7_75t_L g1752 ( 
.A(n_1546),
.B(n_474),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1670),
.B(n_23),
.Y(n_1753)
);

AND2x6_ASAP7_75t_L g1754 ( 
.A(n_1645),
.B(n_1677),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_SL g1755 ( 
.A1(n_1661),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1755)
);

BUFx8_ASAP7_75t_L g1756 ( 
.A(n_1576),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1580),
.B(n_475),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1571),
.A2(n_1027),
.B(n_943),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1561),
.B(n_939),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1578),
.B(n_476),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1577),
.B(n_26),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1659),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1562),
.A2(n_954),
.B(n_943),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1588),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1647),
.B(n_27),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1659),
.B(n_944),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1573),
.B(n_1574),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1591),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1594),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1769)
);

O2A1O1Ixp5_ASAP7_75t_L g1770 ( 
.A1(n_1636),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1677),
.B(n_944),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1613),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1526),
.Y(n_1773)
);

AOI22x1_ASAP7_75t_SL g1774 ( 
.A1(n_1642),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1614),
.B(n_949),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1592),
.B(n_478),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1616),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1575),
.B(n_31),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1675),
.A2(n_950),
.B1(n_954),
.B2(n_949),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1676),
.A2(n_954),
.B(n_950),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1556),
.B(n_32),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1601),
.B(n_33),
.Y(n_1782)
);

INVx3_ASAP7_75t_SL g1783 ( 
.A(n_1609),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1676),
.A2(n_954),
.B(n_950),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1633),
.B(n_35),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1667),
.B(n_35),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1673),
.Y(n_1787)
);

NOR2xp67_ASAP7_75t_L g1788 ( 
.A(n_1604),
.B(n_480),
.Y(n_1788)
);

OR2x6_ASAP7_75t_SL g1789 ( 
.A(n_1566),
.B(n_36),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1526),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1679),
.A2(n_584),
.B(n_483),
.Y(n_1791)
);

OAI21xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1637),
.A2(n_484),
.B(n_481),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1663),
.B(n_1669),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1618),
.B(n_1623),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1608),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_L g1796 ( 
.A1(n_1599),
.A2(n_36),
.B(n_37),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1644),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1634),
.B(n_38),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1639),
.B(n_39),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1572),
.B(n_485),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1569),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1638),
.B(n_486),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_1569),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1679),
.A2(n_583),
.B(n_490),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1610),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1569),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1585),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1582),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1685),
.B(n_1611),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1612),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1810)
);

CKINVDCx8_ASAP7_75t_R g1811 ( 
.A(n_1585),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1558),
.A2(n_582),
.B(n_491),
.Y(n_1812)
);

NAND2xp33_ASAP7_75t_SL g1813 ( 
.A(n_1671),
.B(n_47),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1674),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1620),
.B(n_487),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1560),
.A2(n_581),
.B(n_494),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1671),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1657),
.A2(n_580),
.B(n_495),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1622),
.B(n_493),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1682),
.B(n_52),
.C(n_53),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1662),
.B(n_1572),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1643),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1657),
.A2(n_579),
.B(n_496),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1585),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1681),
.B(n_55),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1624),
.B(n_1625),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1648),
.A2(n_500),
.B(n_498),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1632),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1678),
.B(n_56),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1649),
.A2(n_504),
.B(n_503),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1590),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1626),
.B(n_58),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1630),
.B(n_59),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1683),
.B(n_59),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1665),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1553),
.A2(n_578),
.B(n_509),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1583),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1583),
.B(n_63),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_SL g1839 ( 
.A1(n_1721),
.A2(n_1684),
.B(n_1629),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1691),
.A2(n_1564),
.B(n_1552),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1708),
.A2(n_1570),
.B1(n_1567),
.B2(n_1619),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1711),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1809),
.B(n_1662),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1688),
.A2(n_1658),
.B(n_1581),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1694),
.B(n_1619),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1767),
.B(n_1664),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1701),
.A2(n_1563),
.B(n_1664),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1826),
.B(n_1671),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1687),
.A2(n_1590),
.B(n_1666),
.Y(n_1849)
);

AO31x2_ASAP7_75t_L g1850 ( 
.A1(n_1703),
.A2(n_1666),
.A3(n_1590),
.B(n_1621),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1717),
.B(n_64),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1697),
.A2(n_510),
.B(n_505),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1699),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1689),
.B(n_64),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1757),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1726),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1747),
.A2(n_66),
.B(n_68),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1764),
.Y(n_1858)
);

INVx5_ASAP7_75t_L g1859 ( 
.A(n_1742),
.Y(n_1859)
);

NAND3xp33_ASAP7_75t_L g1860 ( 
.A(n_1820),
.B(n_69),
.C(n_70),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1698),
.A2(n_1784),
.B(n_1780),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1821),
.B(n_511),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1700),
.A2(n_514),
.B(n_512),
.Y(n_1863)
);

AOI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1775),
.A2(n_516),
.B(n_515),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1716),
.B(n_69),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1692),
.A2(n_518),
.B(n_517),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1786),
.A2(n_70),
.B(n_71),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1722),
.A2(n_521),
.B(n_519),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1723),
.A2(n_72),
.B(n_73),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1706),
.A2(n_75),
.B(n_72),
.C(n_74),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1754),
.B(n_74),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_SL g1872 ( 
.A(n_1771),
.B(n_523),
.Y(n_1872)
);

OAI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1724),
.A2(n_526),
.B(n_525),
.Y(n_1873)
);

NAND2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1696),
.B(n_528),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1772),
.Y(n_1875)
);

AOI21x1_ASAP7_75t_SL g1876 ( 
.A1(n_1733),
.A2(n_1765),
.B(n_1753),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1735),
.A2(n_75),
.B(n_76),
.Y(n_1877)
);

BUFx2_ASAP7_75t_SL g1878 ( 
.A(n_1803),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1791),
.A2(n_1804),
.B(n_1818),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1729),
.B(n_78),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1713),
.B(n_532),
.Y(n_1881)
);

AO31x2_ASAP7_75t_L g1882 ( 
.A1(n_1709),
.A2(n_534),
.A3(n_535),
.B(n_533),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1754),
.B(n_79),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1754),
.B(n_79),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1731),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1756),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1740),
.Y(n_1887)
);

AOI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1704),
.A2(n_538),
.B(n_537),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1749),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1802),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1793),
.A2(n_81),
.B(n_82),
.Y(n_1891)
);

O2A1O1Ixp5_ASAP7_75t_L g1892 ( 
.A1(n_1823),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1808),
.A2(n_85),
.B(n_87),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1768),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1758),
.A2(n_540),
.B(n_539),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1739),
.A2(n_88),
.B(n_89),
.Y(n_1896)
);

A2O1A1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1796),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1835),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1760),
.B(n_543),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1686),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1827),
.A2(n_545),
.B(n_544),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1763),
.A2(n_1771),
.B(n_1759),
.Y(n_1902)
);

OAI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1830),
.A2(n_547),
.B(n_546),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1743),
.A2(n_549),
.B(n_548),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1815),
.A2(n_91),
.B(n_92),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1707),
.B(n_550),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1736),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1812),
.A2(n_552),
.B(n_551),
.Y(n_1908)
);

AO21x2_ASAP7_75t_L g1909 ( 
.A1(n_1816),
.A2(n_93),
.B(n_95),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1795),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1718),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1713),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1836),
.A2(n_554),
.B(n_553),
.Y(n_1913)
);

AND2x4_ASAP7_75t_SL g1914 ( 
.A(n_1762),
.B(n_555),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1754),
.B(n_96),
.Y(n_1915)
);

OAI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1738),
.A2(n_558),
.B(n_556),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1819),
.A2(n_96),
.B(n_97),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1822),
.A2(n_562),
.B(n_561),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1696),
.B(n_564),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1762),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1769),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1817),
.Y(n_1922)
);

BUFx3_ASAP7_75t_L g1923 ( 
.A(n_1745),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1737),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1817),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1777),
.B(n_568),
.Y(n_1926)
);

AOI211x1_ASAP7_75t_L g1927 ( 
.A1(n_1797),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_L g1928 ( 
.A(n_1783),
.B(n_1744),
.Y(n_1928)
);

NAND2x1p5_ASAP7_75t_L g1929 ( 
.A(n_1696),
.B(n_1790),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1734),
.B(n_102),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1828),
.A2(n_105),
.B(n_108),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1712),
.B(n_1750),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1811),
.B(n_570),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1751),
.A2(n_574),
.B(n_573),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1779),
.A2(n_576),
.B(n_575),
.Y(n_1935)
);

OAI21x1_ASAP7_75t_L g1936 ( 
.A1(n_1770),
.A2(n_108),
.B(n_109),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1693),
.A2(n_109),
.B(n_111),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1710),
.B(n_451),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1794),
.A2(n_112),
.B(n_113),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1801),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1773),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1800),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1761),
.A2(n_112),
.B(n_113),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1785),
.A2(n_114),
.B(n_115),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1728),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1778),
.B(n_116),
.Y(n_1946)
);

OA21x2_ASAP7_75t_L g1947 ( 
.A1(n_1814),
.A2(n_117),
.B(n_118),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1781),
.B(n_1787),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_L g1949 ( 
.A1(n_1798),
.A2(n_118),
.B(n_119),
.Y(n_1949)
);

NAND2x1p5_ASAP7_75t_L g1950 ( 
.A(n_1859),
.B(n_1806),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1853),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1948),
.B(n_1690),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1869),
.B(n_1752),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1912),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1853),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1846),
.B(n_1715),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1920),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1875),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1856),
.B(n_1742),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1856),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1940),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1879),
.A2(n_1755),
.B(n_1788),
.Y(n_1962)
);

CKINVDCx6p67_ASAP7_75t_R g1963 ( 
.A(n_1878),
.Y(n_1963)
);

BUFx4f_ASAP7_75t_L g1964 ( 
.A(n_1926),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1858),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1885),
.B(n_1773),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1921),
.A2(n_1805),
.B1(n_1810),
.B2(n_1746),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1885),
.B(n_1773),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1893),
.A2(n_1855),
.B1(n_1932),
.B2(n_1877),
.Y(n_1969)
);

OR2x6_ASAP7_75t_L g1970 ( 
.A(n_1843),
.B(n_1849),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1887),
.B(n_1807),
.Y(n_1971)
);

NAND2x1p5_ASAP7_75t_L g1972 ( 
.A(n_1859),
.B(n_1800),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1887),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1923),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1889),
.B(n_1705),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1889),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1941),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1870),
.A2(n_1931),
.B1(n_1890),
.B2(n_1897),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1905),
.B(n_1725),
.C(n_1720),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1848),
.B(n_1834),
.Y(n_1980)
);

AOI21xp33_ASAP7_75t_SL g1981 ( 
.A1(n_1886),
.A2(n_1695),
.B(n_1782),
.Y(n_1981)
);

AO21x2_ASAP7_75t_L g1982 ( 
.A1(n_1847),
.A2(n_1829),
.B(n_1714),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1917),
.B(n_1776),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1841),
.B(n_1748),
.Y(n_1984)
);

BUFx3_ASAP7_75t_L g1985 ( 
.A(n_1898),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1842),
.B(n_1911),
.Y(n_1986)
);

NOR2x1_ASAP7_75t_SL g1987 ( 
.A(n_1909),
.B(n_1766),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1894),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1926),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1928),
.A2(n_1813),
.B1(n_1833),
.B2(n_1832),
.Y(n_1990)
);

O2A1O1Ixp33_ASAP7_75t_SL g1991 ( 
.A1(n_1907),
.A2(n_1837),
.B(n_1702),
.C(n_1730),
.Y(n_1991)
);

NAND2x1_ASAP7_75t_L g1992 ( 
.A(n_1894),
.B(n_1766),
.Y(n_1992)
);

AO21x1_ASAP7_75t_L g1993 ( 
.A1(n_1891),
.A2(n_1838),
.B(n_1825),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1941),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1910),
.B(n_1789),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1910),
.B(n_1799),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1845),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1854),
.B(n_1719),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1922),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1906),
.B(n_1774),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1865),
.B(n_1807),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1922),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1939),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1942),
.B(n_1946),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1882),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1938),
.A2(n_1741),
.B1(n_1824),
.B2(n_1807),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1930),
.B(n_1880),
.Y(n_2007)
);

BUFx12f_ASAP7_75t_L g2008 ( 
.A(n_1881),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1857),
.A2(n_1756),
.B1(n_1792),
.B2(n_1824),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1925),
.Y(n_2010)
);

INVx5_ASAP7_75t_L g2011 ( 
.A(n_1862),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1859),
.B(n_1824),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1860),
.A2(n_1831),
.B1(n_1727),
.B2(n_1732),
.Y(n_2013)
);

AOI222xp33_ASAP7_75t_L g2014 ( 
.A1(n_1867),
.A2(n_123),
.B1(n_125),
.B2(n_120),
.C1(n_121),
.C2(n_124),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1943),
.B(n_1831),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1937),
.Y(n_2016)
);

AO21x2_ASAP7_75t_L g2017 ( 
.A1(n_1844),
.A2(n_1831),
.B(n_120),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1882),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1925),
.Y(n_2019)
);

A2O1A1Ixp33_ASAP7_75t_SL g2020 ( 
.A1(n_1944),
.A2(n_1896),
.B(n_1924),
.C(n_1900),
.Y(n_2020)
);

INVx5_ASAP7_75t_L g2021 ( 
.A(n_1862),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1850),
.B(n_123),
.Y(n_2022)
);

OAI321xp33_ASAP7_75t_L g2023 ( 
.A1(n_1945),
.A2(n_126),
.A3(n_127),
.B1(n_128),
.B2(n_130),
.C(n_131),
.Y(n_2023)
);

BUFx4_ASAP7_75t_SL g2024 ( 
.A(n_1958),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_1954),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1951),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1951),
.Y(n_2027)
);

INVx6_ASAP7_75t_L g2028 ( 
.A(n_1961),
.Y(n_2028)
);

INVx6_ASAP7_75t_L g2029 ( 
.A(n_1961),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1963),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1955),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1967),
.A2(n_1969),
.B1(n_1978),
.B2(n_1979),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1983),
.A2(n_1927),
.B1(n_1947),
.B2(n_1871),
.Y(n_2033)
);

OAI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_2011),
.A2(n_1883),
.B1(n_1915),
.B2(n_1884),
.Y(n_2034)
);

CKINVDCx8_ASAP7_75t_R g2035 ( 
.A(n_1961),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1955),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_1965),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_SL g2038 ( 
.A1(n_1995),
.A2(n_1947),
.B1(n_1861),
.B2(n_1902),
.Y(n_2038)
);

INVx6_ASAP7_75t_L g2039 ( 
.A(n_1985),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1988),
.Y(n_2040)
);

INVx1_ASAP7_75t_SL g2041 ( 
.A(n_1954),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1974),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_2014),
.A2(n_1899),
.B1(n_1909),
.B2(n_1839),
.Y(n_2043)
);

CKINVDCx11_ASAP7_75t_R g2044 ( 
.A(n_2008),
.Y(n_2044)
);

BUFx12f_ASAP7_75t_L g2045 ( 
.A(n_1989),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1953),
.A2(n_1933),
.B1(n_1934),
.B2(n_1851),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1960),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_1964),
.A2(n_1927),
.B1(n_1863),
.B2(n_1904),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1973),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1976),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1957),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_1994),
.Y(n_2052)
);

CKINVDCx20_ASAP7_75t_R g2053 ( 
.A(n_1952),
.Y(n_2053)
);

NAND2x1p5_ASAP7_75t_L g2054 ( 
.A(n_2011),
.B(n_1866),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1997),
.Y(n_2055)
);

INVx4_ASAP7_75t_L g2056 ( 
.A(n_2012),
.Y(n_2056)
);

CKINVDCx11_ASAP7_75t_R g2057 ( 
.A(n_1994),
.Y(n_2057)
);

BUFx12f_ASAP7_75t_L g2058 ( 
.A(n_1989),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1964),
.A2(n_1874),
.B1(n_1919),
.B2(n_1935),
.Y(n_2059)
);

INVx6_ASAP7_75t_L g2060 ( 
.A(n_1994),
.Y(n_2060)
);

AOI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_1984),
.A2(n_1949),
.B1(n_1936),
.B2(n_1918),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1993),
.A2(n_1881),
.B1(n_1840),
.B2(n_1901),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_1957),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1970),
.A2(n_1903),
.B1(n_1908),
.B2(n_1913),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1966),
.Y(n_2065)
);

CKINVDCx6p67_ASAP7_75t_R g2066 ( 
.A(n_2001),
.Y(n_2066)
);

INVxp67_ASAP7_75t_SL g2067 ( 
.A(n_2010),
.Y(n_2067)
);

INVx4_ASAP7_75t_L g2068 ( 
.A(n_2012),
.Y(n_2068)
);

INVx6_ASAP7_75t_L g2069 ( 
.A(n_1989),
.Y(n_2069)
);

BUFx10_ASAP7_75t_L g2070 ( 
.A(n_2022),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1986),
.Y(n_2071)
);

BUFx12f_ASAP7_75t_L g2072 ( 
.A(n_2007),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2055),
.B(n_2071),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2047),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_2032),
.A2(n_1962),
.B(n_2020),
.Y(n_2075)
);

BUFx8_ASAP7_75t_L g2076 ( 
.A(n_2037),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2067),
.B(n_2050),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_SL g2078 ( 
.A1(n_2032),
.A2(n_1987),
.B(n_1970),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2026),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_2028),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_2048),
.A2(n_1991),
.B(n_1892),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_2048),
.A2(n_1987),
.B(n_1982),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2025),
.B(n_1956),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_2025),
.Y(n_2084)
);

AOI31xp33_ASAP7_75t_L g2085 ( 
.A1(n_2030),
.A2(n_1981),
.A3(n_1972),
.B(n_1998),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_2028),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2043),
.A2(n_2009),
.B1(n_1990),
.B2(n_2011),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2027),
.Y(n_2088)
);

O2A1O1Ixp5_ASAP7_75t_L g2089 ( 
.A1(n_2033),
.A2(n_1992),
.B(n_2016),
.C(n_2022),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2041),
.B(n_2005),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2041),
.B(n_2005),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2031),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2051),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2063),
.B(n_2018),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2046),
.A2(n_2021),
.B1(n_2015),
.B2(n_2013),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2049),
.B(n_2018),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2046),
.A2(n_2021),
.B1(n_1980),
.B2(n_2000),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2040),
.B(n_2003),
.Y(n_2098)
);

NOR2xp67_ASAP7_75t_L g2099 ( 
.A(n_2063),
.B(n_2021),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2079),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2075),
.A2(n_2062),
.B1(n_2033),
.B2(n_2061),
.Y(n_2101)
);

NOR3xp33_ASAP7_75t_SL g2102 ( 
.A(n_2097),
.B(n_2034),
.C(n_2023),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_R g2103 ( 
.A(n_2076),
.B(n_2044),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2098),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2085),
.B(n_2053),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_R g2106 ( 
.A(n_2076),
.B(n_2035),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2083),
.B(n_2065),
.Y(n_2107)
);

NOR2x1p5_ASAP7_75t_L g2108 ( 
.A(n_2080),
.B(n_2072),
.Y(n_2108)
);

AO31x2_ASAP7_75t_L g2109 ( 
.A1(n_2082),
.A2(n_2036),
.A3(n_2068),
.B(n_2056),
.Y(n_2109)
);

NAND3xp33_ASAP7_75t_L g2110 ( 
.A(n_2081),
.B(n_2038),
.C(n_2061),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2084),
.B(n_2093),
.Y(n_2111)
);

AO21x2_ASAP7_75t_L g2112 ( 
.A1(n_2110),
.A2(n_2078),
.B(n_2099),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_2110),
.Y(n_2113)
);

AOI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2101),
.A2(n_2087),
.B1(n_2078),
.B2(n_2089),
.C(n_2095),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2100),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_2108),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2111),
.B(n_2080),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2104),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2109),
.B(n_2086),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2115),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2112),
.B(n_2109),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2113),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2112),
.B(n_2109),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2113),
.Y(n_2124)
);

AOI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_2113),
.A2(n_2105),
.B1(n_2066),
.B2(n_2059),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2112),
.B(n_2086),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2118),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2113),
.B(n_2102),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2116),
.B(n_2090),
.Y(n_2129)
);

AOI21xp5_ASAP7_75t_L g2130 ( 
.A1(n_2128),
.A2(n_2113),
.B(n_2114),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2124),
.Y(n_2131)
);

NAND2xp33_ASAP7_75t_SL g2132 ( 
.A(n_2124),
.B(n_2113),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2129),
.B(n_2116),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2129),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_SL g2135 ( 
.A1(n_2122),
.A2(n_2103),
.B1(n_2039),
.B2(n_2024),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2126),
.B(n_2117),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2127),
.Y(n_2137)
);

INVxp67_ASAP7_75t_L g2138 ( 
.A(n_2120),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2127),
.Y(n_2139)
);

AOI221xp5_ASAP7_75t_L g2140 ( 
.A1(n_2120),
.A2(n_2114),
.B1(n_2118),
.B2(n_2119),
.C(n_2117),
.Y(n_2140)
);

OAI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2125),
.A2(n_2119),
.B1(n_2038),
.B2(n_2099),
.C(n_2073),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2136),
.B(n_2126),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_2135),
.B(n_2130),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2133),
.B(n_2106),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2131),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2134),
.B(n_2121),
.Y(n_2146)
);

OR2x2_ASAP7_75t_SL g2147 ( 
.A(n_2131),
.B(n_2039),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2137),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2138),
.B(n_2121),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2138),
.B(n_2132),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2145),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2150),
.B(n_2142),
.Y(n_2152)
);

NAND2x1_ASAP7_75t_L g2153 ( 
.A(n_2144),
.B(n_2123),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2143),
.B(n_2140),
.Y(n_2154)
);

NAND2x1p5_ASAP7_75t_L g2155 ( 
.A(n_2153),
.B(n_2143),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_2152),
.B(n_2147),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_2154),
.B(n_2141),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2151),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2156),
.B(n_2155),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2157),
.B(n_2146),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2158),
.Y(n_2161)
);

INVxp67_ASAP7_75t_L g2162 ( 
.A(n_2156),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2155),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2155),
.Y(n_2164)
);

INVx1_ASAP7_75t_SL g2165 ( 
.A(n_2159),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2162),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2163),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2163),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2164),
.B(n_2132),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2162),
.B(n_2149),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2160),
.Y(n_2171)
);

INVxp67_ASAP7_75t_L g2172 ( 
.A(n_2161),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2163),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2162),
.B(n_2149),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2165),
.B(n_2148),
.Y(n_2175)
);

AOI211x1_ASAP7_75t_SL g2176 ( 
.A1(n_2169),
.A2(n_2139),
.B(n_2123),
.C(n_2006),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2165),
.B(n_2042),
.Y(n_2177)
);

OAI22xp33_ASAP7_75t_L g2178 ( 
.A1(n_2171),
.A2(n_2029),
.B1(n_2074),
.B2(n_2077),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2167),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2166),
.B(n_2107),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2168),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2173),
.B(n_2076),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_2170),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2174),
.A2(n_2029),
.B1(n_2058),
.B2(n_2045),
.Y(n_2184)
);

AOI322xp5_ASAP7_75t_L g2185 ( 
.A1(n_2172),
.A2(n_2091),
.A3(n_2090),
.B1(n_2094),
.B2(n_2004),
.C1(n_2064),
.C2(n_2003),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2167),
.Y(n_2186)
);

AOI31xp33_ASAP7_75t_L g2187 ( 
.A1(n_2165),
.A2(n_1929),
.A3(n_1950),
.B(n_1975),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2179),
.B(n_2098),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2186),
.B(n_2079),
.Y(n_2189)
);

NAND3xp33_ASAP7_75t_L g2190 ( 
.A(n_2177),
.B(n_2057),
.C(n_126),
.Y(n_2190)
);

A2O1A1Ixp33_ASAP7_75t_L g2191 ( 
.A1(n_2183),
.A2(n_2181),
.B(n_2182),
.C(n_2175),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_2180),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2176),
.Y(n_2193)
);

OAI21xp33_ASAP7_75t_L g2194 ( 
.A1(n_2187),
.A2(n_2184),
.B(n_2178),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2185),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2179),
.B(n_2088),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2177),
.Y(n_2197)
);

OAI221xp5_ASAP7_75t_L g2198 ( 
.A1(n_2182),
.A2(n_2059),
.B1(n_2054),
.B2(n_1996),
.C(n_2069),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2179),
.B(n_2088),
.Y(n_2199)
);

AOI21xp33_ASAP7_75t_L g2200 ( 
.A1(n_2182),
.A2(n_127),
.B(n_128),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2179),
.Y(n_2201)
);

INVx1_ASAP7_75t_SL g2202 ( 
.A(n_2177),
.Y(n_2202)
);

NAND2xp33_ASAP7_75t_R g2203 ( 
.A(n_2197),
.B(n_131),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2201),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2202),
.B(n_2092),
.Y(n_2205)
);

CKINVDCx16_ASAP7_75t_R g2206 ( 
.A(n_2193),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2190),
.B(n_132),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2195),
.A2(n_2060),
.B1(n_2017),
.B2(n_2069),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2188),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2192),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2189),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2191),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_2200),
.B(n_132),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2194),
.B(n_2092),
.Y(n_2214)
);

NOR2x1_ASAP7_75t_L g2215 ( 
.A(n_2196),
.B(n_133),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2199),
.B(n_2091),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2215),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_2204),
.B(n_2198),
.Y(n_2218)
);

OAI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2208),
.A2(n_2060),
.B1(n_2052),
.B2(n_2056),
.Y(n_2219)
);

AND3x1_ASAP7_75t_L g2220 ( 
.A(n_2213),
.B(n_133),
.C(n_134),
.Y(n_2220)
);

NAND3xp33_ASAP7_75t_L g2221 ( 
.A(n_2203),
.B(n_134),
.C(n_135),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2207),
.Y(n_2222)
);

NOR2x1_ASAP7_75t_L g2223 ( 
.A(n_2212),
.B(n_135),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_2209),
.B(n_2070),
.Y(n_2224)
);

NOR3xp33_ASAP7_75t_L g2225 ( 
.A(n_2210),
.B(n_1876),
.C(n_136),
.Y(n_2225)
);

NOR3xp33_ASAP7_75t_L g2226 ( 
.A(n_2206),
.B(n_136),
.C(n_137),
.Y(n_2226)
);

AND4x1_ASAP7_75t_L g2227 ( 
.A(n_2214),
.B(n_139),
.C(n_137),
.D(n_138),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2205),
.A2(n_1872),
.B(n_1914),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2211),
.Y(n_2229)
);

NAND4xp75_ASAP7_75t_L g2230 ( 
.A(n_2216),
.B(n_141),
.C(n_138),
.D(n_140),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2207),
.B(n_140),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2212),
.B(n_141),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2212),
.B(n_142),
.Y(n_2233)
);

NAND4xp25_ASAP7_75t_SL g2234 ( 
.A(n_2208),
.B(n_2094),
.C(n_2096),
.D(n_144),
.Y(n_2234)
);

AOI211xp5_ASAP7_75t_SL g2235 ( 
.A1(n_2212),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2235)
);

NAND2xp33_ASAP7_75t_L g2236 ( 
.A(n_2215),
.B(n_143),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2212),
.B(n_145),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2212),
.B(n_145),
.Y(n_2238)
);

AOI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2236),
.A2(n_146),
.B(n_147),
.Y(n_2239)
);

O2A1O1Ixp33_ASAP7_75t_L g2240 ( 
.A1(n_2217),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2227),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2235),
.B(n_2070),
.Y(n_2242)
);

NAND4xp25_ASAP7_75t_L g2243 ( 
.A(n_2218),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2221),
.B(n_149),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2226),
.B(n_150),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2220),
.A2(n_1977),
.B1(n_2068),
.B2(n_2096),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_2230),
.Y(n_2247)
);

AND4x1_ASAP7_75t_L g2248 ( 
.A(n_2231),
.B(n_153),
.C(n_151),
.D(n_152),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_SL g2249 ( 
.A(n_2223),
.B(n_152),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2222),
.B(n_153),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2229),
.B(n_154),
.Y(n_2251)
);

NAND3xp33_ASAP7_75t_L g2252 ( 
.A(n_2232),
.B(n_154),
.C(n_155),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2233),
.Y(n_2253)
);

NOR2xp67_ASAP7_75t_L g2254 ( 
.A(n_2234),
.B(n_2237),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2224),
.B(n_156),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2238),
.Y(n_2256)
);

AOI211xp5_ASAP7_75t_SL g2257 ( 
.A1(n_2225),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_2257)
);

NAND3xp33_ASAP7_75t_SL g2258 ( 
.A(n_2228),
.B(n_157),
.C(n_158),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_2219),
.Y(n_2259)
);

O2A1O1Ixp33_ASAP7_75t_L g2260 ( 
.A1(n_2236),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2260)
);

NOR2x1_ASAP7_75t_SL g2261 ( 
.A(n_2230),
.B(n_1864),
.Y(n_2261)
);

NAND5xp2_ASAP7_75t_L g2262 ( 
.A(n_2229),
.B(n_161),
.C(n_159),
.D(n_160),
.E(n_162),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2217),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2223),
.B(n_162),
.C(n_163),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2217),
.Y(n_2265)
);

OAI221xp5_ASAP7_75t_L g2266 ( 
.A1(n_2225),
.A2(n_166),
.B1(n_163),
.B2(n_165),
.C(n_167),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2230),
.Y(n_2267)
);

NAND2x1p5_ASAP7_75t_L g2268 ( 
.A(n_2217),
.B(n_1916),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2217),
.Y(n_2269)
);

INVx1_ASAP7_75t_SL g2270 ( 
.A(n_2230),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2235),
.B(n_165),
.Y(n_2271)
);

INVxp67_ASAP7_75t_L g2272 ( 
.A(n_2220),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_L g2273 ( 
.A(n_2223),
.B(n_166),
.C(n_167),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2235),
.B(n_168),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2217),
.Y(n_2275)
);

NAND3xp33_ASAP7_75t_L g2276 ( 
.A(n_2249),
.B(n_168),
.C(n_169),
.Y(n_2276)
);

NAND4xp75_ASAP7_75t_L g2277 ( 
.A(n_2254),
.B(n_172),
.C(n_169),
.D(n_170),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2242),
.B(n_170),
.Y(n_2278)
);

NOR3x1_ASAP7_75t_L g2279 ( 
.A(n_2243),
.B(n_172),
.C(n_173),
.Y(n_2279)
);

NAND3xp33_ASAP7_75t_SL g2280 ( 
.A(n_2260),
.B(n_173),
.C(n_174),
.Y(n_2280)
);

NAND4xp25_ASAP7_75t_L g2281 ( 
.A(n_2257),
.B(n_177),
.C(n_175),
.D(n_176),
.Y(n_2281)
);

AND4x1_ASAP7_75t_L g2282 ( 
.A(n_2264),
.B(n_181),
.C(n_179),
.D(n_180),
.Y(n_2282)
);

NAND3xp33_ASAP7_75t_SL g2283 ( 
.A(n_2247),
.B(n_182),
.C(n_183),
.Y(n_2283)
);

NOR4xp25_ASAP7_75t_L g2284 ( 
.A(n_2270),
.B(n_186),
.C(n_184),
.D(n_185),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2239),
.A2(n_185),
.B(n_186),
.Y(n_2285)
);

AOI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2266),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_2286)
);

NOR3xp33_ASAP7_75t_SL g2287 ( 
.A(n_2258),
.B(n_187),
.C(n_188),
.Y(n_2287)
);

NAND4xp25_ASAP7_75t_L g2288 ( 
.A(n_2241),
.B(n_2272),
.C(n_2267),
.D(n_2271),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2250),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2274),
.B(n_1966),
.Y(n_2290)
);

NOR3xp33_ASAP7_75t_L g2291 ( 
.A(n_2263),
.B(n_190),
.C(n_192),
.Y(n_2291)
);

NAND3xp33_ASAP7_75t_L g2292 ( 
.A(n_2264),
.B(n_193),
.C(n_194),
.Y(n_2292)
);

NOR2x1_ASAP7_75t_L g2293 ( 
.A(n_2273),
.B(n_193),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2248),
.B(n_194),
.Y(n_2294)
);

NOR4xp25_ASAP7_75t_L g2295 ( 
.A(n_2265),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_2295)
);

NAND4xp25_ASAP7_75t_L g2296 ( 
.A(n_2269),
.B(n_198),
.C(n_195),
.D(n_197),
.Y(n_2296)
);

NOR2x1_ASAP7_75t_L g2297 ( 
.A(n_2273),
.B(n_199),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2262),
.B(n_200),
.Y(n_2298)
);

NAND3xp33_ASAP7_75t_L g2299 ( 
.A(n_2244),
.B(n_200),
.C(n_201),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2275),
.B(n_201),
.Y(n_2300)
);

NAND3xp33_ASAP7_75t_SL g2301 ( 
.A(n_2255),
.B(n_202),
.C(n_203),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2259),
.A2(n_1968),
.B1(n_1971),
.B2(n_1959),
.Y(n_2302)
);

NAND3xp33_ASAP7_75t_L g2303 ( 
.A(n_2252),
.B(n_202),
.C(n_203),
.Y(n_2303)
);

AOI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_2253),
.A2(n_2256),
.B1(n_2245),
.B2(n_2251),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2240),
.A2(n_205),
.B(n_206),
.Y(n_2305)
);

NOR3xp33_ASAP7_75t_L g2306 ( 
.A(n_2246),
.B(n_205),
.C(n_207),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2268),
.A2(n_1971),
.B1(n_1968),
.B2(n_1959),
.Y(n_2307)
);

NAND4xp75_ASAP7_75t_L g2308 ( 
.A(n_2261),
.B(n_209),
.C(n_207),
.D(n_208),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_L g2309 ( 
.A(n_2272),
.B(n_208),
.C(n_209),
.Y(n_2309)
);

NAND4xp25_ASAP7_75t_L g2310 ( 
.A(n_2288),
.B(n_212),
.C(n_210),
.D(n_211),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2298),
.B(n_211),
.Y(n_2311)
);

AOI221x1_ASAP7_75t_L g2312 ( 
.A1(n_2278),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.C(n_215),
.Y(n_2312)
);

XOR2x1_ASAP7_75t_L g2313 ( 
.A(n_2289),
.B(n_213),
.Y(n_2313)
);

NOR3xp33_ASAP7_75t_L g2314 ( 
.A(n_2299),
.B(n_214),
.C(n_216),
.Y(n_2314)
);

OAI211xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2304),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2295),
.B(n_217),
.Y(n_2316)
);

NOR3xp33_ASAP7_75t_L g2317 ( 
.A(n_2301),
.B(n_218),
.C(n_219),
.Y(n_2317)
);

NOR4xp75_ASAP7_75t_L g2318 ( 
.A(n_2308),
.B(n_222),
.C(n_220),
.D(n_221),
.Y(n_2318)
);

NOR4xp75_ASAP7_75t_L g2319 ( 
.A(n_2280),
.B(n_226),
.C(n_223),
.D(n_224),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2294),
.Y(n_2320)
);

NOR3x1_ASAP7_75t_L g2321 ( 
.A(n_2281),
.B(n_226),
.C(n_227),
.Y(n_2321)
);

NOR2x1_ASAP7_75t_L g2322 ( 
.A(n_2277),
.B(n_227),
.Y(n_2322)
);

OAI211xp5_ASAP7_75t_SL g2323 ( 
.A1(n_2287),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2323)
);

AOI211xp5_ASAP7_75t_L g2324 ( 
.A1(n_2284),
.A2(n_2283),
.B(n_2292),
.C(n_2303),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2282),
.B(n_228),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2296),
.B(n_230),
.Y(n_2326)
);

NAND3xp33_ASAP7_75t_SL g2327 ( 
.A(n_2286),
.B(n_231),
.C(n_232),
.Y(n_2327)
);

NOR4xp25_ASAP7_75t_L g2328 ( 
.A(n_2276),
.B(n_234),
.C(n_232),
.D(n_233),
.Y(n_2328)
);

NOR4xp25_ASAP7_75t_L g2329 ( 
.A(n_2300),
.B(n_236),
.C(n_234),
.D(n_235),
.Y(n_2329)
);

AO21x1_ASAP7_75t_L g2330 ( 
.A1(n_2285),
.A2(n_235),
.B(n_236),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2293),
.Y(n_2331)
);

NOR4xp25_ASAP7_75t_L g2332 ( 
.A(n_2290),
.B(n_2297),
.C(n_2279),
.D(n_2306),
.Y(n_2332)
);

NOR2x1_ASAP7_75t_L g2333 ( 
.A(n_2305),
.B(n_237),
.Y(n_2333)
);

NAND3xp33_ASAP7_75t_L g2334 ( 
.A(n_2309),
.B(n_238),
.C(n_239),
.Y(n_2334)
);

NOR2x1_ASAP7_75t_L g2335 ( 
.A(n_2291),
.B(n_238),
.Y(n_2335)
);

AOI322xp5_ASAP7_75t_L g2336 ( 
.A1(n_2302),
.A2(n_2019),
.A3(n_241),
.B1(n_242),
.B2(n_243),
.C1(n_244),
.C2(n_245),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2307),
.B(n_239),
.C(n_241),
.Y(n_2337)
);

AOI211x1_ASAP7_75t_SL g2338 ( 
.A1(n_2288),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_2338)
);

NOR3xp33_ASAP7_75t_SL g2339 ( 
.A(n_2288),
.B(n_245),
.C(n_246),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2277),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2284),
.B(n_247),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2284),
.B(n_247),
.Y(n_2342)
);

AOI32xp33_ASAP7_75t_L g2343 ( 
.A1(n_2293),
.A2(n_248),
.A3(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_SL g2344 ( 
.A(n_2284),
.B(n_248),
.C(n_249),
.Y(n_2344)
);

NOR3xp33_ASAP7_75t_L g2345 ( 
.A(n_2288),
.B(n_250),
.C(n_251),
.Y(n_2345)
);

AOI211xp5_ASAP7_75t_L g2346 ( 
.A1(n_2284),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_2346)
);

NOR4xp25_ASAP7_75t_L g2347 ( 
.A(n_2288),
.B(n_256),
.C(n_252),
.D(n_255),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2278),
.A2(n_255),
.B(n_256),
.Y(n_2348)
);

NAND4xp25_ASAP7_75t_L g2349 ( 
.A(n_2288),
.B(n_259),
.C(n_257),
.D(n_258),
.Y(n_2349)
);

AOI21xp33_ASAP7_75t_L g2350 ( 
.A1(n_2278),
.A2(n_258),
.B(n_260),
.Y(n_2350)
);

NOR4xp25_ASAP7_75t_L g2351 ( 
.A(n_2288),
.B(n_262),
.C(n_260),
.D(n_261),
.Y(n_2351)
);

NOR3xp33_ASAP7_75t_L g2352 ( 
.A(n_2288),
.B(n_261),
.C(n_262),
.Y(n_2352)
);

NOR2x1_ASAP7_75t_L g2353 ( 
.A(n_2277),
.B(n_263),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2298),
.B(n_263),
.Y(n_2354)
);

NAND3xp33_ASAP7_75t_L g2355 ( 
.A(n_2282),
.B(n_264),
.C(n_265),
.Y(n_2355)
);

OAI211xp5_ASAP7_75t_SL g2356 ( 
.A1(n_2304),
.A2(n_267),
.B(n_264),
.C(n_265),
.Y(n_2356)
);

NOR3xp33_ASAP7_75t_L g2357 ( 
.A(n_2288),
.B(n_267),
.C(n_268),
.Y(n_2357)
);

AOI211x1_ASAP7_75t_L g2358 ( 
.A1(n_2305),
.A2(n_1888),
.B(n_271),
.C(n_269),
.Y(n_2358)
);

NOR2x1_ASAP7_75t_L g2359 ( 
.A(n_2277),
.B(n_270),
.Y(n_2359)
);

NAND3xp33_ASAP7_75t_SL g2360 ( 
.A(n_2284),
.B(n_270),
.C(n_271),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2298),
.B(n_272),
.Y(n_2361)
);

AOI22xp33_ASAP7_75t_L g2362 ( 
.A1(n_2317),
.A2(n_2002),
.B1(n_1999),
.B2(n_1868),
.Y(n_2362)
);

A2O1A1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2343),
.A2(n_2326),
.B(n_2348),
.C(n_2336),
.Y(n_2363)
);

NAND5xp2_ASAP7_75t_L g2364 ( 
.A(n_2324),
.B(n_273),
.C(n_274),
.D(n_275),
.E(n_276),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2345),
.B(n_2357),
.C(n_2352),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_R g2366 ( 
.A(n_2344),
.B(n_273),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2313),
.Y(n_2367)
);

AOI221xp5_ASAP7_75t_L g2368 ( 
.A1(n_2347),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.C(n_277),
.Y(n_2368)
);

INVx1_ASAP7_75t_SL g2369 ( 
.A(n_2318),
.Y(n_2369)
);

AOI222xp33_ASAP7_75t_L g2370 ( 
.A1(n_2360),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.C1(n_281),
.C2(n_282),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2329),
.B(n_279),
.Y(n_2371)
);

OAI322xp33_ASAP7_75t_L g2372 ( 
.A1(n_2340),
.A2(n_280),
.A3(n_281),
.B1(n_283),
.B2(n_285),
.C1(n_286),
.C2(n_288),
.Y(n_2372)
);

OAI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2355),
.A2(n_2353),
.B(n_2322),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2351),
.B(n_283),
.Y(n_2374)
);

NOR2x1_ASAP7_75t_L g2375 ( 
.A(n_2310),
.B(n_286),
.Y(n_2375)
);

INVx1_ASAP7_75t_SL g2376 ( 
.A(n_2319),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2316),
.Y(n_2377)
);

OAI211xp5_ASAP7_75t_L g2378 ( 
.A1(n_2328),
.A2(n_288),
.B(n_289),
.C(n_290),
.Y(n_2378)
);

NOR3xp33_ASAP7_75t_L g2379 ( 
.A(n_2361),
.B(n_289),
.C(n_290),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2341),
.A2(n_291),
.B(n_293),
.Y(n_2380)
);

OAI211xp5_ASAP7_75t_SL g2381 ( 
.A1(n_2340),
.A2(n_293),
.B(n_294),
.C(n_295),
.Y(n_2381)
);

INVx1_ASAP7_75t_SL g2382 ( 
.A(n_2325),
.Y(n_2382)
);

O2A1O1Ixp33_ASAP7_75t_L g2383 ( 
.A1(n_2342),
.A2(n_295),
.B(n_296),
.C(n_297),
.Y(n_2383)
);

OAI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_2349),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_2384)
);

OAI311xp33_ASAP7_75t_L g2385 ( 
.A1(n_2331),
.A2(n_298),
.A3(n_299),
.B1(n_300),
.C1(n_301),
.Y(n_2385)
);

OAI21xp33_ASAP7_75t_SL g2386 ( 
.A1(n_2359),
.A2(n_300),
.B(n_301),
.Y(n_2386)
);

O2A1O1Ixp33_ASAP7_75t_L g2387 ( 
.A1(n_2311),
.A2(n_302),
.B(n_304),
.C(n_305),
.Y(n_2387)
);

OAI32xp33_ASAP7_75t_L g2388 ( 
.A1(n_2338),
.A2(n_302),
.A3(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2330),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2354),
.Y(n_2390)
);

OAI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2346),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2333),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2339),
.B(n_2332),
.Y(n_2393)
);

AOI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_2327),
.A2(n_308),
.B(n_309),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2312),
.B(n_310),
.Y(n_2395)
);

BUFx2_ASAP7_75t_L g2396 ( 
.A(n_2335),
.Y(n_2396)
);

OAI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2334),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_2397)
);

INVx1_ASAP7_75t_SL g2398 ( 
.A(n_2350),
.Y(n_2398)
);

NOR2x1p5_ASAP7_75t_L g2399 ( 
.A(n_2337),
.B(n_311),
.Y(n_2399)
);

XOR2x2_ASAP7_75t_L g2400 ( 
.A(n_2314),
.B(n_312),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_2320),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_2323),
.B(n_314),
.Y(n_2402)
);

CKINVDCx20_ASAP7_75t_R g2403 ( 
.A(n_2321),
.Y(n_2403)
);

NAND4xp25_ASAP7_75t_L g2404 ( 
.A(n_2315),
.B(n_2356),
.C(n_2358),
.D(n_317),
.Y(n_2404)
);

AOI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_2341),
.A2(n_315),
.B(n_316),
.Y(n_2405)
);

CKINVDCx20_ASAP7_75t_R g2406 ( 
.A(n_2339),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2339),
.B(n_315),
.Y(n_2407)
);

NAND2xp33_ASAP7_75t_SL g2408 ( 
.A(n_2339),
.B(n_318),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2310),
.B(n_319),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2313),
.B(n_319),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2407),
.B(n_320),
.Y(n_2411)
);

XNOR2xp5_ASAP7_75t_L g2412 ( 
.A(n_2406),
.B(n_321),
.Y(n_2412)
);

XNOR2xp5_ASAP7_75t_L g2413 ( 
.A(n_2400),
.B(n_321),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2373),
.B(n_322),
.Y(n_2414)
);

AOI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2408),
.A2(n_1873),
.B1(n_1852),
.B2(n_1895),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2395),
.Y(n_2416)
);

XNOR2x1_ASAP7_75t_L g2417 ( 
.A(n_2375),
.B(n_322),
.Y(n_2417)
);

XOR2x1_ASAP7_75t_L g2418 ( 
.A(n_2389),
.B(n_323),
.Y(n_2418)
);

NAND4xp75_ASAP7_75t_L g2419 ( 
.A(n_2393),
.B(n_323),
.C(n_324),
.D(n_325),
.Y(n_2419)
);

NOR2x1_ASAP7_75t_L g2420 ( 
.A(n_2410),
.B(n_324),
.Y(n_2420)
);

NOR2x1_ASAP7_75t_L g2421 ( 
.A(n_2372),
.B(n_325),
.Y(n_2421)
);

NOR2x1_ASAP7_75t_L g2422 ( 
.A(n_2371),
.B(n_326),
.Y(n_2422)
);

OAI211xp5_ASAP7_75t_L g2423 ( 
.A1(n_2386),
.A2(n_326),
.B(n_327),
.C(n_328),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2403),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_2424)
);

OR2x2_ASAP7_75t_L g2425 ( 
.A(n_2364),
.B(n_329),
.Y(n_2425)
);

NOR2x1p5_ASAP7_75t_L g2426 ( 
.A(n_2374),
.B(n_330),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2399),
.B(n_330),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2402),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2376),
.B(n_331),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2396),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_2381),
.B(n_332),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2367),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_2432)
);

NOR2xp67_ASAP7_75t_L g2433 ( 
.A(n_2378),
.B(n_334),
.Y(n_2433)
);

AO22x2_ASAP7_75t_L g2434 ( 
.A1(n_2369),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2383),
.Y(n_2435)
);

XNOR2x1_ASAP7_75t_L g2436 ( 
.A(n_2401),
.B(n_337),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2370),
.B(n_338),
.Y(n_2437)
);

BUFx4f_ASAP7_75t_SL g2438 ( 
.A(n_2382),
.Y(n_2438)
);

OAI221xp5_ASAP7_75t_L g2439 ( 
.A1(n_2368),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.C(n_342),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2409),
.Y(n_2440)
);

NAND4xp75_ASAP7_75t_L g2441 ( 
.A(n_2380),
.B(n_339),
.C(n_340),
.D(n_341),
.Y(n_2441)
);

NAND3xp33_ASAP7_75t_L g2442 ( 
.A(n_2379),
.B(n_342),
.C(n_343),
.Y(n_2442)
);

INVxp33_ASAP7_75t_L g2443 ( 
.A(n_2366),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2365),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_2444)
);

NAND4xp75_ASAP7_75t_L g2445 ( 
.A(n_2405),
.B(n_346),
.C(n_347),
.D(n_348),
.Y(n_2445)
);

OAI221xp5_ASAP7_75t_L g2446 ( 
.A1(n_2368),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.C(n_350),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2377),
.Y(n_2447)
);

XNOR2xp5_ASAP7_75t_L g2448 ( 
.A(n_2384),
.B(n_349),
.Y(n_2448)
);

NOR2x1_ASAP7_75t_L g2449 ( 
.A(n_2387),
.B(n_2397),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2388),
.Y(n_2450)
);

NOR3xp33_ASAP7_75t_L g2451 ( 
.A(n_2411),
.B(n_2392),
.C(n_2398),
.Y(n_2451)
);

NOR4xp25_ASAP7_75t_L g2452 ( 
.A(n_2450),
.B(n_2363),
.C(n_2390),
.D(n_2391),
.Y(n_2452)
);

NAND4xp75_ASAP7_75t_L g2453 ( 
.A(n_2422),
.B(n_2394),
.C(n_2385),
.D(n_2404),
.Y(n_2453)
);

O2A1O1Ixp33_ASAP7_75t_L g2454 ( 
.A1(n_2437),
.A2(n_2362),
.B(n_351),
.C(n_352),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2425),
.B(n_350),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2414),
.B(n_351),
.Y(n_2456)
);

AND4x1_ASAP7_75t_L g2457 ( 
.A(n_2429),
.B(n_352),
.C(n_353),
.D(n_354),
.Y(n_2457)
);

BUFx3_ASAP7_75t_L g2458 ( 
.A(n_2427),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2418),
.B(n_353),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_L g2460 ( 
.A(n_2448),
.B(n_354),
.C(n_355),
.Y(n_2460)
);

NOR3xp33_ASAP7_75t_SL g2461 ( 
.A(n_2423),
.B(n_355),
.C(n_356),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2436),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2417),
.A2(n_356),
.B(n_357),
.Y(n_2463)
);

NAND4xp25_ASAP7_75t_L g2464 ( 
.A(n_2433),
.B(n_357),
.C(n_358),
.D(n_359),
.Y(n_2464)
);

NOR2x1_ASAP7_75t_L g2465 ( 
.A(n_2419),
.B(n_2420),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2434),
.Y(n_2466)
);

NOR2x1_ASAP7_75t_L g2467 ( 
.A(n_2426),
.B(n_358),
.Y(n_2467)
);

NAND4xp25_ASAP7_75t_SL g2468 ( 
.A(n_2431),
.B(n_360),
.C(n_361),
.D(n_362),
.Y(n_2468)
);

NAND3xp33_ASAP7_75t_SL g2469 ( 
.A(n_2430),
.B(n_360),
.C(n_361),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2434),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2412),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2438),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_2472)
);

XNOR2x1_ASAP7_75t_L g2473 ( 
.A(n_2413),
.B(n_363),
.Y(n_2473)
);

OAI211xp5_ASAP7_75t_SL g2474 ( 
.A1(n_2421),
.A2(n_365),
.B(n_366),
.C(n_368),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_SL g2475 ( 
.A(n_2435),
.B(n_365),
.C(n_368),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2441),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2432),
.B(n_369),
.Y(n_2477)
);

NOR4xp25_ASAP7_75t_L g2478 ( 
.A(n_2416),
.B(n_370),
.C(n_371),
.D(n_372),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2445),
.B(n_371),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2470),
.Y(n_2480)
);

CKINVDCx20_ASAP7_75t_R g2481 ( 
.A(n_2471),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2455),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2478),
.B(n_2444),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2459),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_2467),
.Y(n_2485)
);

CKINVDCx6p67_ASAP7_75t_R g2486 ( 
.A(n_2458),
.Y(n_2486)
);

XNOR2xp5_ASAP7_75t_L g2487 ( 
.A(n_2473),
.B(n_2442),
.Y(n_2487)
);

AOI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2465),
.A2(n_2443),
.B(n_2447),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2456),
.Y(n_2489)
);

OR2x2_ASAP7_75t_L g2490 ( 
.A(n_2464),
.B(n_2439),
.Y(n_2490)
);

BUFx2_ASAP7_75t_L g2491 ( 
.A(n_2475),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_2462),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2479),
.Y(n_2493)
);

INVxp67_ASAP7_75t_L g2494 ( 
.A(n_2468),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2466),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2476),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2477),
.Y(n_2497)
);

XNOR2xp5_ASAP7_75t_L g2498 ( 
.A(n_2453),
.B(n_2457),
.Y(n_2498)
);

CKINVDCx16_ASAP7_75t_R g2499 ( 
.A(n_2452),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2460),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2469),
.Y(n_2501)
);

OAI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2499),
.A2(n_2446),
.B1(n_2461),
.B2(n_2428),
.Y(n_2502)
);

A2O1A1Ixp33_ASAP7_75t_L g2503 ( 
.A1(n_2488),
.A2(n_2463),
.B(n_2454),
.C(n_2474),
.Y(n_2503)
);

AOI221xp5_ASAP7_75t_L g2504 ( 
.A1(n_2480),
.A2(n_2451),
.B1(n_2440),
.B2(n_2472),
.C(n_2424),
.Y(n_2504)
);

AOI322xp5_ASAP7_75t_L g2505 ( 
.A1(n_2495),
.A2(n_2449),
.A3(n_2415),
.B1(n_374),
.B2(n_375),
.C1(n_376),
.C2(n_377),
.Y(n_2505)
);

AOI322xp5_ASAP7_75t_L g2506 ( 
.A1(n_2501),
.A2(n_372),
.A3(n_373),
.B1(n_374),
.B2(n_375),
.C1(n_376),
.C2(n_377),
.Y(n_2506)
);

AOI322xp5_ASAP7_75t_L g2507 ( 
.A1(n_2494),
.A2(n_373),
.A3(n_378),
.B1(n_379),
.B2(n_380),
.C1(n_381),
.C2(n_382),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2486),
.B(n_378),
.Y(n_2508)
);

AOI322xp5_ASAP7_75t_L g2509 ( 
.A1(n_2500),
.A2(n_380),
.A3(n_381),
.B1(n_382),
.B2(n_383),
.C1(n_384),
.C2(n_385),
.Y(n_2509)
);

AOI221xp5_ASAP7_75t_L g2510 ( 
.A1(n_2496),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.C(n_387),
.Y(n_2510)
);

AOI322xp5_ASAP7_75t_L g2511 ( 
.A1(n_2481),
.A2(n_386),
.A3(n_388),
.B1(n_389),
.B2(n_390),
.C1(n_391),
.C2(n_392),
.Y(n_2511)
);

AOI221xp5_ASAP7_75t_L g2512 ( 
.A1(n_2485),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.C(n_391),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2482),
.Y(n_2513)
);

O2A1O1Ixp33_ASAP7_75t_L g2514 ( 
.A1(n_2493),
.A2(n_392),
.B(n_393),
.C(n_394),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2491),
.B(n_395),
.Y(n_2515)
);

NAND3xp33_ASAP7_75t_SL g2516 ( 
.A(n_2492),
.B(n_395),
.C(n_396),
.Y(n_2516)
);

INVx4_ASAP7_75t_L g2517 ( 
.A(n_2484),
.Y(n_2517)
);

AOI322xp5_ASAP7_75t_L g2518 ( 
.A1(n_2483),
.A2(n_396),
.A3(n_397),
.B1(n_398),
.B2(n_399),
.C1(n_400),
.C2(n_401),
.Y(n_2518)
);

OAI221xp5_ASAP7_75t_L g2519 ( 
.A1(n_2498),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.C(n_401),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2513),
.A2(n_2487),
.B1(n_2489),
.B2(n_2497),
.Y(n_2520)
);

OAI22x1_ASAP7_75t_L g2521 ( 
.A1(n_2515),
.A2(n_2490),
.B1(n_403),
.B2(n_404),
.Y(n_2521)
);

AO22x2_ASAP7_75t_L g2522 ( 
.A1(n_2502),
.A2(n_402),
.B1(n_403),
.B2(n_404),
.Y(n_2522)
);

AOI211xp5_ASAP7_75t_SL g2523 ( 
.A1(n_2504),
.A2(n_402),
.B(n_405),
.C(n_406),
.Y(n_2523)
);

AO22x2_ASAP7_75t_L g2524 ( 
.A1(n_2516),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2508),
.Y(n_2525)
);

AOI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2517),
.A2(n_408),
.B1(n_409),
.B2(n_412),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2519),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2503),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_2528)
);

HB1xp67_ASAP7_75t_L g2529 ( 
.A(n_2510),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2518),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2514),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2507),
.Y(n_2532)
);

OAI21x1_ASAP7_75t_L g2533 ( 
.A1(n_2530),
.A2(n_2512),
.B(n_2505),
.Y(n_2533)
);

AOI221xp5_ASAP7_75t_L g2534 ( 
.A1(n_2524),
.A2(n_2506),
.B1(n_2509),
.B2(n_2511),
.C(n_417),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2522),
.Y(n_2535)
);

NAND5xp2_ASAP7_75t_L g2536 ( 
.A(n_2520),
.B(n_413),
.C(n_415),
.D(n_416),
.E(n_417),
.Y(n_2536)
);

NAND3xp33_ASAP7_75t_L g2537 ( 
.A(n_2523),
.B(n_415),
.C(n_416),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2521),
.B(n_418),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2538),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2534),
.B(n_2525),
.Y(n_2540)
);

XNOR2xp5_ASAP7_75t_L g2541 ( 
.A(n_2537),
.B(n_2532),
.Y(n_2541)
);

AOI21xp33_ASAP7_75t_L g2542 ( 
.A1(n_2535),
.A2(n_2531),
.B(n_2529),
.Y(n_2542)
);

OAI22xp5_ASAP7_75t_SL g2543 ( 
.A1(n_2541),
.A2(n_2527),
.B1(n_2528),
.B2(n_2526),
.Y(n_2543)
);

AOI22xp5_ASAP7_75t_L g2544 ( 
.A1(n_2540),
.A2(n_2533),
.B1(n_2536),
.B2(n_420),
.Y(n_2544)
);

OAI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2539),
.A2(n_2542),
.B1(n_419),
.B2(n_421),
.Y(n_2545)
);

AOI22xp5_ASAP7_75t_L g2546 ( 
.A1(n_2541),
.A2(n_418),
.B1(n_419),
.B2(n_421),
.Y(n_2546)
);

OAI22x1_ASAP7_75t_L g2547 ( 
.A1(n_2541),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2543),
.A2(n_423),
.B(n_424),
.Y(n_2548)
);

OAI21xp33_ASAP7_75t_L g2549 ( 
.A1(n_2544),
.A2(n_425),
.B(n_426),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2545),
.B(n_426),
.Y(n_2550)
);

OAI22xp5_ASAP7_75t_SL g2551 ( 
.A1(n_2547),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_2551)
);

AOI21xp5_ASAP7_75t_L g2552 ( 
.A1(n_2550),
.A2(n_2546),
.B(n_428),
.Y(n_2552)
);

XNOR2xp5_ASAP7_75t_L g2553 ( 
.A(n_2551),
.B(n_427),
.Y(n_2553)
);

AOI222xp33_ASAP7_75t_L g2554 ( 
.A1(n_2549),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.C1(n_432),
.C2(n_433),
.Y(n_2554)
);

AO22x2_ASAP7_75t_L g2555 ( 
.A1(n_2552),
.A2(n_2548),
.B1(n_431),
.B2(n_432),
.Y(n_2555)
);

OA21x2_ASAP7_75t_L g2556 ( 
.A1(n_2555),
.A2(n_2553),
.B(n_2554),
.Y(n_2556)
);

OAI31xp33_ASAP7_75t_L g2557 ( 
.A1(n_2556),
.A2(n_430),
.A3(n_433),
.B(n_434),
.Y(n_2557)
);

AOI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2557),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.C(n_437),
.Y(n_2558)
);

AOI221xp5_ASAP7_75t_L g2559 ( 
.A1(n_2558),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.C(n_438),
.Y(n_2559)
);

AOI211xp5_ASAP7_75t_L g2560 ( 
.A1(n_2559),
.A2(n_438),
.B(n_439),
.C(n_440),
.Y(n_2560)
);


endmodule