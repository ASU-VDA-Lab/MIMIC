module fake_jpeg_30823_n_74 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_20),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_24),
.B1(n_23),
.B2(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_37),
.B(n_39),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_44),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_28),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_4),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_56),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_31),
.B(n_3),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_1),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_4),
.B(n_5),
.Y(n_55)
);

AOI21x1_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_48),
.B(n_7),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_6),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_10),
.B(n_11),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_57),
.B(n_54),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_64),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_55),
.B(n_12),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_68),
.B(n_60),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B(n_67),
.C(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_62),
.B1(n_11),
.B2(n_16),
.C(n_14),
.Y(n_74)
);


endmodule