module real_aes_8726_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g479 ( .A1(n_0), .A2(n_183), .B(n_480), .C(n_483), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_1), .B(n_474), .Y(n_485) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g232 ( .A(n_3), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_4), .B(n_171), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_5), .A2(n_458), .B(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_6), .A2(n_9), .B1(n_441), .B2(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_6), .Y(n_753) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_7), .A2(n_188), .B(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_8), .A2(n_38), .B1(n_144), .B2(n_156), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_9), .A2(n_128), .B1(n_129), .B2(n_441), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_9), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_10), .B(n_188), .Y(n_221) );
AND2x6_ASAP7_75t_L g159 ( .A(n_11), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_12), .A2(n_159), .B(n_461), .C(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_13), .B(n_39), .Y(n_113) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_15), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g226 ( .A(n_16), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_17), .B(n_171), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_18), .B(n_186), .Y(n_204) );
AO32x2_ASAP7_75t_L g180 ( .A1(n_19), .A2(n_181), .A3(n_185), .B1(n_187), .B2(n_188), .Y(n_180) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_20), .A2(n_92), .B1(n_125), .B2(n_739), .C1(n_740), .C2(n_742), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_20), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_21), .B(n_144), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_22), .B(n_186), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_23), .A2(n_54), .B1(n_144), .B2(n_156), .Y(n_184) );
AOI22xp33_ASAP7_75t_SL g197 ( .A1(n_24), .A2(n_79), .B1(n_144), .B2(n_148), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_25), .B(n_144), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_26), .A2(n_187), .B(n_461), .C(n_463), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_27), .A2(n_187), .B(n_461), .C(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_29), .B(n_136), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_30), .A2(n_458), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_31), .B(n_136), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_32), .A2(n_101), .B1(n_114), .B2(n_756), .Y(n_100) );
INVx2_ASAP7_75t_L g146 ( .A(n_33), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_34), .A2(n_492), .B(n_493), .C(n_497), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_35), .B(n_144), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_36), .B(n_136), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_37), .B(n_151), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_40), .B(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_41), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_42), .B(n_171), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_43), .B(n_458), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_44), .A2(n_492), .B(n_497), .C(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_45), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_46), .B(n_144), .Y(n_214) );
INVx1_ASAP7_75t_L g481 ( .A(n_47), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_48), .A2(n_88), .B1(n_156), .B2(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g520 ( .A(n_49), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_50), .B(n_144), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_51), .B(n_144), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_52), .B(n_458), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_53), .B(n_219), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g208 ( .A1(n_55), .A2(n_59), .B1(n_144), .B2(n_148), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_56), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_57), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_58), .B(n_144), .Y(n_245) );
INVx1_ASAP7_75t_L g160 ( .A(n_60), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_61), .B(n_458), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_62), .B(n_474), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_63), .A2(n_219), .B(n_229), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_64), .B(n_144), .Y(n_233) );
INVx1_ASAP7_75t_L g139 ( .A(n_65), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_67), .B(n_171), .Y(n_495) );
AO32x2_ASAP7_75t_L g193 ( .A1(n_68), .A2(n_187), .A3(n_188), .B1(n_194), .B2(n_198), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_69), .B(n_172), .Y(n_551) );
INVx1_ASAP7_75t_L g244 ( .A(n_70), .Y(n_244) );
INVx1_ASAP7_75t_L g169 ( .A(n_71), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_72), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_73), .B(n_465), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_74), .A2(n_461), .B(n_497), .C(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_75), .B(n_148), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_76), .Y(n_529) );
INVx1_ASAP7_75t_L g106 ( .A(n_77), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_78), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_80), .B(n_156), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_81), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_82), .B(n_148), .Y(n_175) );
INVx2_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_84), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_85), .B(n_158), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_86), .B(n_148), .Y(n_215) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g122 ( .A(n_87), .B(n_110), .Y(n_122) );
OR2x2_ASAP7_75t_L g444 ( .A(n_87), .B(n_111), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_89), .A2(n_99), .B1(n_148), .B2(n_149), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_90), .B(n_458), .Y(n_490) );
INVx1_ASAP7_75t_L g494 ( .A(n_91), .Y(n_494) );
INVxp67_ASAP7_75t_L g532 ( .A(n_93), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_94), .B(n_148), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_95), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g507 ( .A(n_96), .Y(n_507) );
INVx1_ASAP7_75t_L g547 ( .A(n_97), .Y(n_547) );
AND2x2_ASAP7_75t_L g522 ( .A(n_98), .B(n_136), .Y(n_522) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx12_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g757 ( .A(n_104), .Y(n_757) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx3_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g743 ( .A(n_108), .Y(n_743) );
NOR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g738 ( .A(n_109), .B(n_111), .Y(n_738) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AOI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_124), .B1(n_744), .B2(n_745), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g744 ( .A(n_118), .Y(n_744) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_120), .A2(n_746), .B(n_754), .Y(n_745) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_123), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g755 ( .A(n_122), .Y(n_755) );
OAI22x1_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_442), .B1(n_445), .B2(n_736), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_127), .A2(n_446), .B1(n_736), .B2(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_128), .A2(n_129), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_363), .Y(n_129) );
NAND5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_282), .C(n_297), .D(n_323), .E(n_345), .Y(n_130) );
NOR2xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_262), .Y(n_131) );
OAI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_199), .B1(n_235), .B2(n_251), .C(n_252), .Y(n_132) );
NOR2xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_189), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_134), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g439 ( .A(n_134), .Y(n_439) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_162), .Y(n_134) );
INVx1_ASAP7_75t_L g279 ( .A(n_135), .Y(n_279) );
AND2x2_ASAP7_75t_L g281 ( .A(n_135), .B(n_180), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_135), .B(n_179), .Y(n_291) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_135), .Y(n_309) );
INVx1_ASAP7_75t_L g319 ( .A(n_135), .Y(n_319) );
OR2x2_ASAP7_75t_L g357 ( .A(n_135), .B(n_256), .Y(n_357) );
INVx2_ASAP7_75t_L g407 ( .A(n_135), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_135), .B(n_255), .Y(n_424) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .B(n_161), .Y(n_135) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_136), .A2(n_166), .B(n_178), .Y(n_165) );
INVx2_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
INVx1_ASAP7_75t_L g471 ( .A(n_136), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_136), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_136), .A2(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_L g186 ( .A(n_137), .B(n_138), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_153), .B(n_159), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_147), .B(n_150), .Y(n_142) );
INVx3_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_144), .Y(n_509) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
BUFx3_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
AND2x6_ASAP7_75t_L g461 ( .A(n_145), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx1_ASAP7_75t_L g220 ( .A(n_146), .Y(n_220) );
INVx2_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx3_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
AND2x2_ASAP7_75t_L g459 ( .A(n_152), .B(n_220), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_152), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_157), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_157), .A2(n_231), .B(n_244), .C(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_158), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_158), .A2(n_172), .B1(n_195), .B2(n_197), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_158), .A2(n_183), .B1(n_207), .B2(n_208), .Y(n_206) );
INVx4_ASAP7_75t_L g482 ( .A(n_158), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_167), .B(n_173), .Y(n_166) );
BUFx3_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_159), .A2(n_213), .B(n_216), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_159), .A2(n_225), .B(n_230), .Y(n_224) );
AND2x4_ASAP7_75t_L g458 ( .A(n_159), .B(n_459), .Y(n_458) );
INVx4_ASAP7_75t_SL g484 ( .A(n_159), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_159), .B(n_459), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g162 ( .A(n_163), .B(n_179), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_164), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_164), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_SL g339 ( .A(n_164), .B(n_279), .Y(n_339) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
INVx2_ASAP7_75t_L g256 ( .A(n_165), .Y(n_256) );
OR2x2_ASAP7_75t_L g318 ( .A(n_165), .B(n_319), .Y(n_318) );
O2A1O1Ixp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_171), .Y(n_167) );
INVx2_ASAP7_75t_L g183 ( .A(n_171), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_171), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_171), .A2(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_171), .B(n_532), .Y(n_531) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .Y(n_173) );
INVx1_ASAP7_75t_L g229 ( .A(n_176), .Y(n_229) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g465 ( .A(n_177), .Y(n_465) );
AND2x2_ASAP7_75t_L g257 ( .A(n_179), .B(n_193), .Y(n_257) );
AND2x2_ASAP7_75t_L g274 ( .A(n_179), .B(n_254), .Y(n_274) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g192 ( .A(n_180), .B(n_193), .Y(n_192) );
BUFx2_ASAP7_75t_L g277 ( .A(n_180), .Y(n_277) );
AND2x2_ASAP7_75t_L g406 ( .A(n_180), .B(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_183), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_183), .A2(n_231), .B(n_232), .C(n_233), .Y(n_230) );
INVx2_ASAP7_75t_L g223 ( .A(n_185), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_185), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_186), .Y(n_188) );
NAND3xp33_ASAP7_75t_L g205 ( .A(n_187), .B(n_206), .C(n_209), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_187), .A2(n_240), .B(n_243), .Y(n_239) );
INVx4_ASAP7_75t_L g209 ( .A(n_188), .Y(n_209) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_188), .A2(n_212), .B(n_221), .Y(n_211) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_188), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_188), .A2(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g251 ( .A(n_189), .Y(n_251) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_192), .Y(n_189) );
AND2x2_ASAP7_75t_L g369 ( .A(n_190), .B(n_257), .Y(n_369) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g370 ( .A(n_191), .B(n_281), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_192), .A2(n_338), .B(n_340), .C(n_342), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_192), .B(n_338), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_192), .A2(n_268), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g254 ( .A(n_193), .Y(n_254) );
INVx1_ASAP7_75t_L g290 ( .A(n_193), .Y(n_290) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_193), .Y(n_299) );
INVx2_ASAP7_75t_L g483 ( .A(n_196), .Y(n_483) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_196), .Y(n_496) );
INVx1_ASAP7_75t_L g468 ( .A(n_198), .Y(n_468) );
INVx1_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_210), .Y(n_200) );
AND2x2_ASAP7_75t_L g316 ( .A(n_201), .B(n_261), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_201), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_202), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g408 ( .A(n_202), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g440 ( .A(n_202), .Y(n_440) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g270 ( .A(n_203), .Y(n_270) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_250), .Y(n_296) );
NOR2x1_ASAP7_75t_L g305 ( .A(n_203), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g312 ( .A(n_203), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
AO21x1_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_209), .B(n_248), .Y(n_247) );
INVx3_ASAP7_75t_L g474 ( .A(n_209), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_209), .B(n_499), .Y(n_498) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_209), .A2(n_504), .B(n_511), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_209), .B(n_512), .Y(n_511) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_209), .A2(n_546), .B(n_553), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_210), .B(n_352), .Y(n_387) );
INVx1_ASAP7_75t_SL g391 ( .A(n_210), .Y(n_391) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_222), .Y(n_210) );
INVx3_ASAP7_75t_L g250 ( .A(n_211), .Y(n_250) );
AND2x2_ASAP7_75t_L g261 ( .A(n_211), .B(n_238), .Y(n_261) );
AND2x2_ASAP7_75t_L g283 ( .A(n_211), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g328 ( .A(n_211), .B(n_322), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_211), .B(n_260), .Y(n_409) );
INVx2_ASAP7_75t_L g231 ( .A(n_219), .Y(n_231) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g249 ( .A(n_222), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_222), .B(n_238), .Y(n_285) );
AND2x2_ASAP7_75t_L g321 ( .A(n_222), .B(n_322), .Y(n_321) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_234), .Y(n_222) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_223), .A2(n_239), .B(n_246), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .C(n_229), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_227), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_227), .A2(n_551), .B(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_229), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_231), .A2(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_249), .Y(n_236) );
INVx1_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
AND2x2_ASAP7_75t_L g343 ( .A(n_237), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_237), .B(n_264), .Y(n_349) );
AOI21xp5_ASAP7_75t_SL g423 ( .A1(n_237), .A2(n_255), .B(n_278), .Y(n_423) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_247), .Y(n_237) );
OR2x2_ASAP7_75t_L g266 ( .A(n_238), .B(n_247), .Y(n_266) );
AND2x2_ASAP7_75t_L g313 ( .A(n_238), .B(n_250), .Y(n_313) );
INVx2_ASAP7_75t_L g322 ( .A(n_238), .Y(n_322) );
INVx1_ASAP7_75t_L g428 ( .A(n_238), .Y(n_428) );
AND2x2_ASAP7_75t_L g352 ( .A(n_247), .B(n_322), .Y(n_352) );
INVx1_ASAP7_75t_L g377 ( .A(n_247), .Y(n_377) );
AND2x2_ASAP7_75t_L g286 ( .A(n_249), .B(n_270), .Y(n_286) );
AND2x2_ASAP7_75t_L g298 ( .A(n_249), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_SL g416 ( .A(n_249), .Y(n_416) );
INVx2_ASAP7_75t_L g306 ( .A(n_250), .Y(n_306) );
AND2x2_ASAP7_75t_L g344 ( .A(n_250), .B(n_260), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_250), .B(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B(n_258), .Y(n_252) );
AND2x2_ASAP7_75t_L g359 ( .A(n_253), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g413 ( .A(n_253), .Y(n_413) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g333 ( .A(n_254), .Y(n_333) );
BUFx2_ASAP7_75t_L g432 ( .A(n_254), .Y(n_432) );
BUFx2_ASAP7_75t_L g303 ( .A(n_255), .Y(n_303) );
AND2x2_ASAP7_75t_L g405 ( .A(n_255), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g388 ( .A(n_256), .Y(n_388) );
AND2x4_ASAP7_75t_L g315 ( .A(n_257), .B(n_278), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_257), .B(n_339), .Y(n_351) );
AOI32xp33_ASAP7_75t_L g275 ( .A1(n_258), .A2(n_276), .A3(n_278), .B1(n_280), .B2(n_281), .Y(n_275) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
INVx3_ASAP7_75t_L g264 ( .A(n_259), .Y(n_264) );
OR2x2_ASAP7_75t_L g400 ( .A(n_259), .B(n_356), .Y(n_400) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g269 ( .A(n_260), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g376 ( .A(n_260), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g268 ( .A(n_261), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g280 ( .A(n_261), .B(n_270), .Y(n_280) );
INVx1_ASAP7_75t_L g401 ( .A(n_261), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_261), .B(n_376), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B(n_271), .C(n_275), .Y(n_262) );
OAI322xp33_ASAP7_75t_L g371 ( .A1(n_263), .A2(n_308), .A3(n_372), .B1(n_374), .B2(n_378), .C1(n_379), .C2(n_383), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVxp67_ASAP7_75t_L g336 ( .A(n_264), .Y(n_336) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g390 ( .A(n_266), .B(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_266), .B(n_306), .Y(n_437) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
OR2x2_ASAP7_75t_L g415 ( .A(n_270), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_273), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g324 ( .A(n_274), .B(n_303), .Y(n_324) );
AND2x2_ASAP7_75t_L g395 ( .A(n_274), .B(n_308), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_274), .B(n_382), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_276), .A2(n_283), .B1(n_286), .B2(n_287), .C(n_292), .Y(n_282) );
OR2x2_ASAP7_75t_L g293 ( .A(n_276), .B(n_289), .Y(n_293) );
AND2x2_ASAP7_75t_L g381 ( .A(n_276), .B(n_382), .Y(n_381) );
AOI32xp33_ASAP7_75t_L g420 ( .A1(n_276), .A2(n_306), .A3(n_421), .B1(n_422), .B2(n_425), .Y(n_420) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_277), .B(n_313), .C(n_336), .Y(n_354) );
AND2x2_ASAP7_75t_L g380 ( .A(n_277), .B(n_373), .Y(n_380) );
INVxp67_ASAP7_75t_L g360 ( .A(n_278), .Y(n_360) );
BUFx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_281), .B(n_333), .Y(n_389) );
INVx2_ASAP7_75t_L g399 ( .A(n_281), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_281), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g368 ( .A(n_284), .Y(n_368) );
OR2x2_ASAP7_75t_L g294 ( .A(n_285), .B(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_287), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_290), .Y(n_373) );
AND2x2_ASAP7_75t_L g332 ( .A(n_291), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_291), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AOI21xp33_ASAP7_75t_SL g317 ( .A1(n_293), .A2(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g411 ( .A(n_296), .B(n_321), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_300), .B(n_310), .C(n_317), .Y(n_297) );
AND2x2_ASAP7_75t_L g341 ( .A(n_299), .B(n_309), .Y(n_341) );
INVx2_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
OR2x2_ASAP7_75t_L g394 ( .A(n_299), .B(n_357), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_299), .B(n_437), .Y(n_436) );
AOI211xp5_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_302), .B(n_304), .C(n_307), .Y(n_300) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_303), .B(n_341), .Y(n_340) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_304), .A2(n_399), .B(n_423), .C(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_305), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g362 ( .A(n_306), .B(n_352), .Y(n_362) );
INVx1_ASAP7_75t_L g367 ( .A(n_306), .Y(n_367) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVxp33_ASAP7_75t_L g418 ( .A(n_312), .Y(n_418) );
AND2x2_ASAP7_75t_L g397 ( .A(n_313), .B(n_376), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_318), .A2(n_380), .B(n_381), .Y(n_379) );
OAI322xp33_ASAP7_75t_L g398 ( .A1(n_320), .A2(n_399), .A3(n_400), .B1(n_401), .B2(n_402), .C1(n_404), .C2(n_408), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_330), .B2(n_334), .C(n_337), .Y(n_323) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g375 ( .A(n_328), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g419 ( .A(n_332), .Y(n_419) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_335), .B(n_355), .Y(n_421) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g384 ( .A(n_344), .B(n_352), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B1(n_350), .B2(n_352), .C(n_353), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_348), .A2(n_365), .B1(n_369), .B2(n_370), .C(n_371), .Y(n_364) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_352), .B(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_358), .B2(n_361), .Y(n_353) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx2_ASAP7_75t_SL g382 ( .A(n_357), .Y(n_382) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND5xp2_ASAP7_75t_L g363 ( .A(n_364), .B(n_385), .C(n_410), .D(n_420), .E(n_430), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_366), .B(n_368), .Y(n_365) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_367), .B(n_373), .C(n_439), .D(n_440), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_370), .A2(n_431), .B1(n_433), .B2(n_435), .C(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
OAI322xp33_ASAP7_75t_L g386 ( .A1(n_380), .A2(n_387), .A3(n_388), .B1(n_389), .B2(n_390), .C1(n_392), .C2(n_396), .Y(n_386) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_398), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g431 ( .A(n_406), .B(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B1(n_418), .B2(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g741 ( .A(n_443), .Y(n_741) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_SL g446 ( .A(n_447), .B(n_691), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_626), .Y(n_447) );
NAND4xp25_ASAP7_75t_SL g448 ( .A(n_449), .B(n_571), .C(n_595), .D(n_618), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_513), .B1(n_543), .B2(n_555), .C(n_558), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_486), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_452), .A2(n_472), .B1(n_514), .B2(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_452), .B(n_487), .Y(n_629) );
AND2x2_ASAP7_75t_L g648 ( .A(n_452), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_452), .B(n_632), .Y(n_718) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_472), .Y(n_452) );
AND2x2_ASAP7_75t_L g586 ( .A(n_453), .B(n_487), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_453), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g609 ( .A(n_453), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g614 ( .A(n_453), .B(n_473), .Y(n_614) );
INVx2_ASAP7_75t_L g646 ( .A(n_453), .Y(n_646) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_453), .Y(n_690) );
AND2x2_ASAP7_75t_L g707 ( .A(n_453), .B(n_584), .Y(n_707) );
INVx5_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g625 ( .A(n_454), .B(n_584), .Y(n_625) );
AND2x4_ASAP7_75t_L g639 ( .A(n_454), .B(n_472), .Y(n_639) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_454), .Y(n_643) );
AND2x2_ASAP7_75t_L g663 ( .A(n_454), .B(n_578), .Y(n_663) );
AND2x2_ASAP7_75t_L g713 ( .A(n_454), .B(n_488), .Y(n_713) );
AND2x2_ASAP7_75t_L g723 ( .A(n_454), .B(n_473), .Y(n_723) );
OR2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_469), .Y(n_454) );
AOI21xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_460), .B(n_468), .Y(n_455) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx5_ASAP7_75t_L g478 ( .A(n_461), .Y(n_478) );
INVx2_ASAP7_75t_L g467 ( .A(n_465), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_467), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_467), .A2(n_496), .B(n_520), .C(n_521), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x2_ASAP7_75t_L g579 ( .A(n_472), .B(n_487), .Y(n_579) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_472), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_472), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g669 ( .A(n_472), .Y(n_669) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g557 ( .A(n_473), .B(n_502), .Y(n_557) );
AND2x2_ASAP7_75t_L g584 ( .A(n_473), .B(n_503), .Y(n_584) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_485), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_478), .B(n_479), .C(n_484), .Y(n_476) );
INVx2_ASAP7_75t_L g492 ( .A(n_478), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_478), .A2(n_484), .B(n_529), .C(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g497 ( .A(n_484), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_486), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_500), .Y(n_486) );
OR2x2_ASAP7_75t_L g610 ( .A(n_487), .B(n_501), .Y(n_610) );
AND2x2_ASAP7_75t_L g647 ( .A(n_487), .B(n_557), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_487), .B(n_578), .Y(n_658) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_487), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_487), .B(n_614), .Y(n_731) );
INVx5_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g556 ( .A(n_488), .Y(n_556) );
AND2x2_ASAP7_75t_L g565 ( .A(n_488), .B(n_501), .Y(n_565) );
AND2x2_ASAP7_75t_L g681 ( .A(n_488), .B(n_576), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_488), .B(n_614), .Y(n_703) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_501), .Y(n_649) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_502), .Y(n_601) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g578 ( .A(n_503), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_514), .B(n_591), .Y(n_710) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_515), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g562 ( .A(n_515), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_SL g570 ( .A(n_515), .Y(n_570) );
OR2x2_ASAP7_75t_L g593 ( .A(n_515), .B(n_563), .Y(n_593) );
OR2x2_ASAP7_75t_L g603 ( .A(n_515), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g666 ( .A(n_515), .B(n_525), .Y(n_666) );
AND2x2_ASAP7_75t_SL g704 ( .A(n_515), .B(n_524), .Y(n_704) );
NOR4xp25_ASAP7_75t_L g725 ( .A(n_515), .B(n_646), .C(n_726), .D(n_727), .Y(n_725) );
AND2x2_ASAP7_75t_L g735 ( .A(n_515), .B(n_567), .Y(n_735) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g560 ( .A(n_524), .B(n_556), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_524), .B(n_562), .Y(n_729) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_534), .Y(n_524) );
OR2x2_ASAP7_75t_L g569 ( .A(n_525), .B(n_570), .Y(n_569) );
INVx3_ASAP7_75t_L g576 ( .A(n_525), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_525), .B(n_545), .Y(n_588) );
INVxp67_ASAP7_75t_L g591 ( .A(n_525), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_525), .B(n_563), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_525), .B(n_535), .Y(n_657) );
AND2x2_ASAP7_75t_L g672 ( .A(n_525), .B(n_567), .Y(n_672) );
OR2x2_ASAP7_75t_L g701 ( .A(n_525), .B(n_535), .Y(n_701) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_533), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_534), .B(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_534), .B(n_570), .Y(n_709) );
OR2x2_ASAP7_75t_L g730 ( .A(n_534), .B(n_607), .Y(n_730) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g544 ( .A(n_535), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g567 ( .A(n_535), .B(n_563), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_535), .B(n_545), .Y(n_582) );
AND2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_576), .Y(n_652) );
AND2x2_ASAP7_75t_L g686 ( .A(n_535), .B(n_570), .Y(n_686) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_536), .B(n_570), .Y(n_589) );
AND2x2_ASAP7_75t_L g617 ( .A(n_536), .B(n_545), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_543), .B(n_625), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_544), .A2(n_632), .B1(n_668), .B2(n_685), .C(n_687), .Y(n_684) );
INVx5_ASAP7_75t_SL g563 ( .A(n_545), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OAI33xp33_ASAP7_75t_L g583 ( .A1(n_556), .A2(n_584), .A3(n_585), .B1(n_587), .B2(n_590), .B3(n_594), .Y(n_583) );
OR2x2_ASAP7_75t_L g599 ( .A(n_556), .B(n_600), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g708 ( .A1(n_556), .A2(n_625), .A3(n_632), .B1(n_709), .B2(n_710), .C1(n_711), .C2(n_714), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_556), .B(n_584), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_SL g732 ( .A1(n_556), .A2(n_584), .B(n_733), .C(n_735), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_557), .A2(n_572), .B1(n_577), .B2(n_580), .C(n_583), .Y(n_571) );
INVx1_ASAP7_75t_L g664 ( .A(n_557), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_557), .B(n_713), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_561), .B1(n_564), .B2(n_566), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g641 ( .A(n_562), .B(n_576), .Y(n_641) );
AND2x2_ASAP7_75t_L g699 ( .A(n_562), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g607 ( .A(n_563), .B(n_570), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_563), .B(n_576), .Y(n_635) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_565), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_565), .B(n_643), .Y(n_697) );
OAI321xp33_ASAP7_75t_L g716 ( .A1(n_565), .A2(n_638), .A3(n_717), .B1(n_718), .B2(n_719), .C(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g683 ( .A(n_566), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_567), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g622 ( .A(n_567), .B(n_570), .Y(n_622) );
AOI321xp33_ASAP7_75t_L g680 ( .A1(n_567), .A2(n_584), .A3(n_681), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g597 ( .A(n_569), .B(n_582), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_570), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_570), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_570), .B(n_656), .Y(n_693) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g616 ( .A(n_574), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g581 ( .A(n_575), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g689 ( .A(n_576), .Y(n_689) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_579), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g612 ( .A(n_584), .Y(n_612) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_586), .B(n_621), .Y(n_670) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
OR2x2_ASAP7_75t_L g634 ( .A(n_589), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g679 ( .A(n_589), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_590), .A2(n_637), .B1(n_640), .B2(n_642), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g734 ( .A(n_593), .B(n_657), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B1(n_602), .B2(n_608), .C(n_611), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx2_ASAP7_75t_L g632 ( .A(n_601), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_SL g678 ( .A(n_604), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_606), .B(n_656), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_606), .A2(n_674), .B(n_676), .Y(n_673) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g719 ( .A(n_607), .B(n_701), .Y(n_719) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_SL g621 ( .A(n_610), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_615), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g665 ( .A(n_617), .B(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g727 ( .A(n_617), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_621), .B(n_639), .Y(n_675) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g696 ( .A(n_625), .Y(n_696) );
NAND5xp2_ASAP7_75t_L g626 ( .A(n_627), .B(n_644), .C(n_653), .D(n_673), .E(n_680), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B(n_633), .C(n_636), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g668 ( .A(n_632), .Y(n_668) );
CKINVDCx16_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_640), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g682 ( .A(n_642), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_648), .B(n_650), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_645), .A2(n_699), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_698) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AOI321xp33_ASAP7_75t_L g653 ( .A1(n_646), .A2(n_654), .A3(n_658), .B1(n_659), .B2(n_665), .C(n_667), .Y(n_653) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g724 ( .A(n_658), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_660), .B(n_664), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g676 ( .A(n_661), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NOR2xp67_ASAP7_75t_SL g688 ( .A(n_662), .B(n_669), .Y(n_688) );
AOI321xp33_ASAP7_75t_SL g720 ( .A1(n_665), .A2(n_721), .A3(n_722), .B1(n_723), .B2(n_724), .C(n_725), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_670), .C(n_671), .Y(n_667) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_678), .B(n_686), .Y(n_715) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .C(n_690), .Y(n_687) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_716), .C(n_728), .Y(n_691) );
OAI211xp5_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_694), .B(n_698), .C(n_708), .Y(n_692) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_696), .B(n_697), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_697), .A2(n_729), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g717 ( .A(n_699), .Y(n_717) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g721 ( .A(n_719), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx14_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
endmodule