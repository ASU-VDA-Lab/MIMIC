module fake_netlist_6_4073_n_186 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_186);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_186;

wire n_52;
wire n_119;
wire n_91;
wire n_46;
wire n_163;
wire n_146;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_130;
wire n_85;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp33_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_3),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_4),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_5),
.Y(n_73)
);

AND3x2_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_6),
.C(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_32),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_52),
.Y(n_77)
);

AND2x6_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2x1p5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_R g84 ( 
.A(n_63),
.B(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_54),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_49),
.B1(n_41),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_76),
.B1(n_61),
.B2(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

O2A1O1Ixp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_57),
.B(n_59),
.C(n_69),
.Y(n_96)
);

AO31x2_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_60),
.A3(n_56),
.B(n_66),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_60),
.B(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_57),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_64),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_59),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_89),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_92),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_93),
.B1(n_82),
.B2(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_87),
.Y(n_111)
);

AOI21x1_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_75),
.B(n_78),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_82),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_96),
.B(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_106),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_114),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_114),
.Y(n_129)
);

NAND2x1_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_117),
.B1(n_82),
.B2(n_113),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_41),
.B1(n_108),
.B2(n_74),
.Y(n_139)
);

AOI31xp33_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_129),
.A3(n_126),
.B(n_136),
.Y(n_140)
);

AOI222xp33_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_72),
.B1(n_68),
.B2(n_78),
.C1(n_37),
.C2(n_33),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_119),
.B1(n_111),
.B2(n_104),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_68),
.B1(n_72),
.B2(n_92),
.C(n_91),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_100),
.B(n_96),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_130),
.C(n_85),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_135),
.B(n_134),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_132),
.B(n_102),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_74),
.A3(n_70),
.B1(n_91),
.B2(n_86),
.C1(n_85),
.C2(n_14),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_67),
.Y(n_150)
);

AOI211xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_70),
.B(n_86),
.C(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_133),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_102),
.B(n_133),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_70),
.B(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_97),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_97),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_102),
.B(n_103),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_67),
.C(n_64),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_97),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_97),
.Y(n_163)
);

NOR2x1p5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_64),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_147),
.B1(n_151),
.B2(n_64),
.C(n_11),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_64),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_166)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_146),
.Y(n_167)
);

NAND2x1p5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_102),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_8),
.Y(n_169)
);

NAND4xp75_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_9),
.C(n_13),
.D(n_14),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_162),
.B1(n_161),
.B2(n_164),
.C(n_64),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_101),
.B(n_99),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g175 ( 
.A(n_169),
.Y(n_175)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_13),
.A3(n_16),
.B1(n_80),
.B2(n_81),
.C1(n_83),
.C2(n_99),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_97),
.Y(n_177)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_165),
.B1(n_172),
.B2(n_167),
.C(n_170),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_80),
.C(n_83),
.Y(n_179)
);

AOI22x1_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_176),
.B1(n_175),
.B2(n_179),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_168),
.B(n_174),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_177),
.Y(n_182)
);

OAI221xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_81),
.B1(n_83),
.B2(n_28),
.C(n_30),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_81),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_181),
.B(n_180),
.Y(n_185)
);

AOI221xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_183),
.B1(n_20),
.B2(n_17),
.C(n_105),
.Y(n_186)
);


endmodule