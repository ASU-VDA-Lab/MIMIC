module fake_jpeg_14225_n_473 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_44),
.C(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_48),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_53),
.B(n_69),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_74),
.Y(n_91)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_31),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_87),
.Y(n_92)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_16),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_85),
.Y(n_98)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_75),
.B1(n_79),
.B2(n_82),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_93),
.A2(n_106),
.B1(n_5),
.B2(n_8),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_145),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_99),
.B(n_104),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_39),
.B1(n_30),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_102),
.A2(n_127),
.B1(n_41),
.B2(n_2),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_36),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_34),
.B1(n_39),
.B2(n_30),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_105),
.A2(n_117),
.B1(n_123),
.B2(n_5),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_39),
.B1(n_34),
.B2(n_44),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_110),
.B(n_113),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_45),
.C(n_18),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_111),
.B(n_41),
.C(n_13),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_25),
.B1(n_38),
.B2(n_35),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_20),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_35),
.B1(n_25),
.B2(n_23),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_50),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_126),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_55),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_15),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_68),
.B(n_15),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_49),
.B(n_15),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_0),
.Y(n_145)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_147),
.Y(n_247)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_149),
.Y(n_211)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_52),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_199),
.C(n_134),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_0),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_169),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_100),
.A2(n_28),
.B1(n_77),
.B2(n_51),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_165),
.A2(n_166),
.B(n_187),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_100),
.A2(n_41),
.B1(n_14),
.B2(n_13),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_185),
.Y(n_234)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_1),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_171),
.B(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_102),
.B1(n_130),
.B2(n_140),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_91),
.A2(n_13),
.B1(n_41),
.B2(n_3),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_119),
.A2(n_41),
.B1(n_2),
.B2(n_3),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_178),
.A2(n_196),
.B1(n_97),
.B2(n_114),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_98),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_4),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_186),
.Y(n_203)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_130),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_187),
.A2(n_197),
.B1(n_116),
.B2(n_139),
.Y(n_240)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_193),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_138),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_191),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_94),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_146),
.B1(n_112),
.B2(n_96),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_93),
.A2(n_8),
.B1(n_9),
.B2(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_9),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_107),
.A2(n_109),
.B(n_120),
.C(n_134),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_97),
.B(n_94),
.C(n_90),
.Y(n_235)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_151),
.B1(n_171),
.B2(n_175),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_206),
.A2(n_227),
.B1(n_233),
.B2(n_197),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_169),
.Y(n_255)
);

OR2x4_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_94),
.Y(n_215)
);

INVx2_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_151),
.B(n_140),
.C(n_137),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_120),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_137),
.C(n_146),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_165),
.A2(n_109),
.B(n_107),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_222),
.A2(n_236),
.B(n_160),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_181),
.A2(n_112),
.B1(n_116),
.B2(n_139),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_243),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_97),
.B(n_90),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_192),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_244),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_191),
.B1(n_189),
.B2(n_186),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_160),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_251),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_161),
.B(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_157),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_155),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_281),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_255),
.B(n_284),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_173),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_256),
.B(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_214),
.A2(n_182),
.B1(n_190),
.B2(n_201),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_259),
.A2(n_260),
.B1(n_266),
.B2(n_296),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_214),
.A2(n_182),
.B1(n_190),
.B2(n_201),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_194),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_265),
.B(n_270),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_268),
.B(n_285),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_232),
.A2(n_157),
.B1(n_178),
.B2(n_189),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_168),
.C(n_158),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_213),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_226),
.Y(n_316)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_220),
.C(n_210),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_178),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_213),
.B(n_178),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_206),
.A2(n_234),
.B1(n_232),
.B2(n_245),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_283),
.B1(n_243),
.B2(n_208),
.Y(n_299)
);

NAND2x1_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_202),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_234),
.A2(n_185),
.B1(n_191),
.B2(n_200),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_221),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_239),
.B(n_166),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_218),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_211),
.B(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_288),
.B(n_292),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_150),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_156),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_231),
.Y(n_330)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_291),
.Y(n_329)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_205),
.Y(n_293)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_222),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_295),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_242),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_297),
.B(n_304),
.Y(n_356)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_298),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_313),
.B1(n_267),
.B2(n_292),
.Y(n_342)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_253),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_235),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_311),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_280),
.A2(n_243),
.B1(n_233),
.B2(n_211),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_320),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_260),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_241),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_325),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_241),
.Y(n_325)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_243),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_334),
.Y(n_340)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_237),
.Y(n_334)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_258),
.B(n_237),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_281),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_277),
.C(n_263),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_351),
.C(n_355),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_342),
.A2(n_343),
.B1(n_345),
.B2(n_350),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_267),
.B1(n_296),
.B2(n_284),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_254),
.B1(n_269),
.B2(n_283),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_267),
.B(n_281),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_357),
.B(n_358),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_359),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_349),
.A2(n_366),
.B(n_319),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_299),
.A2(n_292),
.B1(n_263),
.B2(n_273),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_289),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_318),
.C(n_302),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_290),
.B(n_207),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_312),
.A2(n_319),
.B(n_308),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_330),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_276),
.Y(n_361)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_274),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_225),
.C(n_209),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_323),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_365),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_301),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_334),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_262),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_367),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_369),
.A2(n_375),
.B(n_385),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_332),
.C(n_322),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_394),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_328),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_393),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_351),
.B(n_335),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_374),
.B(n_364),
.Y(n_404)
);

AO21x1_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_343),
.B(n_342),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_366),
.A2(n_300),
.B1(n_315),
.B2(n_309),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_378),
.A2(n_383),
.B1(n_387),
.B2(n_341),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_381),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_367),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_360),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_340),
.A2(n_300),
.B1(n_315),
.B2(n_309),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_347),
.A2(n_329),
.B(n_305),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_340),
.A2(n_305),
.B1(n_329),
.B2(n_306),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_350),
.A2(n_331),
.B1(n_321),
.B2(n_317),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_390),
.B1(n_225),
.B2(n_209),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_341),
.A2(n_321),
.B1(n_317),
.B2(n_307),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_212),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_354),
.B1(n_365),
.B2(n_344),
.Y(n_395)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_358),
.C(n_357),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_402),
.C(n_388),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_378),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_414),
.Y(n_428)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_362),
.C(n_361),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_404),
.B(n_409),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_382),
.A2(n_348),
.B1(n_375),
.B2(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_370),
.A2(n_339),
.B1(n_352),
.B2(n_346),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_407),
.A2(n_386),
.B1(n_380),
.B2(n_371),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_370),
.A2(n_339),
.B(n_336),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_408),
.A2(n_412),
.B(n_377),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_353),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_387),
.A2(n_336),
.B1(n_346),
.B2(n_337),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_413),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_385),
.B(n_368),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_390),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_228),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_393),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_374),
.B(n_228),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_416),
.B(n_394),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_419),
.C(n_434),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_406),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_418),
.B(n_398),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_SL g421 ( 
.A(n_415),
.B(n_411),
.Y(n_421)
);

AOI21x1_ASAP7_75t_SL g445 ( 
.A1(n_421),
.A2(n_425),
.B(n_428),
.Y(n_445)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_423),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_426),
.A2(n_408),
.B1(n_401),
.B2(n_397),
.Y(n_435)
);

AOI221xp5_ASAP7_75t_L g446 ( 
.A1(n_427),
.A2(n_430),
.B1(n_431),
.B2(n_429),
.C(n_432),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_412),
.A2(n_207),
.B(n_376),
.C(n_310),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_426),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_440),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_425),
.A2(n_397),
.B(n_407),
.C(n_404),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_424),
.C(n_431),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_402),
.C(n_409),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_443),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_422),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_442),
.B(n_444),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_433),
.A2(n_396),
.B(n_411),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_403),
.C(n_416),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_446),
.A2(n_447),
.B1(n_247),
.B2(n_205),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_424),
.A2(n_262),
.B1(n_293),
.B2(n_204),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_454),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_436),
.A2(n_443),
.B1(n_430),
.B2(n_445),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_450),
.B(n_451),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_421),
.C(n_420),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_420),
.C(n_417),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_444),
.C(n_438),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_456),
.A2(n_448),
.B1(n_449),
.B2(n_453),
.Y(n_458)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_458),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_455),
.A2(n_445),
.B(n_440),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_459),
.A2(n_451),
.B(n_452),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_461),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_435),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_463),
.A2(n_460),
.B(n_457),
.Y(n_468)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g464 ( 
.A1(n_458),
.A2(n_438),
.B(n_427),
.C(n_212),
.D(n_224),
.Y(n_464)
);

OAI21x1_ASAP7_75t_SL g467 ( 
.A1(n_464),
.A2(n_438),
.B(n_462),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_467),
.A2(n_468),
.B(n_466),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_468),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_470),
.C(n_465),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_457),
.C(n_464),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g473 ( 
.A(n_472),
.Y(n_473)
);


endmodule