module fake_jpeg_27024_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_29),
.B(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_64),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_47),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_39),
.B1(n_57),
.B2(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_48),
.B1(n_46),
.B2(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_39),
.B1(n_57),
.B2(n_51),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_79),
.B1(n_1),
.B2(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_52),
.B(n_53),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_50),
.B(n_45),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_74),
.B(n_71),
.C(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_50),
.B1(n_56),
.B2(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_0),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_92),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_88),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_71),
.Y(n_91)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_94),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_38),
.C(n_25),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_88),
.B1(n_90),
.B2(n_86),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_102),
.B1(n_89),
.B2(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_24),
.B1(n_35),
.B2(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_4),
.Y(n_107)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_106),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_95),
.C(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_19),
.C(n_26),
.Y(n_121)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_95),
.B1(n_6),
.B2(n_5),
.C(n_9),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_118),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_7),
.A3(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_17),
.B(n_18),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_121),
.B(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_116),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_126),
.B(n_114),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_113),
.B(n_114),
.C(n_123),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_125),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_27),
.B(n_28),
.Y(n_134)
);


endmodule