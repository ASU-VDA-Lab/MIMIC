module real_jpeg_13773_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_253, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_253;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_61),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_61),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_45),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_72),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_72),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_12),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_13),
.B(n_56),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_13),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_13),
.B(n_26),
.C(n_41),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_13),
.B(n_66),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_102),
.B(n_158),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_13),
.A2(n_51),
.B(n_67),
.C(n_185),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_143),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_13),
.B(n_207),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_63),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_63),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_63),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_15),
.Y(n_82)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.C(n_64),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_22),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_23),
.B(n_34),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_24),
.A2(n_29),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_24),
.A2(n_29),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_25),
.B(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_29),
.B(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_30),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_32),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_35),
.Y(n_229)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_37),
.B(n_147),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_38),
.A2(n_68),
.B(n_143),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_46),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_39),
.A2(n_44),
.B1(n_46),
.B2(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_39),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_39),
.B(n_145),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_39),
.A2(n_46),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_43),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_43),
.B(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_43),
.A2(n_155),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_46),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_60),
.B2(n_62),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_62),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_48),
.A2(n_57),
.B(n_143),
.C(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_60),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_49),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_50),
.B(n_52),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_52),
.B1(n_67),
.B2(n_68),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_51),
.A2(n_54),
.A3(n_57),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_69),
.B(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_69),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_65),
.A2(n_70),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_65),
.A2(n_93),
.B1(n_120),
.B2(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_71),
.Y(n_121)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_88),
.B2(n_89),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_87),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_99),
.B2(n_106),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_93),
.A2(n_121),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_97),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_103),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_102),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_102),
.A2(n_103),
.B1(n_128),
.B2(n_187),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_103),
.A2(n_164),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_103),
.B(n_143),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_103),
.A2(n_172),
.B(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_112),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_108),
.B(n_110),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_112),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_122),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_240)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_122),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_125),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_127),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI321xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_236),
.A3(n_245),
.B1(n_250),
.B2(n_251),
.C(n_253),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_218),
.B(n_235),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_197),
.B(n_217),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_180),
.B(n_196),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_160),
.B(n_179),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_138),
.B(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_146),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_140),
.B1(n_146),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B(n_144),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_141),
.A2(n_144),
.B(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_153),
.C(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_168),
.B(n_178),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_166),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_173),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_191),
.C(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_186),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_210),
.B2(n_211),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_213),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_205),
.C(n_209),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_220),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_232),
.C(n_233),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_230),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_227),
.C(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_239),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);


endmodule