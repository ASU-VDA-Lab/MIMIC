module fake_jpeg_27089_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_33),
.B1(n_36),
.B2(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_12),
.B1(n_18),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_11),
.B1(n_17),
.B2(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_12),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_44),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_11),
.A3(n_21),
.B1(n_13),
.B2(n_19),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_45),
.B1(n_28),
.B2(n_19),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_16),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_13),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_31),
.B1(n_40),
.B2(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_31),
.B1(n_34),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_8),
.Y(n_71)
);

OAI22x1_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_52),
.B1(n_45),
.B2(n_15),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_26),
.B1(n_30),
.B2(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_6),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_8),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_10),
.A3(n_9),
.B1(n_5),
.B2(n_4),
.C1(n_3),
.C2(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_1),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_59),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_58),
.C(n_56),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_73),
.A2(n_57),
.B(n_63),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_78),
.B(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_30),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_69),
.B(n_61),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_66),
.C(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_2),
.C(n_3),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_84),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_15),
.A3(n_69),
.B1(n_92),
.B2(n_95),
.C1(n_97),
.C2(n_99),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_15),
.B(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_15),
.Y(n_104)
);


endmodule