module fake_jpeg_2557_n_550 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_550);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_54),
.B(n_73),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_60),
.B(n_66),
.Y(n_148)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_40),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_38),
.B(n_39),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_78),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_0),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_79),
.Y(n_157)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_80),
.Y(n_151)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_83),
.B(n_94),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_43),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_36),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_160),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_29),
.B1(n_47),
.B2(n_36),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_114),
.A2(n_125),
.B1(n_141),
.B2(n_154),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_53),
.A2(n_44),
.B1(n_43),
.B2(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_116),
.A2(n_136),
.B1(n_152),
.B2(n_31),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_29),
.B1(n_47),
.B2(n_36),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_55),
.A2(n_44),
.B1(n_15),
.B2(n_30),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_29),
.B1(n_47),
.B2(n_36),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_65),
.A2(n_44),
.B1(n_15),
.B2(n_30),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_36),
.B1(n_15),
.B2(n_44),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_48),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_161),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_54),
.B(n_74),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_78),
.B(n_24),
.C(n_37),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_42),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_56),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_84),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_76),
.B1(n_31),
.B2(n_72),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_169),
.A2(n_201),
.B1(n_207),
.B2(n_210),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_101),
.B1(n_100),
.B2(n_97),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_188),
.B1(n_202),
.B2(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_175),
.B(n_195),
.Y(n_250)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_42),
.B1(n_28),
.B2(n_25),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_190),
.Y(n_222)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_63),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_192),
.B(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_121),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_59),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_197),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_199),
.Y(n_235)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_203),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_133),
.A2(n_34),
.B1(n_24),
.B2(n_37),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_67),
.B1(n_95),
.B2(n_92),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_212),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_34),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_213),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_118),
.A2(n_46),
.B1(n_61),
.B2(n_28),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_116),
.A2(n_22),
.B1(n_25),
.B2(n_33),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_105),
.B1(n_166),
.B2(n_151),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_106),
.B(n_108),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_46),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

NOR2x1_ASAP7_75t_R g214 ( 
.A(n_139),
.B(n_79),
.Y(n_214)
);

CKINVDCx9p33_ASAP7_75t_R g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_33),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_112),
.B(n_2),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_165),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_162),
.B1(n_138),
.B2(n_131),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_227),
.B1(n_230),
.B2(n_184),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_138),
.B1(n_162),
.B2(n_144),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_181),
.A2(n_141),
.B1(n_125),
.B2(n_114),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_229),
.B1(n_244),
.B2(n_247),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_174),
.A2(n_110),
.B1(n_122),
.B2(n_155),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_177),
.A2(n_165),
.B1(n_127),
.B2(n_120),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_159),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_189),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_169),
.A2(n_179),
.B1(n_192),
.B2(n_211),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_179),
.A2(n_110),
.B1(n_122),
.B2(n_155),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_217),
.B1(n_198),
.B2(n_197),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_192),
.B(n_124),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_167),
.Y(n_259)
);

AO22x2_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_213),
.B1(n_200),
.B2(n_178),
.Y(n_256)
);

AO21x2_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_270),
.B(n_277),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_257),
.A2(n_245),
.B1(n_232),
.B2(n_240),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_260),
.B(n_237),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_219),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_221),
.A2(n_206),
.B1(n_175),
.B2(n_195),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_267),
.B1(n_274),
.B2(n_245),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_194),
.B1(n_180),
.B2(n_193),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_263),
.A2(n_280),
.B1(n_227),
.B2(n_248),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_214),
.B(n_175),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_250),
.B(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_221),
.A2(n_166),
.B1(n_105),
.B2(n_191),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_204),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_272),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_173),
.B(n_170),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_271),
.B(n_254),
.Y(n_292)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_183),
.B(n_96),
.C(n_167),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_185),
.B(n_151),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_186),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_225),
.A2(n_196),
.B1(n_187),
.B2(n_182),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_186),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_278),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_205),
.B1(n_171),
.B2(n_182),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_219),
.B(n_146),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_172),
.C(n_199),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_255),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_244),
.B1(n_229),
.B2(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_190),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_285),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_205),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_235),
.A2(n_142),
.B1(n_128),
.B2(n_117),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_286),
.A2(n_142),
.B1(n_128),
.B2(n_240),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_288),
.A2(n_292),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_306),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_284),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_297),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_294),
.B(n_296),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_222),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_276),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_265),
.B1(n_274),
.B2(n_281),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_250),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_307),
.C(n_241),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_258),
.A2(n_254),
.B1(n_223),
.B2(n_232),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_280),
.B1(n_263),
.B2(n_275),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_222),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_305),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_260),
.B(n_235),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_258),
.A2(n_241),
.B1(n_220),
.B2(n_255),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_313),
.B1(n_259),
.B2(n_282),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_258),
.A2(n_280),
.B1(n_285),
.B2(n_267),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_257),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_264),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_268),
.B(n_220),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_241),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_269),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_329),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_327),
.A2(n_331),
.B1(n_334),
.B2(n_343),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_296),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_315),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_288),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_275),
.B1(n_277),
.B2(n_256),
.Y(n_331)
);

OAI21x1_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_289),
.B(n_292),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_332),
.A2(n_264),
.B(n_117),
.C(n_49),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_271),
.B(n_286),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_333),
.A2(n_342),
.B(n_351),
.Y(n_381)
);

AOI21xp33_ASAP7_75t_L g335 ( 
.A1(n_294),
.A2(n_259),
.B(n_270),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_113),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_305),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_293),
.B(n_279),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_350),
.Y(n_380)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_340),
.B(n_300),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_345),
.B1(n_314),
.B2(n_309),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_259),
.B(n_270),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_256),
.B1(n_283),
.B2(n_266),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_218),
.C(n_242),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_325),
.C(n_336),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_309),
.A2(n_256),
.B1(n_264),
.B2(n_230),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_256),
.B1(n_264),
.B2(n_273),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_347),
.A2(n_309),
.B1(n_308),
.B2(n_304),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_349),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_293),
.B(n_256),
.Y(n_350)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_351),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_354),
.Y(n_391)
);

AO21x2_ASAP7_75t_SL g357 ( 
.A1(n_343),
.A2(n_309),
.B(n_289),
.Y(n_357)
);

CKINVDCx6p67_ASAP7_75t_R g394 ( 
.A(n_357),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_358),
.A2(n_369),
.B1(n_370),
.B2(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_321),
.B(n_333),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_362),
.A2(n_374),
.B(n_379),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_363),
.A2(n_365),
.B1(n_373),
.B2(n_331),
.Y(n_386)
);

AO21x2_ASAP7_75t_L g364 ( 
.A1(n_345),
.A2(n_309),
.B(n_350),
.Y(n_364)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_322),
.A2(n_304),
.B1(n_291),
.B2(n_306),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_366),
.Y(n_414)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_346),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_368),
.B(n_372),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_298),
.B1(n_312),
.B2(n_307),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_327),
.A2(n_312),
.B1(n_315),
.B2(n_303),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_302),
.C(n_303),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_300),
.B1(n_264),
.B2(n_234),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_375),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_218),
.Y(n_376)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_218),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_384),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_242),
.B(n_252),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_381),
.A2(n_383),
.B(n_334),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_346),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_386),
.A2(n_388),
.B1(n_405),
.B2(n_409),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_401),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_378),
.A2(n_363),
.B1(n_356),
.B2(n_358),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_342),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_408),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_320),
.Y(n_397)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_320),
.Y(n_400)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_337),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_364),
.B1(n_383),
.B2(n_361),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_406),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_323),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_380),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_380),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_326),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_413),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_326),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_352),
.B(n_329),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_410),
.B(n_49),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_338),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_354),
.C(n_352),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_425),
.C(n_428),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_433),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_362),
.B(n_357),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_426),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_412),
.A2(n_364),
.B1(n_324),
.B2(n_357),
.Y(n_422)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_422),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_386),
.A2(n_388),
.B1(n_406),
.B2(n_389),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_379),
.C(n_341),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_355),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_397),
.A2(n_364),
.B1(n_357),
.B2(n_371),
.Y(n_427)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_367),
.C(n_359),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_361),
.C(n_373),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_431),
.C(n_435),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_383),
.C(n_364),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_383),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_117),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_440),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_234),
.C(n_239),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_234),
.C(n_239),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_439),
.C(n_385),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_226),
.C(n_251),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_416),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_457),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_448),
.A2(n_437),
.B1(n_433),
.B2(n_461),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_408),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_453),
.Y(n_481)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_400),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_398),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_459),
.Y(n_483)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_436),
.A2(n_398),
.B1(n_387),
.B2(n_392),
.Y(n_457)
);

INVx11_ASAP7_75t_L g458 ( 
.A(n_435),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_421),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_460),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_415),
.A2(n_394),
.B1(n_414),
.B2(n_395),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_461),
.A2(n_463),
.B1(n_447),
.B2(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_417),
.B(n_394),
.C(n_395),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_438),
.C(n_437),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_432),
.A2(n_394),
.B1(n_414),
.B2(n_385),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_464),
.A2(n_465),
.B1(n_466),
.B2(n_449),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_446),
.A2(n_420),
.B1(n_437),
.B2(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_478),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_434),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_473),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_463),
.A2(n_437),
.B(n_396),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_474),
.C(n_253),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_442),
.C(n_455),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_472),
.B(n_477),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_454),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_450),
.A2(n_396),
.B(n_440),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_226),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_476),
.A2(n_253),
.B1(n_168),
.B2(n_45),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_226),
.C(n_251),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_252),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_445),
.A2(n_251),
.B(n_176),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_459),
.Y(n_487)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_480),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_489),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_449),
.B(n_454),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_486),
.A2(n_468),
.B(n_45),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_499),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_252),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_491),
.B(n_495),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_251),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_458),
.C(n_171),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_497),
.C(n_481),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_253),
.C(n_168),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_471),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_501),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_499),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_479),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_494),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_469),
.B(n_474),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_515),
.B(n_516),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_481),
.Y(n_508)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_508),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_512),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_488),
.A2(n_476),
.B1(n_464),
.B2(n_465),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_514),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_478),
.C(n_477),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_486),
.A2(n_45),
.B(n_3),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_492),
.A2(n_45),
.B(n_3),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_2),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_518),
.B(n_520),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_492),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_497),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_523),
.B(n_524),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_504),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_45),
.C(n_3),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_525),
.B(n_509),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_505),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_526),
.A2(n_521),
.B(n_520),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_2),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_522),
.C(n_527),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_530),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_2),
.B(n_4),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_535),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_503),
.C(n_514),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_SL g536 ( 
.A1(n_519),
.A2(n_512),
.B(n_4),
.C(n_7),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_SL g537 ( 
.A1(n_536),
.A2(n_11),
.B(n_4),
.C(n_7),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_541),
.B(n_8),
.Y(n_544)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_533),
.C(n_9),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_2),
.C(n_8),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_539),
.B(n_533),
.C(n_9),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_542),
.A2(n_538),
.B(n_9),
.Y(n_545)
);

AO21x1_ASAP7_75t_L g546 ( 
.A1(n_543),
.A2(n_544),
.B(n_8),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_545),
.B(n_546),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_547),
.A2(n_11),
.B(n_9),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_10),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_10),
.B(n_11),
.Y(n_550)
);


endmodule