module fake_ariane_1299_n_166 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_166);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_166;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_156;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_121;
wire n_118;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

INVxp33_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_1),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_5),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_7),
.B1(n_8),
.B2(n_16),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_42),
.B1(n_46),
.B2(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_42),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_52),
.B1(n_62),
.B2(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_60),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_58),
.Y(n_92)
);

NAND2x1p5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_89),
.B(n_95),
.C(n_81),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_76),
.B(n_55),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_79),
.Y(n_102)
);

HB1xp67_ASAP7_75t_SL g103 ( 
.A(n_89),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_80),
.B(n_56),
.C(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_97),
.B(n_94),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_90),
.B1(n_83),
.B2(n_81),
.C(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_100),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_99),
.B(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_83),
.B1(n_90),
.B2(n_89),
.Y(n_111)
);

AND4x1_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_84),
.C(n_50),
.D(n_92),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_111),
.Y(n_117)
);

AO21x2_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_104),
.B(n_107),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_122),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_119),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_129),
.Y(n_142)
);

OAI221xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_121),
.B1(n_120),
.B2(n_50),
.C(n_56),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_135),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2x1_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_146),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_121),
.C(n_56),
.Y(n_151)
);

AND2x4_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_136),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_139),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_140),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_57),
.C(n_138),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_71),
.B(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_118),
.Y(n_157)
);

OR5x1_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_152),
.C(n_150),
.D(n_149),
.E(n_8),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_156),
.B(n_46),
.C(n_41),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_152),
.B(n_71),
.Y(n_160)
);

AOI211xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_155),
.B(n_61),
.C(n_53),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_84),
.B1(n_33),
.B2(n_93),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_159),
.Y(n_163)
);

NAND4xp25_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_96),
.C(n_106),
.D(n_18),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_17),
.Y(n_165)
);

AOI31xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_164),
.A3(n_106),
.B(n_107),
.Y(n_166)
);


endmodule