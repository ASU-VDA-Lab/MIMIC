module real_aes_571_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g590 ( .A(n_0), .B(n_245), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_1), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g168 ( .A(n_2), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_3), .B(n_527), .Y(n_526) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_4), .B(n_185), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_5), .B(n_229), .Y(n_237) );
INVx1_ASAP7_75t_L g575 ( .A(n_6), .Y(n_575) );
INVx1_ASAP7_75t_L g176 ( .A(n_7), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_8), .Y(n_116) );
AOI22xp5_ASAP7_75t_SL g134 ( .A1(n_9), .A2(n_135), .B1(n_136), .B2(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_9), .Y(n_135) );
OAI22x1_ASAP7_75t_R g137 ( .A1(n_10), .A2(n_79), .B1(n_138), .B2(n_139), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_10), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_11), .Y(n_202) );
AND2x2_ASAP7_75t_L g524 ( .A(n_12), .B(n_217), .Y(n_524) );
INVx2_ASAP7_75t_L g158 ( .A(n_13), .Y(n_158) );
AND3x1_ASAP7_75t_L g113 ( .A(n_14), .B(n_39), .C(n_114), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_14), .Y(n_128) );
INVx1_ASAP7_75t_L g246 ( .A(n_15), .Y(n_246) );
AOI221x1_ASAP7_75t_L g578 ( .A1(n_16), .A2(n_189), .B1(n_529), .B2(n_579), .C(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_17), .B(n_527), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_18), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g132 ( .A(n_18), .Y(n_132) );
INVx1_ASAP7_75t_L g243 ( .A(n_19), .Y(n_243) );
INVx1_ASAP7_75t_SL g258 ( .A(n_20), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_21), .B(n_179), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_22), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_23), .A2(n_30), .B1(n_515), .B2(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_23), .Y(n_843) );
AOI33xp33_ASAP7_75t_L g283 ( .A1(n_24), .A2(n_53), .A3(n_163), .B1(n_171), .B2(n_284), .B3(n_285), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_25), .A2(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_26), .B(n_245), .Y(n_531) );
AOI221xp5_ASAP7_75t_SL g554 ( .A1(n_27), .A2(n_44), .B1(n_527), .B2(n_529), .C(n_555), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_28), .A2(n_830), .B(n_845), .Y(n_829) );
INVx1_ASAP7_75t_L g848 ( .A(n_28), .Y(n_848) );
INVx1_ASAP7_75t_L g194 ( .A(n_29), .Y(n_194) );
NOR3xp33_ASAP7_75t_L g147 ( .A(n_30), .B(n_148), .C(n_339), .Y(n_147) );
INVx1_ASAP7_75t_SL g515 ( .A(n_30), .Y(n_515) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_31), .A2(n_91), .B(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g218 ( .A(n_31), .B(n_91), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_32), .B(n_248), .Y(n_566) );
INVxp67_ASAP7_75t_L g577 ( .A(n_33), .Y(n_577) );
AND2x2_ASAP7_75t_L g550 ( .A(n_34), .B(n_216), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_35), .B(n_169), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_36), .A2(n_529), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_37), .B(n_248), .Y(n_556) );
INVx1_ASAP7_75t_L g162 ( .A(n_38), .Y(n_162) );
AND2x2_ASAP7_75t_L g174 ( .A(n_38), .B(n_165), .Y(n_174) );
AND2x2_ASAP7_75t_L g185 ( .A(n_38), .B(n_168), .Y(n_185) );
OR2x6_ASAP7_75t_L g130 ( .A(n_39), .B(n_131), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_40), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_41), .B(n_169), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_42), .A2(n_190), .B1(n_225), .B2(n_229), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_43), .B(n_234), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_45), .A2(n_83), .B1(n_160), .B2(n_529), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_46), .B(n_179), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_47), .B(n_245), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_48), .B(n_156), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_49), .B(n_179), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_50), .Y(n_228) );
AND2x2_ASAP7_75t_L g593 ( .A(n_51), .B(n_216), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_52), .B(n_216), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_54), .B(n_179), .Y(n_214) );
INVx1_ASAP7_75t_L g167 ( .A(n_55), .Y(n_167) );
INVx1_ASAP7_75t_L g181 ( .A(n_55), .Y(n_181) );
AND2x2_ASAP7_75t_L g215 ( .A(n_56), .B(n_216), .Y(n_215) );
AOI221xp5_ASAP7_75t_L g159 ( .A1(n_57), .A2(n_75), .B1(n_160), .B2(n_169), .C(n_175), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_58), .B(n_169), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_59), .B(n_527), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_60), .B(n_190), .Y(n_204) );
AOI21xp5_ASAP7_75t_SL g267 ( .A1(n_61), .A2(n_160), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g541 ( .A(n_62), .B(n_216), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_63), .B(n_248), .Y(n_591) );
INVx1_ASAP7_75t_L g240 ( .A(n_64), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_65), .B(n_245), .Y(n_539) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_66), .B(n_217), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_67), .A2(n_529), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g213 ( .A(n_68), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_69), .B(n_248), .Y(n_532) );
AND2x2_ASAP7_75t_SL g605 ( .A(n_70), .B(n_156), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_71), .A2(n_160), .B(n_212), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_72), .A2(n_134), .B1(n_819), .B2(n_823), .Y(n_818) );
INVx1_ASAP7_75t_L g165 ( .A(n_73), .Y(n_165) );
INVx1_ASAP7_75t_L g183 ( .A(n_73), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_74), .B(n_169), .Y(n_286) );
AND2x2_ASAP7_75t_L g260 ( .A(n_76), .B(n_189), .Y(n_260) );
INVx1_ASAP7_75t_L g241 ( .A(n_77), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_78), .A2(n_160), .B(n_257), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_79), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_80), .A2(n_160), .B(n_231), .C(n_235), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_81), .B(n_527), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_82), .A2(n_86), .B1(n_169), .B2(n_527), .Y(n_603) );
INVx1_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_85), .B(n_189), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_87), .A2(n_160), .B1(n_281), .B2(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_88), .B(n_245), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_89), .B(n_245), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_90), .A2(n_529), .B(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_92), .Y(n_850) );
INVx1_ASAP7_75t_L g269 ( .A(n_93), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_94), .B(n_248), .Y(n_538) );
AND2x2_ASAP7_75t_L g287 ( .A(n_95), .B(n_189), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_96), .A2(n_192), .B(n_193), .C(n_196), .Y(n_191) );
INVxp67_ASAP7_75t_L g580 ( .A(n_97), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_98), .B(n_527), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_99), .B(n_248), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_100), .A2(n_529), .B(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_102), .B(n_179), .Y(n_270) );
OAI22xp5_ASAP7_75t_SL g840 ( .A1(n_103), .A2(n_841), .B1(n_842), .B2(n_844), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_103), .Y(n_841) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_117), .B(n_849), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_108), .Y(n_852) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_111), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_133), .B1(n_827), .B2(n_829), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
CKINVDCx11_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g828 ( .A(n_120), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp33_ASAP7_75t_L g845 ( .A1(n_124), .A2(n_846), .B(n_847), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g834 ( .A(n_127), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x6_ASAP7_75t_SL g145 ( .A(n_128), .B(n_130), .Y(n_145) );
OR2x6_ASAP7_75t_SL g817 ( .A(n_128), .B(n_129), .Y(n_817) );
OR2x2_ASAP7_75t_L g826 ( .A(n_128), .B(n_130), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_818), .Y(n_133) );
INVxp33_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B1(n_517), .B2(n_815), .Y(n_141) );
CKINVDCx6p67_ASAP7_75t_R g142 ( .A(n_143), .Y(n_142) );
CKINVDCx11_ASAP7_75t_R g822 ( .A(n_143), .Y(n_822) );
INVx3_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_145), .Y(n_144) );
AOI211xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_410), .B(n_513), .C(n_516), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_147), .A2(n_410), .B(n_513), .Y(n_820) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_149), .A2(n_411), .B(n_515), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_149), .B(n_488), .Y(n_838) );
NOR2x1_ASAP7_75t_L g149 ( .A(n_150), .B(n_317), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_300), .Y(n_150) );
AOI221xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_219), .B1(n_261), .B2(n_275), .C(n_290), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_206), .Y(n_152) );
NAND2x1_ASAP7_75t_SL g326 ( .A(n_153), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_153), .B(n_323), .Y(n_353) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_153), .Y(n_399) );
AND2x2_ASAP7_75t_L g407 ( .A(n_153), .B(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g511 ( .A(n_153), .Y(n_511) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_187), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_155), .Y(n_289) );
INVx1_ASAP7_75t_L g305 ( .A(n_155), .Y(n_305) );
AND2x4_ASAP7_75t_L g312 ( .A(n_155), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g322 ( .A(n_155), .B(n_187), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_155), .B(n_308), .Y(n_349) );
INVx1_ASAP7_75t_L g360 ( .A(n_155), .Y(n_360) );
INVxp67_ASAP7_75t_L g394 ( .A(n_155), .Y(n_394) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_186), .Y(n_155) );
INVx2_ASAP7_75t_SL g235 ( .A(n_156), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_156), .A2(n_562), .B(n_563), .Y(n_561) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_158), .B(n_218), .Y(n_217) );
AND2x4_ASAP7_75t_L g229 ( .A(n_158), .B(n_218), .Y(n_229) );
INVxp67_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_160), .A2(n_169), .B1(n_574), .B2(n_576), .Y(n_573) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_166), .Y(n_160) );
NOR2x1p5_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx1_ASAP7_75t_L g285 ( .A(n_163), .Y(n_285) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OR2x6_ASAP7_75t_L g177 ( .A(n_164), .B(n_171), .Y(n_177) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x6_ASAP7_75t_L g245 ( .A(n_165), .B(n_180), .Y(n_245) );
AND2x6_ASAP7_75t_L g529 ( .A(n_166), .B(n_174), .Y(n_529) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx2_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
AND2x4_ASAP7_75t_L g248 ( .A(n_167), .B(n_182), .Y(n_248) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_168), .Y(n_172) );
INVx1_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_173), .Y(n_169) );
INVx1_ASAP7_75t_L g226 ( .A(n_170), .Y(n_226) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVxp33_ASAP7_75t_L g284 ( .A(n_171), .Y(n_284) );
INVx1_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_184), .Y(n_175) );
INVxp67_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_177), .A2(n_184), .B(n_213), .C(n_214), .Y(n_212) );
INVx2_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_177), .A2(n_195), .B1(n_240), .B2(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_177), .A2(n_184), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_177), .A2(n_184), .B(n_269), .C(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g195 ( .A(n_179), .Y(n_195) );
AND2x4_ASAP7_75t_L g527 ( .A(n_179), .B(n_185), .Y(n_527) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_182), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_184), .A2(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_184), .B(n_229), .Y(n_249) );
INVx1_ASAP7_75t_L g281 ( .A(n_184), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_184), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_184), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_184), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_184), .A2(n_556), .B(n_557), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_184), .A2(n_565), .B(n_566), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_184), .A2(n_590), .B(n_591), .Y(n_589) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_185), .Y(n_196) );
INVx2_ASAP7_75t_L g277 ( .A(n_187), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_187), .B(n_208), .Y(n_293) );
INVx1_ASAP7_75t_L g311 ( .A(n_187), .Y(n_311) );
INVx1_ASAP7_75t_L g358 ( .A(n_187), .Y(n_358) );
OR2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_191), .B1(n_197), .B2(n_198), .Y(n_188) );
INVx3_ASAP7_75t_L g198 ( .A(n_189), .Y(n_198) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_190), .B(n_201), .Y(n_200) );
AOI21x1_ASAP7_75t_L g586 ( .A1(n_190), .A2(n_587), .B(n_593), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_195), .B(n_229), .C(n_582), .Y(n_581) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_198), .A2(n_209), .B(n_215), .Y(n_208) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_198), .A2(n_209), .B(n_215), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_199) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_206), .B(n_330), .Y(n_335) );
AND2x2_ASAP7_75t_L g347 ( .A(n_206), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g366 ( .A(n_206), .B(n_312), .Y(n_366) );
INVx1_ASAP7_75t_L g375 ( .A(n_206), .Y(n_375) );
AND2x2_ASAP7_75t_L g423 ( .A(n_206), .B(n_322), .Y(n_423) );
OR2x2_ASAP7_75t_L g466 ( .A(n_206), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g306 ( .A(n_207), .B(n_307), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_207), .B(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g288 ( .A(n_208), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_208), .B(n_308), .Y(n_386) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_208), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_216), .Y(n_253) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_216), .A2(n_554), .B(n_558), .Y(n_553) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_250), .Y(n_220) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_221), .B(n_345), .Y(n_390) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g352 ( .A(n_222), .B(n_343), .Y(n_352) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
INVx1_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
AND2x4_ASAP7_75t_L g298 ( .A(n_223), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g302 ( .A(n_223), .Y(n_302) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_223), .Y(n_338) );
AND2x2_ASAP7_75t_L g508 ( .A(n_223), .B(n_264), .Y(n_508) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
NOR3xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .C(n_228), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_229), .A2(n_267), .B(n_271), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_229), .A2(n_526), .B(n_528), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_229), .B(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_229), .B(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_229), .B(n_580), .Y(n_579) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_235), .A2(n_279), .B(n_287), .Y(n_278) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_235), .A2(n_279), .B(n_287), .Y(n_308) );
AOI21x1_ASAP7_75t_L g601 ( .A1(n_235), .A2(n_602), .B(n_605), .Y(n_601) );
INVx3_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
INVx2_ASAP7_75t_L g316 ( .A(n_236), .Y(n_316) );
NOR2x1_ASAP7_75t_SL g333 ( .A(n_236), .B(n_264), .Y(n_333) );
AND2x2_ASAP7_75t_L g371 ( .A(n_236), .B(n_252), .Y(n_371) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_242), .B(n_249), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B1(n_246), .B2(n_247), .Y(n_242) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g445 ( .A(n_250), .Y(n_445) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g274 ( .A(n_251), .Y(n_274) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
INVx1_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
INVx1_ASAP7_75t_L g403 ( .A(n_252), .Y(n_403) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_252), .Y(n_422) );
OR2x2_ASAP7_75t_L g428 ( .A(n_252), .B(n_264), .Y(n_428) );
AND2x2_ASAP7_75t_L g472 ( .A(n_252), .B(n_299), .Y(n_472) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_260), .Y(n_252) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_253), .A2(n_535), .B(n_541), .Y(n_534) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_253), .A2(n_544), .B(n_550), .Y(n_543) );
AO21x2_ASAP7_75t_L g682 ( .A1(n_253), .A2(n_544), .B(n_550), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_273), .Y(n_262) );
AND2x2_ASAP7_75t_L g314 ( .A(n_263), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g468 ( .A(n_263), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g473 ( .A(n_263), .Y(n_473) );
AND2x2_ASAP7_75t_L g485 ( .A(n_263), .B(n_371), .Y(n_485) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_272), .Y(n_263) );
INVx4_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
INVx2_ASAP7_75t_L g346 ( .A(n_264), .Y(n_346) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_264), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_264), .B(n_404), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_264), .B(n_274), .Y(n_477) );
AND2x2_ASAP7_75t_L g503 ( .A(n_264), .B(n_316), .Y(n_503) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x4_ASAP7_75t_L g405 ( .A(n_272), .B(n_296), .Y(n_405) );
AND2x2_ASAP7_75t_L g332 ( .A(n_273), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g350 ( .A(n_273), .B(n_337), .Y(n_350) );
INVx1_ASAP7_75t_L g384 ( .A(n_273), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_273), .B(n_298), .Y(n_440) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_274), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_275), .A2(n_357), .B1(n_501), .B2(n_504), .Y(n_500) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_288), .Y(n_275) );
INVx1_ASAP7_75t_L g430 ( .A(n_276), .Y(n_430) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g453 ( .A(n_277), .B(n_325), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g462 ( .A(n_277), .B(n_325), .Y(n_462) );
INVx2_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x4_ASAP7_75t_L g323 ( .A(n_278), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g327 ( .A(n_278), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_286), .Y(n_279) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_289), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_292), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g397 ( .A(n_292), .B(n_312), .Y(n_397) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g435 ( .A(n_293), .B(n_349), .Y(n_435) );
INVxp33_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g416 ( .A(n_295), .Y(n_416) );
NOR2x1_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_296), .B(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_296), .Y(n_362) );
INVx2_ASAP7_75t_L g426 ( .A(n_297), .Y(n_426) );
NAND2xp33_ASAP7_75t_SL g501 ( .A(n_297), .B(n_502), .Y(n_501) );
INVx4_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g367 ( .A(n_298), .B(n_346), .Y(n_367) );
AND2x2_ASAP7_75t_L g301 ( .A(n_299), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g404 ( .A(n_299), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B1(n_309), .B2(n_314), .Y(n_300) );
AND2x2_ASAP7_75t_L g329 ( .A(n_301), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g434 ( .A(n_301), .Y(n_434) );
INVx1_ASAP7_75t_L g383 ( .A(n_302), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_303), .A2(n_342), .B1(n_347), .B2(n_350), .Y(n_341) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx2_ASAP7_75t_L g467 ( .A(n_304), .Y(n_467) );
BUFx3_ASAP7_75t_L g432 ( .A(n_305), .Y(n_432) );
INVx1_ASAP7_75t_L g455 ( .A(n_306), .Y(n_455) );
AND2x2_ASAP7_75t_L g393 ( .A(n_307), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g460 ( .A(n_307), .B(n_325), .Y(n_460) );
INVx1_ASAP7_75t_L g494 ( .A(n_307), .Y(n_494) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI21xp33_ASAP7_75t_L g331 ( .A1(n_309), .A2(n_332), .B(n_334), .Y(n_331) );
OA21x2_ASAP7_75t_L g365 ( .A1(n_309), .A2(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g442 ( .A(n_311), .Y(n_442) );
AND2x2_ASAP7_75t_L g459 ( .A(n_311), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g449 ( .A(n_312), .B(n_408), .Y(n_449) );
AND2x2_ASAP7_75t_L g452 ( .A(n_312), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g461 ( .A(n_312), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g406 ( .A(n_315), .B(n_405), .Y(n_406) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_316), .B(n_345), .Y(n_344) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_316), .B(n_421), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_328), .B(n_331), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_326), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_321), .A2(n_337), .B1(n_362), .B2(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_325), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_327), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_327), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g469 ( .A(n_330), .Y(n_469) );
AND2x2_ASAP7_75t_L g456 ( .A(n_333), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_R g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_337), .B(n_420), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_339), .Y(n_514) );
OR3x2_ASAP7_75t_L g837 ( .A(n_339), .B(n_412), .C(n_838), .Y(n_837) );
NAND3x1_ASAP7_75t_SL g339 ( .A(n_340), .B(n_354), .C(n_368), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_351), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_342), .A2(n_452), .B1(n_454), .B2(n_456), .Y(n_451) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_343), .B(n_382), .Y(n_396) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_348), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g417 ( .A(n_348), .B(n_358), .Y(n_417) );
AND2x2_ASAP7_75t_L g441 ( .A(n_348), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_352), .A2(n_448), .B(n_449), .Y(n_447) );
AND2x2_ASAP7_75t_L g499 ( .A(n_352), .B(n_378), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_353), .A2(n_506), .B1(n_509), .B2(n_512), .Y(n_505) );
AOI21xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_361), .B(n_365), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
BUFx2_ASAP7_75t_L g475 ( .A(n_358), .Y(n_475) );
INVx1_ASAP7_75t_SL g482 ( .A(n_358), .Y(n_482) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_359), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_388), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B(n_376), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g377 ( .A(n_371), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_371), .B(n_382), .Y(n_463) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_379), .B(n_385), .Y(n_376) );
OR2x6_ASAP7_75t_L g433 ( .A(n_378), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g483 ( .A(n_386), .Y(n_483) );
OR2x2_ASAP7_75t_L g510 ( .A(n_386), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_387), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_398), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_395), .B2(n_397), .Y(n_389) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_392), .Y(n_490) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_406), .B2(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
AND2x4_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_486), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_436), .C(n_464), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_424), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_418), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp33_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_429), .B1(n_433), .B2(n_435), .Y(n_424) );
NAND2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_426), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_428), .B(n_434), .Y(n_504) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx3_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
INVx2_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_450), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_447), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_441), .B1(n_443), .B2(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_446), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_458), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_453), .B(n_494), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g478 ( .A(n_461), .Y(n_478) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B(n_470), .C(n_479), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI211xp5_ASAP7_75t_L g497 ( .A1(n_467), .A2(n_498), .B(n_500), .C(n_505), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_474), .B1(n_476), .B2(n_478), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_SL g513 ( .A1(n_486), .A2(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp67_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .Y(n_488) );
AOI21xp33_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B(n_495), .Y(n_489) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVxp33_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_516), .B(n_822), .Y(n_821) );
AO22x2_ASAP7_75t_L g819 ( .A1(n_517), .A2(n_816), .B1(n_820), .B2(n_821), .Y(n_819) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_726), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_648), .C(n_698), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_615), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_551), .B1(n_568), .B2(n_598), .C(n_607), .Y(n_521) );
INVx1_ASAP7_75t_SL g697 ( .A(n_522), .Y(n_697) );
AND2x4_ASAP7_75t_SL g522 ( .A(n_523), .B(n_533), .Y(n_522) );
INVx2_ASAP7_75t_L g619 ( .A(n_523), .Y(n_619) );
OR2x2_ASAP7_75t_L g641 ( .A(n_523), .B(n_632), .Y(n_641) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_523), .Y(n_656) );
INVx5_ASAP7_75t_L g663 ( .A(n_523), .Y(n_663) );
AND2x4_ASAP7_75t_L g669 ( .A(n_523), .B(n_543), .Y(n_669) );
AND2x2_ASAP7_75t_SL g672 ( .A(n_523), .B(n_600), .Y(n_672) );
OR2x2_ASAP7_75t_L g681 ( .A(n_523), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g688 ( .A(n_523), .B(n_534), .Y(n_688) );
AND2x2_ASAP7_75t_L g789 ( .A(n_523), .B(n_542), .Y(n_789) );
OR2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx3_ASAP7_75t_SL g640 ( .A(n_533), .Y(n_640) );
AND2x2_ASAP7_75t_L g684 ( .A(n_533), .B(n_600), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_533), .A2(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g725 ( .A(n_533), .B(n_663), .Y(n_725) );
AND2x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_542), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_534), .B(n_543), .Y(n_606) );
OR2x2_ASAP7_75t_L g610 ( .A(n_534), .B(n_543), .Y(n_610) );
INVx1_ASAP7_75t_L g618 ( .A(n_534), .Y(n_618) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_534), .Y(n_630) );
INVx2_ASAP7_75t_L g638 ( .A(n_534), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_534), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g747 ( .A(n_534), .B(n_632), .Y(n_747) );
AND2x2_ASAP7_75t_L g762 ( .A(n_534), .B(n_600), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_540), .Y(n_535) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g631 ( .A(n_543), .B(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_543), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_551), .B(n_755), .Y(n_754) );
NOR2x1p5_ASAP7_75t_L g551 ( .A(n_552), .B(n_559), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g584 ( .A(n_553), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_553), .B(n_560), .Y(n_613) );
INVx1_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
INVx2_ASAP7_75t_L g646 ( .A(n_553), .Y(n_646) );
INVx2_ASAP7_75t_L g652 ( .A(n_553), .Y(n_652) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_553), .Y(n_722) );
OR2x2_ASAP7_75t_L g753 ( .A(n_553), .B(n_560), .Y(n_753) );
OR2x2_ASAP7_75t_L g769 ( .A(n_559), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_SL g571 ( .A(n_560), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g596 ( .A(n_560), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g633 ( .A(n_560), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g645 ( .A(n_560), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g658 ( .A(n_560), .B(n_624), .Y(n_658) );
OR2x2_ASAP7_75t_L g666 ( .A(n_560), .B(n_572), .Y(n_666) );
INVx2_ASAP7_75t_L g693 ( .A(n_560), .Y(n_693) );
INVx1_ASAP7_75t_L g711 ( .A(n_560), .Y(n_711) );
NOR2xp33_ASAP7_75t_R g744 ( .A(n_560), .B(n_585), .Y(n_744) );
OR2x6_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_594), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_569), .A2(n_636), .B1(n_639), .B2(n_642), .Y(n_635) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_583), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g650 ( .A(n_571), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g685 ( .A(n_571), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g764 ( .A(n_571), .B(n_742), .Y(n_764) );
INVx3_ASAP7_75t_L g597 ( .A(n_572), .Y(n_597) );
AND2x4_ASAP7_75t_L g624 ( .A(n_572), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_572), .B(n_585), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_572), .B(n_646), .Y(n_691) );
AND2x2_ASAP7_75t_L g696 ( .A(n_572), .B(n_693), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_572), .B(n_584), .Y(n_733) );
INVx1_ASAP7_75t_L g803 ( .A(n_572), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_572), .B(n_721), .Y(n_814) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g595 ( .A(n_585), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_585), .B(n_597), .Y(n_614) );
INVx2_ASAP7_75t_L g625 ( .A(n_585), .Y(n_625) );
AND2x2_ASAP7_75t_L g651 ( .A(n_585), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g667 ( .A(n_585), .B(n_646), .Y(n_667) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_585), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_585), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g756 ( .A(n_585), .Y(n_756) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_595), .B(n_623), .Y(n_634) );
AOI221x1_ASAP7_75t_SL g728 ( .A1(n_596), .A2(n_729), .B1(n_732), .B2(n_734), .C(n_738), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_596), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g786 ( .A(n_596), .B(n_651), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_596), .B(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_L g717 ( .A(n_597), .B(n_645), .Y(n_717) );
AND2x2_ASAP7_75t_L g755 ( .A(n_597), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_606), .Y(n_599) );
AND2x2_ASAP7_75t_L g608 ( .A(n_600), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g703 ( .A(n_600), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_600), .B(n_619), .Y(n_708) );
AND2x4_ASAP7_75t_L g737 ( .A(n_600), .B(n_638), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_600), .B(n_669), .Y(n_773) );
OR2x2_ASAP7_75t_L g791 ( .A(n_600), .B(n_722), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_600), .B(n_682), .Y(n_801) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g632 ( .A(n_601), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g657 ( .A(n_606), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_606), .A2(n_665), .B1(n_668), .B2(n_670), .Y(n_664) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVx2_ASAP7_75t_L g620 ( .A(n_608), .Y(n_620) );
AND2x2_ASAP7_75t_L g759 ( .A(n_609), .B(n_619), .Y(n_759) );
AND2x2_ASAP7_75t_L g805 ( .A(n_609), .B(n_672), .Y(n_805) );
AND2x2_ASAP7_75t_L g810 ( .A(n_609), .B(n_661), .Y(n_810) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI32xp33_ASAP7_75t_L g779 ( .A1(n_611), .A2(n_681), .A3(n_761), .B1(n_780), .B2(n_782), .Y(n_779) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
AOI211xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_621), .B(n_626), .C(n_635), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_618), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_619), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g799 ( .A(n_619), .Y(n_799) );
AND2x2_ASAP7_75t_L g709 ( .A(n_621), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_622), .B(n_624), .Y(n_621) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_622), .Y(n_809) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_623), .Y(n_678) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_623), .Y(n_778) );
INVx1_ASAP7_75t_L g675 ( .A(n_624), .Y(n_675) );
AND2x2_ASAP7_75t_L g741 ( .A(n_624), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_624), .B(n_752), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_628), .A2(n_708), .B(n_709), .Y(n_707) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g637 ( .A(n_632), .B(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_L g661 ( .A(n_632), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_637), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g768 ( .A(n_637), .Y(n_768) );
AND2x2_ASAP7_75t_L g798 ( .A(n_637), .B(n_799), .Y(n_798) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_638), .Y(n_775) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_640), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g715 ( .A(n_641), .Y(n_715) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g674 ( .A(n_645), .B(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_646), .Y(n_742) );
AND2x2_ASAP7_75t_L g751 ( .A(n_647), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_671), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_658), .B2(n_659), .C(n_664), .Y(n_649) );
INVx1_ASAP7_75t_L g770 ( .A(n_651), .Y(n_770) );
INVxp33_ASAP7_75t_SL g802 ( .A(n_651), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_653), .A2(n_749), .B(n_757), .Y(n_748) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_657), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g670 ( .A(n_658), .Y(n_670) );
AND2x2_ASAP7_75t_L g705 ( .A(n_658), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g724 ( .A(n_658), .B(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_658), .A2(n_786), .B1(n_787), .B2(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OR2x2_ASAP7_75t_L g680 ( .A(n_661), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_661), .B(n_669), .Y(n_719) );
AND2x4_ASAP7_75t_L g736 ( .A(n_663), .B(n_682), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_663), .B(n_737), .Y(n_783) );
AND2x2_ASAP7_75t_L g795 ( .A(n_663), .B(n_747), .Y(n_795) );
NAND2xp33_ASAP7_75t_L g780 ( .A(n_665), .B(n_781), .Y(n_780) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_SL g723 ( .A(n_666), .Y(n_723) );
INVx1_ASAP7_75t_L g794 ( .A(n_667), .Y(n_794) );
INVx2_ASAP7_75t_SL g746 ( .A(n_669), .Y(n_746) );
AOI211xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_673), .B(n_676), .C(n_694), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B(n_683), .C(n_687), .Y(n_676) );
OR2x6_ASAP7_75t_SL g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g706 ( .A(n_678), .Y(n_706) );
INVx1_ASAP7_75t_SL g731 ( .A(n_681), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_681), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_686), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g772 ( .A1(n_690), .A2(n_773), .B1(n_774), .B2(n_776), .Y(n_772) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_704), .B(n_707), .C(n_712), .Y(n_698) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .B1(n_718), .B2(n_720), .C(n_724), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g804 ( .A1(n_723), .A2(n_805), .B1(n_806), .B2(n_810), .C1(n_811), .C2(n_813), .Y(n_804) );
INVx2_ASAP7_75t_L g739 ( .A(n_725), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_765), .C(n_784), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_748), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_736), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_737), .B(n_799), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_743), .B2(n_745), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVxp33_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_746), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_754), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_754), .A2(n_758), .B1(n_760), .B2(n_763), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
CKINVDCx16_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
OAI211xp5_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_769), .B(n_771), .C(n_779), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVxp67_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_792), .C(n_804), .Y(n_784) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI21xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_796), .B(n_803), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_800), .B(n_802), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
INVx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_835), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_832), .B(n_848), .Y(n_847) );
BUFx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_834), .Y(n_833) );
INVxp67_ASAP7_75t_L g846 ( .A(n_835), .Y(n_846) );
AOI22x1_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B1(n_839), .B2(n_840), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g844 ( .A(n_842), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_852), .Y(n_851) );
endmodule