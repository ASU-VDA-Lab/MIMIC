module fake_jpeg_25628_n_204 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_11),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_13),
.B1(n_20),
.B2(n_15),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_33),
.B1(n_24),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_13),
.B1(n_20),
.B2(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_38),
.B1(n_42),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_22),
.B1(n_18),
.B2(n_12),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_20),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_23),
.A2(n_18),
.B1(n_12),
.B2(n_17),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_42),
.B(n_38),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_24),
.B1(n_28),
.B2(n_30),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_50),
.B1(n_53),
.B2(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_29),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx2_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_56),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_11),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_0),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_53),
.B1(n_63),
.B2(n_69),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_54),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_72),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_35),
.B(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_57),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_33),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_35),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_43),
.C(n_44),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_82),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_46),
.B1(n_45),
.B2(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_43),
.B1(n_47),
.B2(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_72),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_44),
.B1(n_55),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_55),
.B1(n_50),
.B2(n_44),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_73),
.B1(n_59),
.B2(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_102),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_73),
.B(n_64),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_77),
.B(n_74),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_80),
.B1(n_81),
.B2(n_76),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_67),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_98),
.C(n_100),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_102),
.C(n_96),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_48),
.B1(n_58),
.B2(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_18),
.B(n_12),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_116),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_93),
.C(n_90),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_60),
.B(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_83),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_95),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_87),
.B1(n_83),
.B2(n_75),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_128),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_131),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_95),
.C(n_96),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_117),
.C(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_51),
.B1(n_34),
.B2(n_40),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_51),
.B1(n_34),
.B2(n_36),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_134),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_133),
.B(n_108),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_17),
.B(n_14),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_17),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_34),
.B1(n_36),
.B2(n_11),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_118),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_111),
.C(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_148),
.Y(n_156)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_147),
.B1(n_109),
.B2(n_124),
.Y(n_155)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_113),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_113),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_110),
.B(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_110),
.C(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_150),
.A2(n_136),
.B1(n_126),
.B2(n_124),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_153),
.C(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_157),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_125),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_131),
.B1(n_121),
.B2(n_133),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_138),
.B1(n_150),
.B2(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_134),
.B1(n_34),
.B2(n_41),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_10),
.B1(n_41),
.B2(n_2),
.Y(n_161)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_10),
.B1(n_17),
.B2(n_14),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_0),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_151),
.C(n_145),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_166),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_151),
.C(n_137),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_41),
.B(n_1),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_174),
.B(n_168),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_0),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_173),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_157),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_2),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_3),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_158),
.Y(n_180)
);

XNOR2x2_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_4),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_182),
.B(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_160),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_164),
.B(n_5),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_165),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_170),
.B(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_6),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_4),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_190),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_187),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_182),
.C(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_191),
.C(n_7),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_6),
.C(n_8),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_196),
.Y(n_202)
);

AOI221xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_8),
.B1(n_9),
.B2(n_199),
.C(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_8),
.Y(n_204)
);


endmodule