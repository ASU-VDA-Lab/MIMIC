module fake_jpeg_13346_n_612 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_612);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_612;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_585;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_1),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_65),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_23),
.B(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_27),
.Y(n_70)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_10),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_9),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_79),
.A2(n_35),
.B1(n_28),
.B2(n_21),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_85),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_86),
.B(n_109),
.Y(n_180)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_27),
.B(n_47),
.CON(n_100),
.SN(n_100)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_100),
.A2(n_13),
.B(n_18),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

BUFx2_ASAP7_75t_SL g215 ( 
.A(n_106),
.Y(n_215)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_20),
.B(n_9),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_110),
.B(n_112),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_20),
.B(n_30),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_120),
.Y(n_199)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_54),
.Y(n_204)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_79),
.B1(n_65),
.B2(n_60),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_134),
.A2(n_136),
.B1(n_158),
.B2(n_174),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_59),
.B(n_57),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_152),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_63),
.B(n_57),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_76),
.B(n_24),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_153),
.B(n_161),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_77),
.A2(n_90),
.B1(n_122),
.B2(n_75),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_154),
.A2(n_194),
.B1(n_195),
.B2(n_106),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_85),
.B(n_53),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_155),
.B(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_62),
.B(n_30),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_162),
.A2(n_190),
.B1(n_26),
.B2(n_6),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_109),
.B(n_44),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_164),
.B(n_170),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_96),
.B(n_44),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_85),
.B(n_33),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_103),
.B(n_33),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_189),
.B(n_206),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_66),
.A2(n_45),
.B1(n_56),
.B2(n_51),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_91),
.B(n_53),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_6),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_68),
.A2(n_41),
.B1(n_51),
.B2(n_48),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_80),
.A2(n_42),
.B1(n_35),
.B2(n_28),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_78),
.A2(n_93),
.B1(n_84),
.B2(n_88),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_200),
.B1(n_125),
.B2(n_89),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_113),
.A2(n_54),
.B1(n_48),
.B2(n_42),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_21),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_6),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_111),
.B(n_99),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_102),
.B(n_11),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_208),
.B(n_3),
.Y(n_286)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

BUFx2_ASAP7_75t_R g210 ( 
.A(n_91),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_216),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_70),
.B(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_SL g298 ( 
.A1(n_221),
.A2(n_249),
.B(n_272),
.C(n_294),
.Y(n_298)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_224),
.A2(n_285),
.B1(n_247),
.B2(n_239),
.Y(n_304)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_129),
.B(n_26),
.C(n_13),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_226),
.B(n_292),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_233),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_230),
.A2(n_252),
.B(n_254),
.Y(n_301)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_159),
.Y(n_232)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_232),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_234),
.B(n_276),
.Y(n_313)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_236),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_199),
.B1(n_134),
.B2(n_216),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_237),
.A2(n_245),
.B1(n_269),
.B2(n_273),
.Y(n_310)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

INVx3_ASAP7_75t_SL g308 ( 
.A(n_238),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_171),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_241),
.B(n_176),
.Y(n_326)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_134),
.A2(n_26),
.B1(n_6),
.B2(n_14),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_248),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_26),
.B1(n_14),
.B2(n_15),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_14),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_250),
.B(n_286),
.Y(n_316)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_132),
.B(n_0),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_0),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_293),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_132),
.B(n_204),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_145),
.Y(n_256)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_184),
.Y(n_259)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_142),
.Y(n_262)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_262),
.Y(n_348)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_169),
.Y(n_267)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_268),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_190),
.A2(n_213),
.B1(n_185),
.B2(n_177),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_178),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_271),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_182),
.B(n_0),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_168),
.A2(n_26),
.B1(n_14),
.B2(n_5),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_198),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_144),
.B(n_1),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_274),
.A2(n_281),
.B(n_290),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_142),
.A2(n_15),
.B1(n_17),
.B2(n_2),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_279),
.B1(n_240),
.B2(n_273),
.Y(n_307)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_149),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_278),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_179),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_160),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_144),
.B(n_3),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_283),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_152),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_200),
.A2(n_3),
.B1(n_141),
.B2(n_197),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_288),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_166),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_186),
.B(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_289),
.B(n_291),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_140),
.B(n_207),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_130),
.B(n_137),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_138),
.B(n_143),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_151),
.A2(n_183),
.B1(n_173),
.B2(n_157),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_256),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_299),
.B(n_311),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_304),
.A2(n_336),
.B1(n_338),
.B2(n_341),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_337),
.B1(n_347),
.B2(n_350),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_292),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_253),
.B(n_223),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_322),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_140),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_167),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_333),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_228),
.B(n_156),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_192),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_224),
.A2(n_192),
.B1(n_160),
.B2(n_171),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_245),
.A2(n_203),
.B1(n_150),
.B2(n_214),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_285),
.A2(n_203),
.B1(n_215),
.B2(n_175),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_290),
.A2(n_211),
.B1(n_292),
.B2(n_254),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_264),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_290),
.A2(n_279),
.B1(n_255),
.B2(n_294),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_254),
.A2(n_220),
.B1(n_226),
.B2(n_244),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_281),
.B(n_231),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_305),
.B(n_252),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_354),
.B(n_355),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_305),
.B(n_299),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_239),
.B(n_312),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_357),
.A2(n_364),
.B(n_339),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_304),
.A2(n_242),
.B1(n_268),
.B2(n_270),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_375),
.B1(n_377),
.B2(n_393),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_373),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_330),
.A2(n_239),
.B(n_252),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_350),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_376),
.C(n_380),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_314),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_368),
.B(n_372),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_310),
.A2(n_347),
.B1(n_307),
.B2(n_337),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_381),
.B1(n_385),
.B2(n_395),
.Y(n_400)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_315),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_302),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_295),
.A2(n_256),
.B1(n_232),
.B2(n_235),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_227),
.C(n_278),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_257),
.B1(n_238),
.B2(n_284),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_378),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_331),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_343),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_318),
.B(n_225),
.C(n_271),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_310),
.A2(n_271),
.B1(n_261),
.B2(n_265),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_219),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_389),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_266),
.C(n_236),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_334),
.C(n_309),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_301),
.A2(n_222),
.B1(n_258),
.B2(n_259),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_302),
.B(n_287),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_386),
.A2(n_388),
.B(n_319),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_322),
.A2(n_246),
.B1(n_251),
.B2(n_288),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_302),
.B(n_276),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_390),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_340),
.B(n_262),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_394),
.Y(n_410)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_392),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_338),
.A2(n_277),
.B1(n_282),
.B2(n_328),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_316),
.B(n_326),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_317),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_329),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_397),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_SL g397 ( 
.A(n_298),
.B(n_329),
.C(n_306),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_399),
.A2(n_373),
.B(n_361),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_298),
.B(n_339),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_401),
.A2(n_368),
.B(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_402),
.B(n_429),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_335),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_406),
.C(n_428),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_335),
.C(n_346),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_370),
.A2(n_298),
.B1(n_297),
.B2(n_308),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_411),
.A2(n_422),
.B1(n_423),
.B2(n_433),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_369),
.A2(n_359),
.B1(n_361),
.B2(n_360),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_413),
.A2(n_415),
.B1(n_388),
.B2(n_385),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_298),
.B1(n_308),
.B2(n_300),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_395),
.A2(n_319),
.B(n_343),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_416),
.A2(n_432),
.B(n_389),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_417),
.B(n_427),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_396),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_427),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_355),
.B(n_345),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_420),
.B(n_425),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_359),
.A2(n_308),
.B1(n_317),
.B2(n_323),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_381),
.A2(n_323),
.B1(n_348),
.B2(n_349),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_345),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_382),
.B(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_358),
.B(n_363),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_380),
.B(n_309),
.C(n_325),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_386),
.C(n_384),
.Y(n_447)
);

NAND2x1_ASAP7_75t_SL g432 ( 
.A(n_397),
.B(n_342),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_356),
.A2(n_323),
.B1(n_348),
.B2(n_349),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_362),
.B1(n_356),
.B2(n_372),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_436),
.A2(n_443),
.B(n_453),
.Y(n_478)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_437),
.Y(n_482)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_434),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_441),
.B(n_445),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_442),
.B(n_444),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_400),
.A2(n_373),
.B1(n_366),
.B2(n_393),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_410),
.B(n_394),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_433),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_413),
.A2(n_415),
.B1(n_432),
.B2(n_407),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_448),
.B1(n_449),
.B2(n_463),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_466),
.C(n_430),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_401),
.A2(n_357),
.B1(n_363),
.B2(n_391),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_405),
.Y(n_451)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_422),
.A2(n_379),
.B1(n_353),
.B2(n_365),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_452),
.A2(n_468),
.B1(n_408),
.B2(n_421),
.Y(n_473)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_456),
.A2(n_459),
.B(n_462),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_432),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_461),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_377),
.B1(n_375),
.B2(n_383),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_460),
.A2(n_405),
.B1(n_428),
.B2(n_414),
.Y(n_472)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_426),
.A2(n_364),
.B(n_371),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_407),
.A2(n_354),
.B1(n_387),
.B2(n_374),
.Y(n_463)
);

OAI211xp5_ASAP7_75t_L g464 ( 
.A1(n_426),
.A2(n_399),
.B(n_403),
.C(n_410),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_465),
.Y(n_494)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_404),
.B(n_398),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_423),
.A2(n_392),
.B1(n_390),
.B2(n_378),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_466),
.B(n_398),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_469),
.B(n_484),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_470),
.B(n_476),
.C(n_480),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_472),
.A2(n_473),
.B1(n_488),
.B2(n_489),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_442),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_487),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_406),
.C(n_424),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_424),
.C(n_425),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_467),
.B(n_420),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_483),
.B(n_449),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_424),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_468),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_443),
.A2(n_416),
.B1(n_421),
.B2(n_402),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_436),
.A2(n_408),
.B1(n_418),
.B2(n_365),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_458),
.A2(n_418),
.B1(n_342),
.B2(n_321),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_491),
.A2(n_448),
.B1(n_446),
.B2(n_437),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_447),
.B(n_325),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_469),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_327),
.C(n_303),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_495),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_467),
.B(n_462),
.C(n_450),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_451),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_463),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_445),
.B(n_327),
.Y(n_497)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_303),
.Y(n_498)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_475),
.Y(n_500)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_474),
.A2(n_460),
.B1(n_458),
.B2(n_452),
.Y(n_501)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_501),
.Y(n_531)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_477),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_510),
.Y(n_537)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_506),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_444),
.Y(n_509)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_481),
.Y(n_512)
);

OAI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_512),
.A2(n_514),
.B(n_520),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_498),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_515),
.B(n_516),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_519),
.A2(n_471),
.B1(n_487),
.B2(n_456),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_472),
.B(n_439),
.Y(n_521)
);

AOI21xp33_ASAP7_75t_L g534 ( 
.A1(n_521),
.A2(n_523),
.B(n_525),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_453),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_476),
.Y(n_532)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_482),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_480),
.B(n_484),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_526),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_471),
.A2(n_439),
.B1(n_450),
.B2(n_457),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_465),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_511),
.C(n_524),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_528),
.B(n_529),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_492),
.C(n_484),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_532),
.B(n_459),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_518),
.B(n_493),
.C(n_495),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_541),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_535),
.A2(n_488),
.B1(n_473),
.B2(n_520),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_499),
.C(n_483),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_513),
.B(n_499),
.C(n_483),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_543),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_506),
.A2(n_494),
.B(n_479),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_513),
.B(n_479),
.C(n_478),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_544),
.B(n_504),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_SL g546 ( 
.A(n_510),
.B(n_478),
.C(n_464),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_546),
.A2(n_497),
.B(n_517),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_519),
.Y(n_548)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_549),
.B(n_558),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_547),
.A2(n_531),
.B1(n_537),
.B2(n_507),
.Y(n_550)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_550),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_539),
.A2(n_500),
.B1(n_502),
.B2(n_505),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_553),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_505),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_537),
.A2(n_507),
.B1(n_538),
.B2(n_496),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_554),
.A2(n_535),
.B1(n_486),
.B2(n_491),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_522),
.C(n_515),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_555),
.B(n_557),
.Y(n_566)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_540),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_556),
.B(n_564),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_529),
.B(n_489),
.C(n_508),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_559),
.B(n_560),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_545),
.B(n_486),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_563),
.B(n_532),
.Y(n_578)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_562),
.B(n_534),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_568),
.B(n_575),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_569),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_545),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_573),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_554),
.A2(n_544),
.B1(n_543),
.B2(n_546),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_561),
.B(n_542),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_523),
.B1(n_512),
.B2(n_541),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_578),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_566),
.B(n_552),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_580),
.B(n_583),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_577),
.B(n_557),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_570),
.B(n_555),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_584),
.B(n_585),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_573),
.B(n_567),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_576),
.A2(n_572),
.B(n_565),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_586),
.A2(n_574),
.B(n_569),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_565),
.B(n_549),
.Y(n_587)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_587),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_558),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_548),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_592),
.A2(n_582),
.B(n_589),
.Y(n_599)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_588),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_593),
.B(n_594),
.Y(n_602)
);

BUFx24_ASAP7_75t_SL g595 ( 
.A(n_579),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g600 ( 
.A1(n_595),
.A2(n_581),
.B(n_553),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_528),
.Y(n_597)
);

INVxp33_ASAP7_75t_L g598 ( 
.A(n_597),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_599),
.A2(n_600),
.B(n_601),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_596),
.A2(n_581),
.B(n_551),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_591),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_590),
.C(n_594),
.Y(n_605)
);

AO21x1_ASAP7_75t_L g607 ( 
.A1(n_605),
.A2(n_553),
.B(n_485),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_598),
.A2(n_602),
.B(n_574),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_606),
.A2(n_530),
.B(n_485),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_607),
.B(n_608),
.C(n_482),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_609),
.B(n_604),
.C(n_435),
.Y(n_610)
);

AOI321xp33_ASAP7_75t_SL g611 ( 
.A1(n_610),
.A2(n_438),
.A3(n_454),
.B1(n_455),
.B2(n_461),
.C(n_530),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_321),
.Y(n_612)
);


endmodule