module fake_jpeg_14344_n_53 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_53);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_16),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_0),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_29),
.Y(n_34)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_24),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_24),
.B(n_19),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_35),
.C(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_19),
.C(n_18),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_18),
.C(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_32),
.C(n_31),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.C(n_1),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_28),
.C(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_4),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_46),
.B(n_47),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_12),
.Y(n_46)
);

XOR2x1_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_3),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_44),
.C(n_6),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_5),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_49),
.B(n_6),
.Y(n_52)
);

AOI321xp33_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_44),
.A3(n_7),
.B1(n_5),
.B2(n_13),
.C(n_17),
.Y(n_53)
);


endmodule