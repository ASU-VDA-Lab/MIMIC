module real_jpeg_12367_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_296, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_296;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_249;
wire n_292;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_52),
.B1(n_59),
.B2(n_62),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_6),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_6),
.A2(n_59),
.B1(n_62),
.B2(n_148),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_148),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_7),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_7),
.B(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_7),
.B(n_62),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_7),
.A2(n_64),
.B(n_187),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_140),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_7),
.A2(n_43),
.B(n_48),
.C(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_7),
.B(n_109),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_7),
.B(n_32),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_7),
.B(n_53),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_7),
.A2(n_62),
.B(n_178),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_9),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_70),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_10),
.A2(n_45),
.B1(n_59),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_10),
.A2(n_45),
.B1(n_64),
.B2(n_65),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_12),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_12),
.A2(n_59),
.B1(n_62),
.B2(n_101),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_101),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_101),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_68),
.Y(n_215)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_15),
.A2(n_36),
.B1(n_59),
.B2(n_62),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_16),
.A2(n_59),
.B1(n_62),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_16),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_16),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_78),
.Y(n_168)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_271),
.B1(n_293),
.B2(n_294),
.Y(n_19)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_124),
.B(n_270),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_22),
.B(n_102),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_86),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_23),
.B(n_80),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_28),
.A2(n_32),
.B(n_37),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_28),
.A2(n_32),
.B1(n_92),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_28),
.A2(n_32),
.B1(n_136),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_32),
.B1(n_168),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_28),
.A2(n_32),
.B1(n_181),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_28),
.A2(n_32),
.B1(n_140),
.B2(n_227),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_28),
.A2(n_32),
.B1(n_220),
.B2(n_227),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_29),
.B(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_31),
.A2(n_34),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_31),
.A2(n_90),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_35),
.A2(n_49),
.B(n_140),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_50),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_44),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_43),
.B(n_75),
.Y(n_179)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_44),
.A2(n_62),
.A3(n_74),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_46),
.A2(n_53),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_46),
.A2(n_53),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_46),
.A2(n_53),
.B1(n_95),
.B2(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_46),
.A2(n_53),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_46),
.A2(n_53),
.B1(n_206),
.B2(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_46),
.A2(n_53),
.B(n_111),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_50),
.A2(n_96),
.B1(n_171),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_57),
.A2(n_58),
.B1(n_147),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_57),
.A2(n_58),
.B1(n_120),
.B2(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_62),
.Y(n_138)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_65),
.B(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_72),
.A2(n_76),
.B1(n_143),
.B2(n_164),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_72),
.A2(n_76),
.B1(n_162),
.B2(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_82),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_82),
.A2(n_119),
.B(n_121),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_88),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_89),
.B(n_93),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_123),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B(n_112),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_109),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_109),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_112),
.A2(n_277),
.B1(n_289),
.B2(n_290),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_112),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_291)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_154),
.B(n_269),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_152),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_126),
.B(n_152),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_132),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_131),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_132),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.C(n_145),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_133),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_139),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_141),
.B(n_145),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI221xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_262),
.B1(n_267),
.B2(n_268),
.C(n_296),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_254),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_198),
.B(n_253),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_182),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_158),
.B(n_182),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.C(n_173),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_159),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_166),
.C(n_167),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_169),
.A2(n_173),
.B1(n_174),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_169),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_193),
.B2(n_197),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_194),
.C(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_185),
.B(n_189),
.C(n_192),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_247),
.B(n_252),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_236),
.B(n_246),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_216),
.B(n_235),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_202),
.B(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_212),
.C(n_214),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_234),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_222),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_233),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_242),
.C(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_292),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_291),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_291),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule