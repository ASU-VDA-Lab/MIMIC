module fake_jpeg_24762_n_267 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_22),
.B(n_26),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_58),
.B(n_34),
.C(n_29),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_14),
.Y(n_72)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_23),
.B1(n_14),
.B2(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_47),
.B1(n_38),
.B2(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_69),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_77),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_31),
.Y(n_75)
);

OR2x4_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_31),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_30),
.C(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g86 ( 
.A(n_80),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_16),
.CI(n_47),
.CON(n_81),
.SN(n_81)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_24),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_23),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_24),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_75),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_52),
.B1(n_42),
.B2(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_52),
.B1(n_15),
.B2(n_28),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_29),
.B1(n_16),
.B2(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_74),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_31),
.B1(n_16),
.B2(n_38),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_69),
.B1(n_43),
.B2(n_45),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_28),
.B1(n_16),
.B2(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_86),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_64),
.C(n_66),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_81),
.B(n_100),
.C(n_91),
.D(n_92),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_64),
.B(n_8),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_121),
.B(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_116),
.B(n_117),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_27),
.B1(n_19),
.B2(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_79),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_119),
.B(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_20),
.B(n_67),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_131),
.C(n_117),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_120),
.B1(n_116),
.B2(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_127),
.B(n_111),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_83),
.B1(n_81),
.B2(n_90),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_100),
.B1(n_93),
.B2(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_43),
.B1(n_57),
.B2(n_96),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_76),
.B1(n_99),
.B2(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_104),
.B1(n_105),
.B2(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_73),
.B1(n_27),
.B2(n_19),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_73),
.B(n_27),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_102),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_160),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_113),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_164),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_143),
.Y(n_163)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_110),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_125),
.C(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_8),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_137),
.B1(n_129),
.B2(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_147),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_184),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_131),
.C(n_127),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_130),
.C(n_139),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_142),
.B1(n_145),
.B2(n_137),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_175),
.A2(n_151),
.B1(n_152),
.B2(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_123),
.C(n_18),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_123),
.C(n_21),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_21),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_187),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_17),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_177),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_17),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_151),
.B1(n_153),
.B2(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_194),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_183),
.B1(n_174),
.B2(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_201),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_147),
.B1(n_166),
.B2(n_163),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_207),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_149),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_205),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_206),
.Y(n_226)
);

BUFx12f_ASAP7_75t_SL g209 ( 
.A(n_199),
.Y(n_209)
);

OAI21x1_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_222),
.B(n_7),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.C(n_0),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_173),
.C(n_17),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_6),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_6),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_5),
.Y(n_232)
);

NAND4xp25_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_6),
.C(n_12),
.D(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_192),
.B1(n_200),
.B2(n_190),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_228),
.B1(n_10),
.B2(n_13),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_233),
.C(n_212),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_235),
.B(n_218),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_12),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_1),
.C(n_2),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_9),
.B(n_12),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_235),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_243),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_232),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_220),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_233),
.B(n_234),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_237),
.B(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_251),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_13),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_13),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_1),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_245),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_250),
.B(n_2),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_256),
.A2(n_257),
.B(n_1),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_244),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_255),
.B1(n_252),
.B2(n_246),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_260),
.B(n_261),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_3),
.B(n_4),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_3),
.B(n_4),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_263),
.C(n_3),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_3),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_4),
.Y(n_267)
);


endmodule