module real_jpeg_2678_n_5 (n_4, n_0, n_1, n_2, n_30, n_28, n_29, n_3, n_31, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_30;
input n_28;
input n_29;
input n_3;
input n_31;

output n_5;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_0),
.A2(n_17),
.B(n_21),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g10 ( 
.A1(n_2),
.A2(n_11),
.B1(n_15),
.B2(n_26),
.Y(n_10)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_7),
.Y(n_6)
);

XNOR2xp5_ASAP7_75t_L g5 ( 
.A(n_6),
.B(n_10),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_9),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND3xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_24),
.C(n_25),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_28),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_29),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_30),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_31),
.Y(n_22)
);


endmodule