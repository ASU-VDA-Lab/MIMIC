module fake_jpeg_5872_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_3),
.Y(n_7)
);

MAJIxp5_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_3),
.C(n_2),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_22),
.B(n_23),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_21),
.B1(n_24),
.B2(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_13),
.B(n_5),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_10),
.B1(n_15),
.B2(n_8),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_11),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_14),
.B(n_12),
.Y(n_23)
);

AO22x1_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_13),
.B1(n_10),
.B2(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_16),
.B1(n_23),
.B2(n_11),
.Y(n_38)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

AND2x6_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_22),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_21),
.C(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_32),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.A3(n_38),
.B1(n_37),
.B2(n_35),
.C1(n_39),
.C2(n_17),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_29),
.Y(n_45)
);

OAI221xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_40),
.B2(n_42),
.C(n_9),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_45),
.B(n_9),
.Y(n_47)
);


endmodule