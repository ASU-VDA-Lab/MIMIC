module real_jpeg_27230_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_244;
wire n_216;
wire n_133;
wire n_179;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_43),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_1),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_57),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_2),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_87)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_67),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_67),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_5),
.A2(n_10),
.B(n_63),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_26),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_6),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_81),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_81),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_10),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_99),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_10),
.B(n_41),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_41),
.B(n_45),
.C(n_180),
.D(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_72),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_25),
.B(n_193),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g221 ( 
.A1(n_10),
.A2(n_64),
.B(n_75),
.C(n_112),
.D(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_10),
.B(n_64),
.Y(n_222)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_21),
.B(n_113),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.C(n_88),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_22),
.B(n_82),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_55),
.C(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_24),
.B(n_39),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_25),
.A2(n_36),
.B1(n_37),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_25),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_25),
.A2(n_34),
.B(n_84),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_25),
.A2(n_34),
.B1(n_105),
.B2(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_25),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_25),
.B(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_26),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_26),
.B(n_46),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_31),
.A2(n_35),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_33),
.A2(n_42),
.A3(n_47),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_33),
.B(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_34),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_34),
.A2(n_200),
.B(n_208),
.Y(n_207)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_35),
.B(n_194),
.Y(n_193)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_36),
.B(n_99),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_40),
.A2(n_52),
.B(n_146),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_46),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_41),
.A2(n_63),
.A3(n_222),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_42),
.B(n_78),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_50),
.B1(n_52),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_44),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_45),
.A2(n_49),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_45),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_45),
.A2(n_49),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_52),
.B(n_148),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_52),
.A2(n_146),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_52),
.B(n_99),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_68),
.B2(n_69),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_58),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_62),
.B(n_99),
.C(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_60),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_61),
.B(n_95),
.Y(n_129)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_64),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_66),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_74),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_71),
.B1(n_108),
.B2(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_80),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_71),
.A2(n_74),
.B(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_72),
.A2(n_75),
.B1(n_110),
.B2(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_78),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_86),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_87),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_88),
.A2(n_89),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.C(n_106),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_91),
.B1(n_106),
.B2(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_93),
.B(n_99),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_103),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_133),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_132),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_172),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_158),
.B(n_171),
.Y(n_137)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_155),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_155),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.C(n_152),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_152),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_159),
.B(n_161),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_162),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_166),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.C(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_167),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_168),
.B(n_170),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_169),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_249),
.C(n_250),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_244),
.B(n_248),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_233),
.B(n_243),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_217),
.B(n_232),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_196),
.B(n_216),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_182),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_204),
.B(n_215),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_209),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_210),
.B(n_214),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_219),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_223),
.C(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_225),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);


endmodule