module fake_jpeg_10640_n_95 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_1),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_2),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_69),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_38),
.C(n_39),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_59),
.B(n_64),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_46),
.C(n_40),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_45),
.B1(n_44),
.B2(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_5),
.B1(n_6),
.B2(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_44),
.B1(n_33),
.B2(n_4),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_2),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_81),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_63),
.B1(n_62),
.B2(n_61),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_71),
.B(n_73),
.C(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_71),
.Y(n_86)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_80),
.A3(n_79),
.B1(n_70),
.B2(n_82),
.C(n_83),
.Y(n_87)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_76),
.B1(n_79),
.B2(n_65),
.C(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

AOI31xp67_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_11),
.A3(n_12),
.B(n_14),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_15),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_16),
.B(n_17),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_19),
.B(n_20),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_24),
.B(n_27),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_28),
.Y(n_95)
);


endmodule