module fake_jpeg_8949_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_25),
.B1(n_32),
.B2(n_29),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_27),
.B1(n_28),
.B2(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_28),
.B1(n_27),
.B2(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_33),
.B(n_30),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_70),
.A2(n_83),
.B1(n_90),
.B2(n_92),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_17),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_89),
.B(n_91),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_88),
.B1(n_25),
.B2(n_26),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_22),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_38),
.B(n_39),
.C(n_45),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_95),
.A3(n_36),
.B1(n_47),
.B2(n_44),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_26),
.B1(n_24),
.B2(n_43),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_43),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_38),
.B1(n_45),
.B2(n_43),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_49),
.B1(n_42),
.B2(n_33),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_24),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_68),
.B1(n_66),
.B2(n_45),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_113),
.B1(n_117),
.B2(n_82),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_91),
.B(n_44),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_105),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_43),
.B1(n_52),
.B2(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_36),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_47),
.B1(n_67),
.B2(n_62),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_69),
.B1(n_49),
.B2(n_36),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_124),
.B1(n_73),
.B2(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_60),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_88),
.B1(n_94),
.B2(n_24),
.Y(n_129)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_130),
.B1(n_136),
.B2(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_113),
.B1(n_100),
.B2(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_138),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_85),
.B1(n_95),
.B2(n_77),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_82),
.B1(n_79),
.B2(n_93),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_79),
.B1(n_84),
.B2(n_81),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_102),
.B1(n_119),
.B2(n_111),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_81),
.B1(n_73),
.B2(n_75),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_140),
.A2(n_156),
.B1(n_21),
.B2(n_19),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_120),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_146),
.B(n_31),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_148),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_106),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_153),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_106),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_44),
.B1(n_41),
.B2(n_33),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_125),
.B1(n_119),
.B2(n_123),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_163),
.B1(n_186),
.B2(n_127),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_172),
.B1(n_127),
.B2(n_19),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_71),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_104),
.B1(n_30),
.B2(n_106),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_99),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_171),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_44),
.B(n_23),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_179),
.B(n_31),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_177),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_131),
.B(n_30),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_19),
.B1(n_104),
.B2(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_178),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_141),
.B(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_23),
.B(n_21),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_21),
.C(n_23),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_31),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_143),
.B(n_132),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_137),
.B1(n_132),
.B2(n_128),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_19),
.Y(n_187)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_155),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_157),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_193),
.B(n_200),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_195),
.A2(n_196),
.B1(n_199),
.B2(n_209),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_21),
.B1(n_9),
.B2(n_16),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_21),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_21),
.A3(n_31),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_206),
.C(n_214),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_162),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_217),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_21),
.B1(n_8),
.B2(n_16),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_1),
.B(n_2),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_31),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_187),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_168),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_178),
.B1(n_174),
.B2(n_181),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_234),
.B1(n_236),
.B2(n_240),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_159),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_237),
.C(n_238),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_235),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_169),
.B1(n_159),
.B2(n_176),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_176),
.B1(n_189),
.B2(n_186),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_166),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_239),
.B(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_183),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_194),
.C(n_197),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_197),
.B1(n_191),
.B2(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_193),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_214),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_209),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_259),
.C(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_201),
.B1(n_203),
.B2(n_172),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_238),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_172),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.C(n_242),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_211),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_202),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_224),
.B(n_223),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_278),
.B(n_280),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_220),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_170),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_267),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_283),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_248),
.A2(n_244),
.B(n_203),
.C(n_220),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_12),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_177),
.C(n_188),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_255),
.C(n_266),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_164),
.B1(n_212),
.B2(n_171),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_283),
.A2(n_284),
.B1(n_273),
.B2(n_276),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_264),
.B1(n_257),
.B2(n_247),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_262),
.B1(n_8),
.B2(n_11),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_278),
.B1(n_6),
.B2(n_14),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_258),
.B1(n_256),
.B2(n_259),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_296),
.B1(n_15),
.B2(n_4),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_294),
.C(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_293),
.B(n_286),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_7),
.C(n_14),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_7),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_15),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_12),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_5),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_12),
.C(n_14),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_278),
.B(n_13),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_15),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_307),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_312),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_286),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_2),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_5),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_300),
.B(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_305),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_290),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_330),
.C(n_320),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_303),
.B(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_310),
.C(n_4),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_325),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_322),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_331),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_318),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_5),
.Y(n_339)
);


endmodule