module fake_netlist_6_2826_n_2366 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2366);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2366;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_2127;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_2250;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_374;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_72),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_178),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_81),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_156),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_54),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_64),
.Y(n_243)
);

BUFx8_ASAP7_75t_SL g244 ( 
.A(n_93),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_139),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_82),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_68),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_85),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_146),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_24),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_193),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_215),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_70),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_150),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_218),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_53),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_226),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_168),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_55),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_123),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_92),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_30),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_51),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_129),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_23),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_38),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_107),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_66),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_67),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_24),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_143),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_144),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_66),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_135),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_195),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_103),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_115),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_5),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_44),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_203),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_106),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_192),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_59),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_59),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_211),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_75),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_174),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_148),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_142),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_2),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_4),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_145),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_113),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_122),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_95),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_172),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_61),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_87),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_48),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_154),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_177),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_190),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_88),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_67),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_65),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_201),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_53),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_126),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_158),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_82),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_216),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_56),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_22),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_175),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_222),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_19),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_58),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_77),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_220),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_93),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_104),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_161),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_85),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_57),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_104),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_33),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_224),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_11),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_69),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_165),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_95),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_65),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_57),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_44),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_151),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_99),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_42),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_204),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_114),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_64),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_181),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_14),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_10),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_69),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_147),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_6),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_125),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_176),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_217),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_17),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_112),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_58),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_23),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_4),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_111),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_138),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_12),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_43),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_131),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_89),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_121),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_92),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_70),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_109),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_52),
.Y(n_389)
);

BUFx8_ASAP7_75t_SL g390 ( 
.A(n_28),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_163),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_127),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_3),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_37),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_36),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_210),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_116),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_81),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_162),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_179),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_137),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_198),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_60),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_149),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_132),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_71),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_109),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_40),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_187),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_49),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_136),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_8),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_35),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_184),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_189),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_90),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_56),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_33),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_2),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_128),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_194),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_37),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_200),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_43),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_71),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_60),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_30),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_169),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_61),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_7),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_183),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_78),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_223),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_73),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_76),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_196),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_91),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_63),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_117),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_170),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_15),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_75),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_96),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_50),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_89),
.Y(n_445)
);

BUFx2_ASAP7_75t_SL g446 ( 
.A(n_96),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_40),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_171),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_94),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_38),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_3),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_155),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_111),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_90),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_231),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_249),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_244),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_247),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_270),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_249),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_355),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_355),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_355),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_343),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_331),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_355),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_343),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_290),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_369),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_390),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_0),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_R g472 ( 
.A(n_234),
.B(n_1),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_237),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_355),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_233),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_235),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_239),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_290),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_355),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_355),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_241),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_355),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_252),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_240),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_355),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_355),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_415),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_260),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_260),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_436),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_260),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_256),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_257),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_240),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_345),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_345),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_260),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_260),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_261),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_242),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_260),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_314),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_293),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_293),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_334),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_293),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_266),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_293),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_264),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_236),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_291),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_281),
.B(n_1),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_293),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_292),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_293),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_248),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_294),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_L g519 ( 
.A(n_281),
.B(n_6),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_305),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_267),
.B(n_7),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_307),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_443),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_266),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_310),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_236),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_282),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_311),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_315),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_245),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_316),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_318),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_322),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_290),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_236),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_328),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_400),
.B(n_8),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_330),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_282),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_273),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_337),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_273),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_338),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_353),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_358),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_254),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_266),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_364),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_383),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_273),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_296),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_385),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_391),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_296),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_396),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_296),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_400),
.B(n_9),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_344),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_404),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_344),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_344),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_348),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_258),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_411),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_414),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_348),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_348),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_420),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_349),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_349),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_421),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_349),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_473),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_489),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_521),
.B(n_471),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_478),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_485),
.B(n_251),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_484),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_456),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_460),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_493),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_521),
.B(n_324),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_494),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_506),
.B(n_243),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_467),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_462),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_455),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_500),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_489),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_512),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_515),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_503),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_492),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_498),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_479),
.B(n_539),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_498),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_503),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_499),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_499),
.Y(n_610)
);

INVxp33_ASAP7_75t_SL g611 ( 
.A(n_457),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_522),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_468),
.B(n_267),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_L g615 ( 
.A(n_552),
.B(n_287),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_502),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_511),
.B(n_373),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_458),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_531),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_504),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_504),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_505),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_505),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_507),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_532),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_535),
.B(n_423),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_536),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_507),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_552),
.B(n_287),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_538),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_543),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_462),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_542),
.B(n_562),
.C(n_519),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_468),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_514),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_548),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_511),
.B(n_373),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_514),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_483),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_516),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_550),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_553),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_483),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_508),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_554),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_516),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_523),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_485),
.B(n_251),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_557),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_508),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_R g659 ( 
.A(n_470),
.B(n_262),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_524),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_529),
.B(n_373),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_495),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_525),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_525),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_527),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_527),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_459),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_534),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_465),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_508),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_469),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_534),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_591),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_602),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_600),
.Y(n_678)
);

AND3x4_ASAP7_75t_L g679 ( 
.A(n_585),
.B(n_519),
.C(n_513),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_581),
.B(n_558),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_600),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_602),
.B(n_529),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_581),
.A2(n_588),
.B1(n_641),
.B2(n_606),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_588),
.B(n_569),
.Y(n_684)
);

AND3x4_ASAP7_75t_L g685 ( 
.A(n_585),
.B(n_513),
.C(n_336),
.Y(n_685)
);

AO22x2_ASAP7_75t_L g686 ( 
.A1(n_641),
.A2(n_243),
.B1(n_301),
.B2(n_287),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_623),
.B(n_570),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_602),
.B(n_537),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_623),
.B(n_510),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_642),
.B(n_537),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_618),
.B(n_301),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_606),
.B(n_518),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_646),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_642),
.Y(n_694)
);

BUFx8_ASAP7_75t_SL g695 ( 
.A(n_593),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_629),
.B(n_530),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_583),
.A2(n_528),
.B1(n_541),
.B2(n_520),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_R g698 ( 
.A(n_659),
.B(n_546),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_592),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_592),
.Y(n_700)
);

NAND3x1_ASAP7_75t_L g701 ( 
.A(n_606),
.B(n_253),
.C(n_245),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_642),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_646),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_600),
.Y(n_704)
);

AO22x2_ASAP7_75t_L g705 ( 
.A1(n_586),
.A2(n_350),
.B1(n_402),
.B2(n_301),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_592),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_618),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_598),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_SL g709 ( 
.A1(n_620),
.A2(n_308),
.B1(n_327),
.B2(n_274),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_618),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_645),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_579),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_598),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_583),
.B(n_501),
.C(n_482),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_582),
.B(n_549),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_651),
.Y(n_716)
);

BUFx4f_ASAP7_75t_L g717 ( 
.A(n_651),
.Y(n_717)
);

INVx6_ASAP7_75t_L g718 ( 
.A(n_608),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_645),
.B(n_540),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_584),
.B(n_560),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_645),
.B(n_540),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_587),
.B(n_306),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_580),
.Y(n_724)
);

AND2x6_ASAP7_75t_L g725 ( 
.A(n_663),
.B(n_350),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_595),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_598),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_595),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_596),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_663),
.B(n_614),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_596),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_601),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_601),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_603),
.Y(n_734)
);

NAND3x1_ASAP7_75t_L g735 ( 
.A(n_614),
.B(n_275),
.C(n_253),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_663),
.B(n_461),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_591),
.B(n_456),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_638),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_638),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_600),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_603),
.B(n_604),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_604),
.B(n_545),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_589),
.B(n_564),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_669),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_629),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_594),
.B(n_573),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_605),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_600),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_605),
.B(n_461),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_671),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_607),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

INVx6_ASAP7_75t_L g753 ( 
.A(n_608),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_656),
.A2(n_576),
.B1(n_497),
.B2(n_496),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_616),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_638),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_616),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_651),
.B(n_314),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_640),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_651),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_612),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_586),
.B(n_464),
.Y(n_764)
);

NOR2x1p5_ASAP7_75t_L g765 ( 
.A(n_597),
.B(n_306),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_599),
.B(n_530),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_607),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_609),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_673),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_651),
.B(n_324),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_609),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_612),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_610),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_640),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_610),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_617),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_640),
.B(n_350),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_664),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_615),
.B(n_545),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_617),
.B(n_547),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_656),
.B(n_544),
.Y(n_781)
);

XOR2xp5_ASAP7_75t_L g782 ( 
.A(n_664),
.B(n_474),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_619),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_619),
.B(n_463),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_613),
.B(n_544),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_621),
.B(n_464),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_622),
.B(n_463),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_402),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_616),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_590),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_622),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_628),
.B(n_517),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_630),
.A2(n_472),
.B1(n_280),
.B2(n_289),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_624),
.B(n_547),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_635),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_651),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_637),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_647),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_624),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_625),
.B(n_555),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_647),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_625),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_616),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_644),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_626),
.A2(n_382),
.B1(n_366),
.B2(n_336),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_626),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_649),
.B(n_551),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_665),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_616),
.Y(n_809)
);

NOR2x1p5_ASAP7_75t_L g810 ( 
.A(n_650),
.B(n_306),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_627),
.B(n_555),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_616),
.Y(n_812)
);

BUFx10_ASAP7_75t_L g813 ( 
.A(n_653),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_627),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_665),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_665),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_657),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_615),
.B(n_556),
.Y(n_818)
);

AND2x6_ASAP7_75t_L g819 ( 
.A(n_631),
.B(n_402),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_666),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_634),
.B(n_556),
.Y(n_821)
);

INVx6_ASAP7_75t_L g822 ( 
.A(n_608),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_611),
.B(n_568),
.Y(n_823)
);

INVx4_ASAP7_75t_SL g824 ( 
.A(n_616),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_666),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_631),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_636),
.B(n_639),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_636),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_639),
.B(n_466),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_643),
.B(n_466),
.Y(n_830)
);

INVx4_ASAP7_75t_SL g831 ( 
.A(n_632),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_643),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_648),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_648),
.B(n_533),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_654),
.B(n_488),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_724),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_707),
.B(n_314),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_730),
.B(n_654),
.Y(n_838)
);

BUFx5_ASAP7_75t_L g839 ( 
.A(n_691),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_730),
.B(n_655),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_707),
.B(n_655),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_676),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_676),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_710),
.A2(n_448),
.B1(n_405),
.B2(n_246),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_772),
.B(n_491),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_797),
.B(n_446),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_693),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_680),
.A2(n_431),
.B1(n_433),
.B2(n_428),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_724),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_SL g850 ( 
.A(n_793),
.B(n_268),
.C(n_263),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_710),
.B(n_711),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_684),
.B(n_255),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_693),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_711),
.B(n_255),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_702),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_719),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_703),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_683),
.B(n_314),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_687),
.B(n_280),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_703),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_682),
.B(n_660),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_736),
.A2(n_441),
.B(n_447),
.C(n_339),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_686),
.A2(n_448),
.B1(n_405),
.B2(n_246),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_692),
.A2(n_452),
.B1(n_440),
.B2(n_250),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_682),
.B(n_660),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_682),
.B(n_661),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_686),
.A2(n_448),
.B1(n_405),
.B2(n_250),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_702),
.B(n_232),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_737),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_677),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_714),
.B(n_835),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_719),
.Y(n_872)
);

AND2x2_ASAP7_75t_SL g873 ( 
.A(n_719),
.B(n_314),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_722),
.B(n_661),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_722),
.B(n_662),
.Y(n_875)
);

BUFx6f_ASAP7_75t_SL g876 ( 
.A(n_712),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_771),
.B(n_662),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_771),
.B(n_668),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_677),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_772),
.B(n_282),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_775),
.B(n_668),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_834),
.B(n_282),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_775),
.B(n_670),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_770),
.B(n_314),
.Y(n_884)
);

INVx8_ASAP7_75t_L g885 ( 
.A(n_691),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_747),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_783),
.B(n_289),
.Y(n_887)
);

AO22x1_ASAP7_75t_L g888 ( 
.A1(n_685),
.A2(n_679),
.B1(n_725),
.B2(n_691),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_L g889 ( 
.A(n_691),
.B(n_725),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_688),
.Y(n_890)
);

BUFx4_ASAP7_75t_L g891 ( 
.A(n_695),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_686),
.A2(n_259),
.B1(n_265),
.B2(n_232),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_747),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_SL g894 ( 
.A1(n_709),
.A2(n_351),
.B1(n_408),
.B2(n_389),
.Y(n_894)
);

BUFx12f_ASAP7_75t_L g895 ( 
.A(n_712),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_690),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_763),
.B(n_418),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_783),
.B(n_319),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_691),
.A2(n_259),
.B1(n_272),
.B2(n_265),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_691),
.B(n_670),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_770),
.B(n_745),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_797),
.B(n_446),
.Y(n_902)
);

NOR2x2_ASAP7_75t_L g903 ( 
.A(n_685),
.B(n_366),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_778),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_767),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_817),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_767),
.Y(n_907)
);

OR2x6_ASAP7_75t_L g908 ( 
.A(n_804),
.B(n_336),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_768),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_804),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_768),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_694),
.B(n_272),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_712),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_764),
.B(n_319),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_725),
.B(n_608),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_773),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_725),
.B(n_578),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_723),
.Y(n_918)
);

AND2x4_ASAP7_75t_SL g919 ( 
.A(n_795),
.B(n_238),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_765),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_773),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_832),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_832),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_828),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_725),
.B(n_578),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_720),
.B(n_726),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_792),
.B(n_271),
.C(n_269),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_725),
.A2(n_276),
.B1(n_283),
.B2(n_277),
.Y(n_928)
);

BUFx5_ASAP7_75t_L g929 ( 
.A(n_819),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_770),
.B(n_745),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_699),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_699),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_728),
.B(n_578),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_700),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_679),
.A2(n_276),
.B1(n_283),
.B2(n_277),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_810),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_828),
.B(n_634),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_742),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_764),
.B(n_389),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_742),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_SL g941 ( 
.A1(n_782),
.A2(n_395),
.B1(n_451),
.B2(n_429),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_828),
.B(n_288),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_729),
.B(n_578),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_833),
.B(n_288),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_731),
.B(n_297),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_833),
.B(n_297),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_833),
.B(n_303),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_686),
.A2(n_303),
.B1(n_361),
.B2(n_342),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_817),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_737),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_732),
.B(n_342),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_675),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_733),
.B(n_361),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_734),
.B(n_371),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_751),
.B(n_371),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_698),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_776),
.B(n_372),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_791),
.B(n_372),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_689),
.B(n_418),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_807),
.A2(n_399),
.B1(n_401),
.B2(n_380),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_696),
.A2(n_399),
.B1(n_401),
.B2(n_380),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_780),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_799),
.B(n_409),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_781),
.B(n_285),
.C(n_284),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_L g965 ( 
.A(n_819),
.B(n_409),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_802),
.B(n_439),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_780),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_823),
.A2(n_439),
.B1(n_480),
.B2(n_475),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_700),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_806),
.B(n_475),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_695),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_794),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_814),
.B(n_674),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_790),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_826),
.B(n_674),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_701),
.A2(n_481),
.B1(n_486),
.B2(n_480),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_794),
.A2(n_441),
.B(n_447),
.C(n_339),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_741),
.B(n_674),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_827),
.B(n_678),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_678),
.B(n_681),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_750),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_678),
.B(n_666),
.Y(n_982)
);

OAI22xp33_ASAP7_75t_L g983 ( 
.A1(n_790),
.A2(n_697),
.B1(n_755),
.B2(n_429),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_800),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_706),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_800),
.Y(n_986)
);

OAI221xp5_ASAP7_75t_L g987 ( 
.A1(n_805),
.A2(n_298),
.B1(n_382),
.B2(n_366),
.C(n_313),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_SL g988 ( 
.A(n_766),
.B(n_395),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_811),
.A2(n_275),
.B(n_313),
.C(n_278),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_701),
.A2(n_786),
.B1(n_705),
.B2(n_785),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_705),
.A2(n_819),
.B1(n_784),
.B2(n_787),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_705),
.A2(n_487),
.B1(n_481),
.B2(n_486),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_706),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_681),
.B(n_667),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_749),
.B(n_451),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_681),
.B(n_667),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_795),
.B(n_418),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_811),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_SL g999 ( 
.A1(n_708),
.A2(n_526),
.B(n_552),
.C(n_487),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_754),
.B(n_667),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_708),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_L g1002 ( 
.A(n_819),
.B(n_632),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_754),
.B(n_658),
.Y(n_1003)
);

AND2x6_ASAP7_75t_SL g1004 ( 
.A(n_715),
.B(n_278),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_L g1005 ( 
.A(n_819),
.B(n_632),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_779),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_713),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_721),
.B(n_407),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_885),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_906),
.B(n_744),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_852),
.A2(n_743),
.B1(n_746),
.B2(n_819),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_836),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_856),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_949),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_856),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_836),
.Y(n_1016)
);

AND2x6_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_754),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_885),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_849),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_894),
.B(n_750),
.C(n_295),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_852),
.B(n_705),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_938),
.B(n_795),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_858),
.A2(n_717),
.B(n_829),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_886),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_859),
.B(n_830),
.Y(n_1025)
);

AOI222xp33_ASAP7_75t_L g1026 ( 
.A1(n_941),
.A2(n_769),
.B1(n_341),
.B2(n_340),
.C1(n_335),
.C2(n_332),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_858),
.A2(n_779),
.B1(n_821),
.B2(n_818),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_904),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_859),
.B(n_813),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_871),
.B(n_813),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_872),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_926),
.B(n_744),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_886),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_845),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_893),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_893),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_907),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_907),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_911),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_950),
.B(n_782),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_911),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_851),
.B(n_713),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_885),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_921),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_921),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_871),
.A2(n_818),
.B(n_821),
.C(n_779),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_995),
.B(n_727),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_901),
.A2(n_821),
.B1(n_818),
.B2(n_718),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_922),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_922),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_SL g1051 ( 
.A(n_983),
.B(n_299),
.C(n_286),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_923),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_995),
.B(n_727),
.Y(n_1053)
);

AND2x6_ASAP7_75t_L g1054 ( 
.A(n_924),
.B(n_803),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_923),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_890),
.B(n_738),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_910),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_855),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_896),
.B(n_738),
.Y(n_1059)
);

BUFx4_ASAP7_75t_SL g1060 ( 
.A(n_910),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_870),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_931),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_924),
.B(n_813),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_931),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_842),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_988),
.B(n_716),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_855),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_838),
.B(n_739),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_940),
.B(n_739),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_855),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_840),
.B(n_758),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_926),
.B(n_824),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_855),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_895),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_926),
.B(n_824),
.Y(n_1075)
);

CKINVDCx8_ASAP7_75t_R g1076 ( 
.A(n_971),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_932),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_932),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_912),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_962),
.B(n_758),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_913),
.B(n_716),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_843),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_895),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_952),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_870),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_901),
.A2(n_718),
.B1(n_822),
.B2(n_753),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_981),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_879),
.B(n_761),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_974),
.B(n_716),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_879),
.B(n_761),
.Y(n_1090)
);

INVx6_ASAP7_75t_L g1091 ( 
.A(n_929),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_864),
.B(n_302),
.C(n_300),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_SL g1093 ( 
.A(n_977),
.B(n_309),
.C(n_304),
.Y(n_1093)
);

AO22x1_ASAP7_75t_L g1094 ( 
.A1(n_948),
.A2(n_788),
.B1(n_777),
.B2(n_317),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_984),
.B(n_998),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_905),
.B(n_774),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_869),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_934),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_839),
.B(n_717),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_934),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_969),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_969),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_985),
.Y(n_1103)
);

CKINVDCx12_ASAP7_75t_R g1104 ( 
.A(n_846),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_880),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_SL g1106 ( 
.A(n_977),
.B(n_320),
.C(n_312),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_985),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_847),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_853),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_935),
.B(n_325),
.C(n_321),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_857),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_846),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_839),
.B(n_717),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_876),
.Y(n_1114)
);

AO22x1_ASAP7_75t_L g1115 ( 
.A1(n_912),
.A2(n_868),
.B1(n_959),
.B2(n_854),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_850),
.B(n_704),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_993),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_993),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_913),
.B(n_752),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_956),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_967),
.B(n_774),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_914),
.B(n_752),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1001),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_846),
.Y(n_1124)
);

OAI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_990),
.A2(n_382),
.B1(n_438),
.B2(n_407),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1001),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_902),
.Y(n_1127)
);

BUFx4f_ASAP7_75t_L g1128 ( 
.A(n_912),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_914),
.B(n_752),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_909),
.B(n_798),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_916),
.B(n_798),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_892),
.A2(n_788),
.B1(n_777),
.B2(n_801),
.Y(n_1132)
);

NAND2x1_ASAP7_75t_L g1133 ( 
.A(n_1007),
.B(n_762),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_873),
.B(n_801),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1007),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_860),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_861),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_SL g1138 ( 
.A(n_960),
.B(n_333),
.C(n_329),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_839),
.B(n_704),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1006),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_863),
.A2(n_788),
.B1(n_777),
.B2(n_808),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_972),
.B(n_808),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_873),
.B(n_854),
.Y(n_1143)
);

CKINVDCx6p67_ASAP7_75t_R g1144 ( 
.A(n_876),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_841),
.B(n_986),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_868),
.B(n_824),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_839),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_839),
.B(n_704),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_918),
.B(n_803),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_874),
.B(n_809),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_917),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_903),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_875),
.B(n_809),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_877),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_865),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_868),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_878),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_839),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_925),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_881),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_939),
.B(n_762),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_866),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_R g1163 ( 
.A(n_920),
.B(n_809),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_980),
.Y(n_1164)
);

CKINVDCx6p67_ASAP7_75t_R g1165 ( 
.A(n_902),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_930),
.A2(n_753),
.B1(n_822),
.B2(n_718),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_936),
.B(n_824),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_939),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_973),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_930),
.A2(n_753),
.B1(n_822),
.B2(n_718),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_882),
.B(n_815),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_964),
.B(n_831),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_887),
.B(n_762),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_915),
.Y(n_1174)
);

AND2x6_ASAP7_75t_L g1175 ( 
.A(n_976),
.B(n_899),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_887),
.B(n_796),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_951),
.B(n_831),
.Y(n_1177)
);

BUFx8_ASAP7_75t_SL g1178 ( 
.A(n_891),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_951),
.B(n_831),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_883),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_862),
.B(n_927),
.C(n_347),
.Y(n_1181)
);

INVx5_ASAP7_75t_L g1182 ( 
.A(n_902),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_975),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_979),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_898),
.B(n_867),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_898),
.B(n_796),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_997),
.B(n_815),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_SL g1188 ( 
.A(n_862),
.B(n_352),
.C(n_346),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_933),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_991),
.A2(n_822),
.B1(n_753),
.B2(n_735),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_943),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_942),
.B(n_704),
.Y(n_1192)
);

CKINVDCx14_ASAP7_75t_R g1193 ( 
.A(n_908),
.Y(n_1193)
);

INVxp67_ASAP7_75t_SL g1194 ( 
.A(n_889),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_903),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_942),
.B(n_816),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_945),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_978),
.B(n_796),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_953),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_908),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1004),
.Y(n_1201)
);

BUFx8_ASAP7_75t_SL g1202 ( 
.A(n_1178),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1133),
.A2(n_1003),
.B(n_994),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1143),
.A2(n_900),
.B(n_837),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1046),
.A2(n_989),
.A3(n_957),
.B(n_963),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1021),
.A2(n_989),
.A3(n_958),
.B(n_982),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1128),
.A2(n_1194),
.B1(n_1011),
.B2(n_1025),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1147),
.A2(n_884),
.B(n_889),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1028),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1128),
.A2(n_844),
.B1(n_928),
.B2(n_968),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1023),
.A2(n_837),
.B(n_884),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1099),
.A2(n_1000),
.B(n_996),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1079),
.B(n_929),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1154),
.B(n_944),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1097),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1116),
.A2(n_946),
.B(n_944),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1133),
.A2(n_970),
.B(n_955),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1113),
.A2(n_970),
.B(n_955),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1147),
.A2(n_961),
.B(n_526),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1173),
.A2(n_937),
.B(n_888),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1128),
.A2(n_848),
.B1(n_947),
.B2(n_946),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1157),
.B(n_947),
.Y(n_1222)
);

AOI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_1029),
.A2(n_1008),
.B(n_897),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1176),
.A2(n_937),
.B(n_954),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1158),
.A2(n_966),
.B(n_820),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1190),
.A2(n_1129),
.A3(n_1161),
.B(n_1122),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1185),
.A2(n_987),
.B(n_919),
.C(n_965),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1057),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1139),
.A2(n_820),
.B(n_816),
.Y(n_1229)
);

BUFx8_ASAP7_75t_SL g1230 ( 
.A(n_1178),
.Y(n_1230)
);

AND2x6_ASAP7_75t_SL g1231 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1012),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1160),
.B(n_1008),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1079),
.A2(n_1008),
.B1(n_908),
.B2(n_919),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1147),
.A2(n_1005),
.B(n_1002),
.Y(n_1235)
);

AND2x6_ASAP7_75t_L g1236 ( 
.A(n_1009),
.B(n_929),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1158),
.A2(n_1005),
.B(n_1002),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1134),
.A2(n_965),
.B(n_735),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1072),
.B(n_831),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1010),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_SL g1241 ( 
.A1(n_1155),
.A2(n_526),
.B(n_326),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1185),
.A2(n_1175),
.B1(n_1137),
.B2(n_1162),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_1009),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1079),
.B(n_929),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1168),
.B(n_354),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1148),
.A2(n_825),
.B(n_552),
.Y(n_1246)
);

AND3x4_ASAP7_75t_L g1247 ( 
.A(n_1032),
.B(n_438),
.C(n_407),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1158),
.A2(n_748),
.B(n_740),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1067),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_L g1250 ( 
.A(n_1144),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1164),
.A2(n_825),
.B(n_561),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1164),
.A2(n_561),
.B(n_559),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1184),
.A2(n_1052),
.B(n_1035),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1180),
.B(n_929),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1072),
.B(n_559),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1042),
.A2(n_565),
.B(n_563),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1009),
.B(n_929),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1035),
.Y(n_1258)
);

AO32x2_ASAP7_75t_L g1259 ( 
.A1(n_1058),
.A2(n_999),
.A3(n_760),
.B1(n_788),
.B2(n_777),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1168),
.B(n_356),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_SL g1261 ( 
.A(n_1026),
.B(n_1051),
.C(n_1201),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1040),
.B(n_563),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1137),
.B(n_929),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1184),
.A2(n_445),
.A3(n_326),
.B(n_332),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1014),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1198),
.A2(n_748),
.B(n_740),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1145),
.A2(n_438),
.B(n_317),
.C(n_335),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1098),
.A2(n_566),
.B(n_565),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1079),
.A2(n_1156),
.B1(n_1162),
.B2(n_1155),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1169),
.A2(n_378),
.B(n_340),
.C(n_341),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1014),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1012),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1052),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1072),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1019),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1019),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1125),
.A2(n_430),
.B1(n_419),
.B2(n_454),
.C(n_417),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1150),
.A2(n_760),
.B(n_999),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1016),
.A2(n_567),
.B(n_566),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1153),
.A2(n_788),
.B(n_777),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1197),
.B(n_740),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1057),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1186),
.A2(n_748),
.B(n_740),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1086),
.A2(n_748),
.B(n_740),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1199),
.B(n_748),
.Y(n_1285)
);

AOI221x1_ASAP7_75t_L g1286 ( 
.A1(n_1116),
.A2(n_442),
.B1(n_378),
.B2(n_386),
.C(n_398),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1047),
.A2(n_571),
.B(n_567),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1016),
.A2(n_572),
.B(n_571),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1189),
.A2(n_574),
.B(n_572),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1183),
.B(n_756),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1079),
.A2(n_812),
.B1(n_789),
.B2(n_756),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1168),
.B(n_418),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1098),
.A2(n_575),
.B(n_574),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1084),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1098),
.A2(n_577),
.B(n_575),
.Y(n_1295)
);

AOI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1053),
.A2(n_577),
.B(n_398),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1166),
.A2(n_757),
.B(n_756),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1169),
.B(n_756),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1040),
.B(n_357),
.Y(n_1299)
);

O2A1O1Ixp5_ASAP7_75t_L g1300 ( 
.A1(n_1115),
.A2(n_442),
.B(n_417),
.C(n_419),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1156),
.A2(n_454),
.B(n_453),
.C(n_449),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1022),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1170),
.A2(n_757),
.B(n_756),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1036),
.Y(n_1305)
);

CKINVDCx12_ASAP7_75t_R g1306 ( 
.A(n_1022),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1068),
.A2(n_788),
.B(n_777),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1037),
.A2(n_386),
.A3(n_410),
.B(n_430),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1034),
.B(n_1105),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1187),
.B(n_444),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1048),
.A2(n_432),
.B(n_410),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1038),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1156),
.A2(n_812),
.B1(n_789),
.B2(n_759),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1171),
.B(n_757),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1071),
.A2(n_652),
.B(n_445),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1032),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1027),
.A2(n_789),
.B1(n_759),
.B2(n_757),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1115),
.B(n_757),
.Y(n_1318)
);

AO32x2_ASAP7_75t_L g1319 ( 
.A1(n_1058),
.A2(n_432),
.A3(n_449),
.B1(n_453),
.B2(n_444),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1065),
.B(n_759),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1039),
.A2(n_789),
.B(n_759),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1067),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1043),
.A2(n_789),
.B(n_759),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1082),
.B(n_812),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1043),
.A2(n_812),
.B(n_633),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1092),
.A2(n_238),
.B1(n_279),
.B2(n_323),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1108),
.B(n_812),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1175),
.A2(n_1110),
.B1(n_1138),
.B2(n_1041),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1016),
.A2(n_652),
.B(n_119),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_1061),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1152),
.B(n_444),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1181),
.A2(n_370),
.B(n_368),
.C(n_367),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1152),
.B(n_359),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1109),
.B(n_360),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1041),
.A2(n_10),
.A3(n_12),
.B(n_13),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1049),
.A2(n_15),
.A3(n_16),
.B(n_18),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1174),
.B(n_238),
.Y(n_1337)
);

NAND2x1_ASAP7_75t_L g1338 ( 
.A(n_1091),
.B(n_632),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1091),
.A2(n_403),
.B1(n_363),
.B2(n_376),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1091),
.A2(n_412),
.B1(n_365),
.B2(n_379),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1049),
.Y(n_1341)
);

BUFx12f_ASAP7_75t_L g1342 ( 
.A(n_1114),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1107),
.A2(n_652),
.B(n_120),
.Y(n_1343)
);

OA22x2_ASAP7_75t_L g1344 ( 
.A1(n_1195),
.A2(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1111),
.B(n_381),
.Y(n_1345)
);

AO22x1_ASAP7_75t_L g1346 ( 
.A1(n_1201),
.A2(n_1087),
.B1(n_1200),
.B2(n_1182),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1043),
.A2(n_633),
.B(n_632),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1196),
.A2(n_652),
.B(n_393),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1050),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1142),
.B(n_384),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1107),
.A2(n_199),
.B(n_124),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1043),
.A2(n_633),
.B(n_632),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1091),
.A2(n_425),
.B1(n_387),
.B2(n_388),
.Y(n_1353)
);

OA21x2_ASAP7_75t_L g1354 ( 
.A1(n_1189),
.A2(n_426),
.B(n_394),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1142),
.B(n_406),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1050),
.A2(n_16),
.A3(n_19),
.B(n_20),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1136),
.B(n_413),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1196),
.A2(n_435),
.B(n_416),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1043),
.A2(n_633),
.B(n_632),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1107),
.A2(n_202),
.B(n_133),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1195),
.B(n_1095),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1055),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1060),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1024),
.A2(n_207),
.B(n_134),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1067),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1249),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1232),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1361),
.B(n_1209),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1215),
.Y(n_1369)
);

NOR4xp25_ASAP7_75t_L g1370 ( 
.A(n_1261),
.B(n_1063),
.C(n_1140),
.D(n_1031),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1247),
.A2(n_1175),
.B1(n_1136),
.B2(n_1066),
.Y(n_1371)
);

BUFx2_ASAP7_75t_SL g1372 ( 
.A(n_1265),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1343),
.A2(n_1130),
.B(n_1096),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1302),
.B(n_1087),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1242),
.B(n_1069),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1232),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1256),
.A2(n_1131),
.B(n_1045),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1304),
.B(n_1069),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1321),
.A2(n_1224),
.B(n_1220),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1242),
.B(n_1080),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1223),
.A2(n_1020),
.B1(n_1112),
.B2(n_1127),
.C(n_1188),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1216),
.A2(n_1055),
.B(n_1056),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1258),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1214),
.B(n_1080),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1208),
.B(n_1067),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1282),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1225),
.A2(n_1033),
.B(n_1024),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1207),
.A2(n_1191),
.B(n_1090),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1274),
.B(n_1075),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1302),
.B(n_1120),
.Y(n_1390)
);

INVx6_ASAP7_75t_L g1391 ( 
.A(n_1228),
.Y(n_1391)
);

AO21x1_ASAP7_75t_L g1392 ( 
.A1(n_1221),
.A2(n_1337),
.B(n_1269),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1227),
.A2(n_1088),
.B(n_1059),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1272),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1273),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1256),
.A2(n_1064),
.B(n_1062),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1227),
.A2(n_1192),
.B(n_1121),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1245),
.A2(n_1193),
.B1(n_1182),
.B2(n_1200),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1211),
.A2(n_1064),
.B(n_1062),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1225),
.A2(n_1329),
.B(n_1288),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1247),
.A2(n_1175),
.B1(n_1121),
.B2(n_1033),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1271),
.B(n_1076),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1274),
.B(n_1075),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1275),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1239),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1276),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1228),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1278),
.A2(n_1078),
.B(n_1077),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1265),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1222),
.B(n_1200),
.Y(n_1410)
);

BUFx4_ASAP7_75t_SL g1411 ( 
.A(n_1271),
.Y(n_1411)
);

BUFx8_ASAP7_75t_L g1412 ( 
.A(n_1342),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1243),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1233),
.A2(n_1061),
.B1(n_1085),
.B2(n_1200),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1239),
.B(n_1075),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1329),
.A2(n_1033),
.B(n_1024),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1286),
.A2(n_1101),
.A3(n_1077),
.B(n_1078),
.Y(n_1417)
);

AO21x1_ASAP7_75t_L g1418 ( 
.A1(n_1337),
.A2(n_1089),
.B(n_1172),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1204),
.A2(n_1015),
.B(n_1172),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1245),
.A2(n_1193),
.B1(n_1182),
.B2(n_1200),
.Y(n_1420)
);

AND2x2_ASAP7_75t_SL g1421 ( 
.A(n_1328),
.B(n_1009),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1238),
.A2(n_1172),
.B(n_1175),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1279),
.A2(n_1044),
.B(n_1117),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1279),
.A2(n_1044),
.B(n_1117),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1306),
.Y(n_1425)
);

AOI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1260),
.A2(n_1013),
.B(n_1182),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1260),
.A2(n_1120),
.B1(n_1104),
.B2(n_1124),
.Y(n_1427)
);

AOI21xp33_ASAP7_75t_L g1428 ( 
.A1(n_1299),
.A2(n_1013),
.B(n_1182),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1262),
.B(n_1165),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1312),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1294),
.B(n_1061),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1252),
.A2(n_1101),
.B(n_1100),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1316),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1250),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1341),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1349),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1362),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1202),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1272),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1305),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1210),
.A2(n_1093),
.B(n_1106),
.C(n_1044),
.Y(n_1441)
);

AOI222xp33_ASAP7_75t_L g1442 ( 
.A1(n_1331),
.A2(n_444),
.B1(n_1124),
.B2(n_434),
.C1(n_450),
.C2(n_422),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1328),
.A2(n_1085),
.B1(n_1174),
.B2(n_1013),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1305),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1326),
.A2(n_1175),
.B1(n_1017),
.B2(n_279),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1288),
.A2(n_1118),
.B(n_1135),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1212),
.A2(n_1251),
.B(n_1203),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1241),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1253),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1294),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1308),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1308),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1350),
.B(n_1085),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1212),
.A2(n_1118),
.B(n_1135),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1355),
.B(n_1085),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_SL g1456 ( 
.A1(n_1332),
.A2(n_1102),
.B(n_1103),
.C(n_1126),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1318),
.A2(n_1123),
.B(n_1100),
.Y(n_1457)
);

INVx4_ASAP7_75t_SL g1458 ( 
.A(n_1249),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1253),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1333),
.B(n_1165),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1240),
.A2(n_1114),
.B1(n_1144),
.B2(n_1074),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1308),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1300),
.A2(n_1132),
.B(n_1141),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1308),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1249),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1250),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1255),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1253),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1330),
.A2(n_1085),
.B1(n_1174),
.B2(n_1070),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1254),
.A2(n_1017),
.B(n_1102),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1246),
.A2(n_1117),
.B(n_1118),
.Y(n_1471)
);

NOR2xp67_ASAP7_75t_L g1472 ( 
.A(n_1240),
.B(n_1058),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1310),
.B(n_1151),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1284),
.A2(n_1135),
.B(n_1103),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1309),
.B(n_1076),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1234),
.A2(n_1083),
.B1(n_1074),
.B2(n_1174),
.Y(n_1476)
);

AOI21xp33_ASAP7_75t_L g1477 ( 
.A1(n_1358),
.A2(n_1159),
.B(n_1151),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1330),
.A2(n_1263),
.B1(n_1174),
.B2(n_1070),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1315),
.A2(n_1123),
.B(n_1126),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1270),
.A2(n_437),
.B1(n_427),
.B2(n_424),
.C(n_1083),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1255),
.B(n_1146),
.Y(n_1481)
);

BUFx4f_ASAP7_75t_L g1482 ( 
.A(n_1239),
.Y(n_1482)
);

INVx5_ASAP7_75t_L g1483 ( 
.A(n_1236),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1297),
.A2(n_1119),
.B(n_1081),
.Y(n_1484)
);

NAND2x1_ASAP7_75t_L g1485 ( 
.A(n_1236),
.B(n_1054),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1255),
.B(n_1146),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1342),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1243),
.B(n_1146),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1292),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1357),
.B(n_1151),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1314),
.A2(n_1070),
.B1(n_1081),
.B2(n_1119),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1303),
.A2(n_1119),
.B(n_1081),
.Y(n_1492)
);

AOI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1283),
.A2(n_1094),
.B(n_1177),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1364),
.A2(n_1179),
.B(n_1177),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1249),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1363),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_SL g1497 ( 
.A1(n_1219),
.A2(n_1017),
.B(n_1054),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1344),
.A2(n_1159),
.B1(n_1151),
.B2(n_1070),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1364),
.A2(n_1179),
.B(n_1177),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1268),
.A2(n_1151),
.B(n_1159),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_SL g1501 ( 
.A1(n_1332),
.A2(n_1301),
.B(n_1270),
.C(n_1267),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1293),
.Y(n_1502)
);

INVx3_ASAP7_75t_SL g1503 ( 
.A(n_1344),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1281),
.A2(n_1070),
.B1(n_1159),
.B2(n_1067),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1226),
.B(n_1159),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1243),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1264),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1295),
.A2(n_1179),
.B(n_1167),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1218),
.A2(n_1017),
.B(n_1054),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1351),
.A2(n_1054),
.B(n_1017),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1360),
.A2(n_1054),
.B(n_1017),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1285),
.A2(n_1073),
.B1(n_1018),
.B2(n_1009),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1202),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1296),
.A2(n_1167),
.B(n_1094),
.Y(n_1514)
);

AOI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1266),
.A2(n_1167),
.B(n_1054),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1264),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1229),
.A2(n_1217),
.B(n_1235),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1226),
.B(n_1334),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1230),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1301),
.A2(n_1104),
.B(n_1149),
.C(n_1163),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1267),
.A2(n_1073),
.B1(n_1018),
.B2(n_362),
.C(n_323),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1243),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1339),
.B(n_1073),
.C(n_1018),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1257),
.A2(n_1018),
.B(n_1073),
.Y(n_1524)
);

INVx4_ASAP7_75t_SL g1525 ( 
.A(n_1322),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1237),
.A2(n_1018),
.B(n_672),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1322),
.B(n_658),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1363),
.A2(n_1345),
.B1(n_1231),
.B2(n_1353),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1340),
.B(n_20),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1348),
.A2(n_1290),
.B(n_1354),
.C(n_1327),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1322),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1322),
.B(n_118),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1307),
.A2(n_238),
.B(n_279),
.Y(n_1533)
);

AO21x1_ASAP7_75t_L g1534 ( 
.A1(n_1317),
.A2(n_1298),
.B(n_1257),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1320),
.A2(n_672),
.B1(n_658),
.B2(n_633),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1365),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1365),
.Y(n_1537)
);

AO31x2_ASAP7_75t_L g1538 ( 
.A1(n_1313),
.A2(n_362),
.A3(n_323),
.B(n_279),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1264),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1264),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_L g1541 ( 
.A(n_1277),
.B(n_362),
.C(n_323),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1248),
.A2(n_672),
.B(n_658),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1354),
.A2(n_362),
.B(n_22),
.C(n_25),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1346),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1311),
.A2(n_672),
.B1(n_658),
.B2(n_633),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1280),
.A2(n_186),
.B(n_153),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1483),
.B(n_1365),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1506),
.Y(n_1548)
);

NAND2x1p5_ASAP7_75t_L g1549 ( 
.A(n_1483),
.B(n_1365),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1367),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1533),
.A2(n_1388),
.B(n_1518),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1505),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1408),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1408),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1482),
.Y(n_1555)
);

INVx6_ASAP7_75t_L g1556 ( 
.A(n_1391),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1529),
.A2(n_1311),
.B1(n_1354),
.B2(n_1287),
.Y(n_1557)
);

BUFx8_ASAP7_75t_L g1558 ( 
.A(n_1487),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1369),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1411),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1418),
.A2(n_1287),
.B(n_1213),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1422),
.A2(n_1226),
.B(n_1324),
.C(n_1213),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1368),
.B(n_1473),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1385),
.A2(n_1244),
.B(n_1323),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1529),
.A2(n_1289),
.B1(n_1244),
.B2(n_1226),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1445),
.A2(n_1289),
.B1(n_1319),
.B2(n_1236),
.Y(n_1566)
);

OR2x6_ASAP7_75t_L g1567 ( 
.A(n_1385),
.B(n_1338),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1445),
.A2(n_1289),
.B1(n_1319),
.B2(n_1236),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1482),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1371),
.A2(n_1291),
.B1(n_1325),
.B2(n_1352),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1383),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1378),
.B(n_1206),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1475),
.B(n_1230),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1385),
.A2(n_1347),
.B(n_1359),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1442),
.A2(n_1528),
.B1(n_1371),
.B2(n_1392),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1384),
.B(n_1206),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1541),
.A2(n_1319),
.B1(n_1236),
.B2(n_1206),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1506),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1503),
.A2(n_1421),
.B1(n_1375),
.B2(n_1380),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1490),
.B(n_1205),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1395),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1490),
.B(n_1206),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1506),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1379),
.A2(n_1259),
.B(n_1205),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1503),
.A2(n_1319),
.B1(n_1336),
.B2(n_1335),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1413),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1386),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1401),
.A2(n_1205),
.B1(n_1259),
.B2(n_672),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1421),
.A2(n_1356),
.B1(n_1336),
.B2(n_1335),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1404),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1406),
.Y(n_1591)
);

NOR3xp33_ASAP7_75t_SL g1592 ( 
.A(n_1476),
.B(n_1356),
.C(n_1336),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1409),
.A2(n_1356),
.B1(n_1336),
.B2(n_1335),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1401),
.A2(n_1205),
.B1(n_1259),
.B2(n_672),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1433),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_R g1596 ( 
.A(n_1402),
.B(n_141),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1481),
.B(n_1390),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1374),
.A2(n_1259),
.B1(n_672),
.B2(n_658),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1480),
.A2(n_658),
.B1(n_1356),
.B2(n_1335),
.C(n_27),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1438),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1430),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1453),
.A2(n_21),
.B(n_25),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1391),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1376),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1433),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1475),
.A2(n_633),
.B1(n_26),
.B2(n_28),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1455),
.B(n_21),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1375),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1391),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1380),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1513),
.Y(n_1611)
);

AND2x6_ASAP7_75t_L g1612 ( 
.A(n_1532),
.B(n_229),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1435),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1546),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1489),
.B(n_32),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1498),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.C(n_41),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1482),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1394),
.Y(n_1618)
);

AO31x2_ASAP7_75t_L g1619 ( 
.A1(n_1507),
.A2(n_41),
.A3(n_42),
.B(n_45),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1441),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1412),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_SL g1622 ( 
.A1(n_1441),
.A2(n_47),
.B(n_51),
.C(n_52),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1374),
.B(n_54),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1390),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1440),
.Y(n_1625)
);

OAI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1381),
.A2(n_1370),
.B1(n_1427),
.B2(n_1429),
.C(n_1460),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1436),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1407),
.B(n_62),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1450),
.B(n_68),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1513),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1398),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1486),
.B(n_228),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1437),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1483),
.B(n_1413),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1501),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.C(n_78),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1372),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1410),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_1637)
);

INVx8_ASAP7_75t_L g1638 ( 
.A(n_1488),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1496),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1483),
.B(n_227),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1496),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1439),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1483),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1444),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1412),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1431),
.B(n_84),
.Y(n_1646)
);

NAND2x1p5_ASAP7_75t_L g1647 ( 
.A(n_1413),
.B(n_225),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1431),
.B(n_86),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1544),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1434),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1440),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1486),
.B(n_219),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1486),
.B(n_213),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1425),
.B(n_97),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1428),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1385),
.A2(n_191),
.B(n_182),
.Y(n_1656)
);

O2A1O1Ixp5_ASAP7_75t_SL g1657 ( 
.A1(n_1516),
.A2(n_98),
.B(n_100),
.C(n_101),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1420),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1434),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1539),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1472),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1426),
.B(n_1477),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1415),
.B(n_1405),
.Y(n_1663)
);

OAI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1543),
.A2(n_1521),
.B1(n_1393),
.B2(n_1501),
.C(n_1520),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1466),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1467),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_1666)
);

OAI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1463),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1397),
.A2(n_110),
.B1(n_159),
.B2(n_160),
.C(n_164),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1524),
.A2(n_166),
.B(n_167),
.Y(n_1669)
);

CKINVDCx6p67_ASAP7_75t_R g1670 ( 
.A(n_1487),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1409),
.A2(n_173),
.B1(n_180),
.B2(n_1412),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1488),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1415),
.B(n_1389),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1523),
.A2(n_1443),
.B1(n_1532),
.B2(n_1466),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1415),
.B(n_1389),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1389),
.B(n_1403),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1540),
.A2(n_1382),
.B1(n_1419),
.B2(n_1448),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1534),
.A2(n_1451),
.B1(n_1462),
.B2(n_1452),
.Y(n_1678)
);

CKINVDCx8_ASAP7_75t_R g1679 ( 
.A(n_1519),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1403),
.B(n_1532),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1403),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1464),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1531),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1497),
.B(n_1485),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1488),
.B(n_1537),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1537),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1447),
.A2(n_1416),
.B(n_1400),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1366),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1536),
.B(n_1538),
.Y(n_1689)
);

OAI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1470),
.A2(n_1530),
.B(n_1414),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1457),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1366),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1461),
.B(n_1538),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1519),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1457),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1538),
.B(n_1495),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1366),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1538),
.B(n_1465),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1458),
.B(n_1525),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1458),
.B(n_1525),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1457),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1417),
.Y(n_1702)
);

OAI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1545),
.A2(n_1522),
.B1(n_1478),
.B2(n_1469),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1458),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1509),
.B(n_1491),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1417),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1447),
.A2(n_1416),
.B(n_1400),
.Y(n_1707)
);

INVx6_ASAP7_75t_L g1708 ( 
.A(n_1525),
.Y(n_1708)
);

AND2x4_ASAP7_75t_SL g1709 ( 
.A(n_1366),
.B(n_1495),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1465),
.B(n_1468),
.Y(n_1710)
);

INVx8_ASAP7_75t_L g1711 ( 
.A(n_1527),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1417),
.B(n_1527),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1408),
.A2(n_1399),
.B1(n_1479),
.B2(n_1514),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1399),
.A2(n_1479),
.B1(n_1514),
.B2(n_1468),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1417),
.B(n_1459),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1504),
.B(n_1456),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1399),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1510),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1479),
.A2(n_1514),
.B1(n_1449),
.B2(n_1377),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1474),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1377),
.A2(n_1494),
.B1(n_1499),
.B2(n_1502),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1512),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1456),
.B(n_1474),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1724)
);

AND2x4_ASAP7_75t_SL g1725 ( 
.A(n_1502),
.B(n_1493),
.Y(n_1725)
);

O2A1O1Ixp5_ASAP7_75t_L g1726 ( 
.A1(n_1515),
.A2(n_1535),
.B(n_1494),
.C(n_1499),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1432),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_R g1728 ( 
.A(n_1511),
.B(n_1499),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1432),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1508),
.B(n_1494),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1508),
.B(n_1377),
.Y(n_1731)
);

NAND2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1508),
.B(n_1492),
.Y(n_1732)
);

AO31x2_ASAP7_75t_L g1733 ( 
.A1(n_1517),
.A2(n_1396),
.A3(n_1526),
.B(n_1454),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1432),
.Y(n_1734)
);

OAI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1396),
.A2(n_1492),
.B1(n_1484),
.B2(n_1387),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1387),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1641),
.B(n_1639),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1575),
.A2(n_1396),
.B1(n_1484),
.B2(n_1500),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1575),
.A2(n_1373),
.B1(n_1454),
.B2(n_1424),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1667),
.A2(n_1373),
.B1(n_1517),
.B2(n_1526),
.C(n_1500),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1624),
.A2(n_1423),
.B1(n_1424),
.B2(n_1446),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1614),
.A2(n_1423),
.B1(n_1471),
.B2(n_1446),
.Y(n_1742)
);

INVxp67_ASAP7_75t_R g1743 ( 
.A(n_1597),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1624),
.A2(n_1471),
.B1(n_1542),
.B2(n_1667),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1726),
.A2(n_1542),
.B(n_1690),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1649),
.A2(n_1614),
.B1(n_1620),
.B2(n_1637),
.C(n_1643),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1608),
.B(n_1563),
.Y(n_1747)
);

OAI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1606),
.A2(n_1649),
.B1(n_1635),
.B2(n_1643),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1664),
.A2(n_1626),
.B(n_1693),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1569),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1571),
.Y(n_1751)
);

BUFx10_ASAP7_75t_L g1752 ( 
.A(n_1560),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1608),
.B(n_1582),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1637),
.A2(n_1610),
.B1(n_1622),
.B2(n_1666),
.C(n_1658),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1581),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1636),
.A2(n_1610),
.B1(n_1666),
.B2(n_1658),
.Y(n_1756)
);

AND2x4_ASAP7_75t_SL g1757 ( 
.A(n_1569),
.B(n_1548),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1590),
.Y(n_1758)
);

OAI211xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1623),
.A2(n_1636),
.B(n_1615),
.C(n_1646),
.Y(n_1759)
);

AOI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1622),
.A2(n_1551),
.B1(n_1602),
.B2(n_1631),
.C(n_1655),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1612),
.A2(n_1573),
.B1(n_1668),
.B2(n_1653),
.Y(n_1761)
);

NOR2xp67_ASAP7_75t_L g1762 ( 
.A(n_1603),
.B(n_1609),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1655),
.A2(n_1671),
.B1(n_1629),
.B2(n_1612),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1596),
.A2(n_1612),
.B1(n_1661),
.B2(n_1648),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1596),
.A2(n_1612),
.B1(n_1640),
.B2(n_1656),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1671),
.A2(n_1629),
.B1(n_1612),
.B2(n_1579),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_SL g1767 ( 
.A(n_1694),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1591),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1567),
.B(n_1684),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1616),
.A2(n_1599),
.B1(n_1585),
.B2(n_1579),
.C(n_1593),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1674),
.A2(n_1559),
.B1(n_1607),
.B2(n_1654),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1674),
.A2(n_1566),
.B1(n_1568),
.B2(n_1645),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1587),
.A2(n_1659),
.B1(n_1605),
.B2(n_1595),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1681),
.B(n_1552),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1659),
.A2(n_1650),
.B1(n_1665),
.B2(n_1617),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1552),
.B(n_1683),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1566),
.A2(n_1568),
.B1(n_1565),
.B2(n_1628),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1557),
.A2(n_1669),
.B1(n_1722),
.B2(n_1662),
.C(n_1565),
.Y(n_1778)
);

OAI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1722),
.A2(n_1569),
.B1(n_1598),
.B2(n_1640),
.Y(n_1779)
);

OAI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1557),
.A2(n_1662),
.B1(n_1647),
.B2(n_1577),
.C(n_1677),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1675),
.A2(n_1632),
.B1(n_1652),
.B2(n_1585),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1647),
.A2(n_1577),
.B1(n_1677),
.B2(n_1562),
.C(n_1676),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1580),
.A2(n_1705),
.B1(n_1562),
.B2(n_1678),
.C(n_1572),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1611),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1675),
.A2(n_1580),
.B1(n_1613),
.B2(n_1601),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1682),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1555),
.B(n_1617),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1670),
.A2(n_1680),
.B1(n_1621),
.B2(n_1555),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1556),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1663),
.B(n_1627),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1633),
.A2(n_1558),
.B1(n_1673),
.B2(n_1570),
.Y(n_1791)
);

INVx5_ASAP7_75t_SL g1792 ( 
.A(n_1699),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1696),
.A2(n_1698),
.B1(n_1705),
.B2(n_1576),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1558),
.A2(n_1589),
.B1(n_1588),
.B2(n_1594),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1589),
.A2(n_1716),
.B1(n_1642),
.B2(n_1644),
.Y(n_1795)
);

AOI33xp33_ASAP7_75t_L g1796 ( 
.A1(n_1678),
.A2(n_1689),
.A3(n_1660),
.B1(n_1686),
.B2(n_1721),
.B3(n_1719),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1630),
.A2(n_1638),
.B(n_1600),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1710),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1716),
.A2(n_1703),
.B1(n_1556),
.B2(n_1672),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1564),
.A2(n_1574),
.B(n_1592),
.C(n_1725),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1556),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1703),
.A2(n_1672),
.B1(n_1638),
.B2(n_1567),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1604),
.B(n_1618),
.Y(n_1803)
);

OAI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1592),
.A2(n_1679),
.B(n_1721),
.C(n_1730),
.Y(n_1804)
);

BUFx4f_ASAP7_75t_L g1805 ( 
.A(n_1708),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1638),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1634),
.A2(n_1548),
.B1(n_1583),
.B2(n_1578),
.C(n_1726),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1625),
.A2(n_1651),
.B1(n_1685),
.B2(n_1578),
.Y(n_1808)
);

AOI222xp33_ASAP7_75t_L g1809 ( 
.A1(n_1583),
.A2(n_1704),
.B1(n_1699),
.B2(n_1700),
.C1(n_1712),
.C2(n_1730),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1553),
.Y(n_1810)
);

OAI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1704),
.A2(n_1708),
.B1(n_1634),
.B2(n_1586),
.Y(n_1811)
);

AO21x2_ASAP7_75t_L g1812 ( 
.A1(n_1735),
.A2(n_1723),
.B(n_1728),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1619),
.B(n_1715),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1731),
.A2(n_1657),
.B(n_1719),
.C(n_1713),
.Y(n_1814)
);

A2O1A1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1700),
.A2(n_1731),
.B(n_1711),
.C(n_1709),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1688),
.B(n_1697),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1735),
.A2(n_1547),
.B(n_1549),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1708),
.A2(n_1561),
.B1(n_1701),
.B2(n_1695),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1561),
.A2(n_1691),
.B1(n_1684),
.B2(n_1586),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1619),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1684),
.A2(n_1720),
.B1(n_1706),
.B2(n_1702),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1547),
.A2(n_1549),
.B1(n_1711),
.B2(n_1697),
.Y(n_1822)
);

CKINVDCx11_ASAP7_75t_R g1823 ( 
.A(n_1688),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1688),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1713),
.A2(n_1553),
.B1(n_1554),
.B2(n_1714),
.C(n_1728),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1711),
.A2(n_1697),
.B1(n_1692),
.B2(n_1688),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1692),
.A2(n_1697),
.B1(n_1584),
.B2(n_1554),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1692),
.Y(n_1828)
);

OAI211xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1714),
.A2(n_1736),
.B(n_1717),
.C(n_1729),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1692),
.A2(n_1718),
.B1(n_1734),
.B2(n_1727),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1718),
.A2(n_1736),
.B1(n_1732),
.B2(n_1619),
.C(n_1724),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1619),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1718),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_SL g1834 ( 
.A1(n_1724),
.A2(n_1718),
.B(n_1732),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1724),
.A2(n_1687),
.B1(n_1707),
.B2(n_1733),
.Y(n_1835)
);

AOI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1733),
.A2(n_1029),
.B(n_852),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1733),
.A2(n_852),
.B1(n_859),
.B2(n_1667),
.C(n_871),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1733),
.A2(n_1029),
.B1(n_1575),
.B2(n_1636),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1641),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1676),
.B(n_769),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1556),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1559),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_852),
.B2(n_1030),
.Y(n_1843)
);

OR2x6_ASAP7_75t_L g1844 ( 
.A(n_1567),
.B(n_1684),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1665),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_1529),
.B2(n_1029),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1606),
.A2(n_1649),
.B1(n_656),
.B2(n_583),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1552),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1575),
.A2(n_1029),
.B(n_1030),
.C(n_871),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1606),
.A2(n_1649),
.B1(n_656),
.B2(n_583),
.Y(n_1851)
);

BUFx12f_ASAP7_75t_L g1852 ( 
.A(n_1560),
.Y(n_1852)
);

BUFx5_ASAP7_75t_L g1853 ( 
.A(n_1720),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1667),
.A2(n_852),
.B1(n_859),
.B2(n_871),
.C(n_680),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_1636),
.B2(n_852),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1668),
.A2(n_1029),
.B1(n_1030),
.B2(n_852),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1667),
.A2(n_852),
.B1(n_859),
.B2(n_871),
.C(n_680),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_852),
.B2(n_1030),
.Y(n_1859)
);

OAI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1624),
.A2(n_852),
.B(n_1026),
.C(n_859),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_852),
.B2(n_1030),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1667),
.A2(n_852),
.B1(n_859),
.B2(n_871),
.C(n_680),
.Y(n_1863)
);

AOI33xp33_ASAP7_75t_L g1864 ( 
.A1(n_1636),
.A2(n_1624),
.A3(n_1649),
.B1(n_983),
.B2(n_959),
.B3(n_1667),
.Y(n_1864)
);

AOI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1667),
.A2(n_852),
.B1(n_859),
.B2(n_871),
.C(n_680),
.Y(n_1865)
);

OAI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1575),
.A2(n_1624),
.B1(n_1614),
.B2(n_1636),
.C1(n_1606),
.C2(n_1610),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1668),
.A2(n_1029),
.B1(n_1030),
.B2(n_852),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_852),
.B2(n_1030),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1606),
.A2(n_1649),
.B1(n_656),
.B2(n_583),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1624),
.A2(n_852),
.B(n_1026),
.C(n_859),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_SL g1871 ( 
.A1(n_1668),
.A2(n_1029),
.B1(n_1030),
.B2(n_852),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1641),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1676),
.B(n_769),
.Y(n_1873)
);

INVx6_ASAP7_75t_L g1874 ( 
.A(n_1704),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1563),
.B(n_1559),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1559),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1550),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1667),
.A2(n_852),
.B1(n_859),
.B2(n_871),
.C(n_680),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1641),
.B(n_1639),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1606),
.A2(n_1649),
.B1(n_656),
.B2(n_583),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_852),
.B2(n_1030),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1667),
.A2(n_852),
.B1(n_859),
.B2(n_871),
.C(n_680),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1575),
.A2(n_1029),
.B1(n_852),
.B2(n_1030),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1885)
);

CKINVDCx6p67_ASAP7_75t_R g1886 ( 
.A(n_1645),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1556),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1552),
.Y(n_1889)
);

OA21x2_ASAP7_75t_L g1890 ( 
.A1(n_1726),
.A2(n_1690),
.B(n_1723),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1556),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1563),
.B(n_1559),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1641),
.B(n_1639),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1575),
.A2(n_852),
.B1(n_859),
.B2(n_1624),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1753),
.B(n_1786),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1786),
.B(n_1813),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1848),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1853),
.Y(n_1899)
);

NOR2x1_ASAP7_75t_L g1900 ( 
.A(n_1807),
.B(n_1811),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1751),
.B(n_1755),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1758),
.B(n_1768),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1820),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1769),
.B(n_1844),
.Y(n_1904)
);

OR2x6_ASAP7_75t_SL g1905 ( 
.A(n_1843),
.B(n_1859),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1832),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1810),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1854),
.B(n_1857),
.Y(n_1908)
);

OAI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1863),
.A2(n_1879),
.B1(n_1883),
.B2(n_1865),
.C(n_1846),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1810),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1889),
.B(n_1747),
.Y(n_1911)
);

AND2x4_ASAP7_75t_SL g1912 ( 
.A(n_1769),
.B(n_1844),
.Y(n_1912)
);

OR2x6_ASAP7_75t_L g1913 ( 
.A(n_1769),
.B(n_1844),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1889),
.B(n_1776),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1876),
.Y(n_1915)
);

OR2x6_ASAP7_75t_L g1916 ( 
.A(n_1817),
.B(n_1834),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1890),
.B(n_1812),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1890),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1833),
.B(n_1835),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1798),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1790),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1745),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1833),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1860),
.A2(n_1870),
.B1(n_1875),
.B2(n_1891),
.C(n_1888),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1812),
.B(n_1893),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1811),
.B(n_1804),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1878),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1793),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1800),
.B(n_1815),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1774),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1814),
.B(n_1821),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1803),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1738),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1842),
.B(n_1877),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1749),
.B(n_1771),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1773),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1795),
.B(n_1783),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1795),
.B(n_1825),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1778),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1821),
.B(n_1819),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1831),
.Y(n_1941)
);

AO21x2_ASAP7_75t_L g1942 ( 
.A1(n_1836),
.A2(n_1827),
.B(n_1780),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1737),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1777),
.B(n_1794),
.Y(n_1944)
);

NAND2x1p5_ASAP7_75t_L g1945 ( 
.A(n_1805),
.B(n_1737),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1777),
.B(n_1794),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1796),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1819),
.B(n_1830),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1771),
.B(n_1840),
.Y(n_1949)
);

INVx5_ASAP7_75t_L g1950 ( 
.A(n_1828),
.Y(n_1950)
);

NAND2x1p5_ASAP7_75t_L g1951 ( 
.A(n_1805),
.B(n_1880),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1880),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1894),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1782),
.Y(n_1954)
);

INVx4_ASAP7_75t_R g1955 ( 
.A(n_1845),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1849),
.B(n_1868),
.C(n_1862),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1818),
.B(n_1785),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1818),
.B(n_1785),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1816),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1827),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1830),
.B(n_1743),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1772),
.B(n_1781),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1829),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1740),
.Y(n_1964)
);

BUFx2_ASAP7_75t_SL g1965 ( 
.A(n_1767),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1826),
.Y(n_1966)
);

NAND2x1_ASAP7_75t_L g1967 ( 
.A(n_1802),
.B(n_1799),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1826),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1772),
.B(n_1781),
.Y(n_1969)
);

AND2x4_ASAP7_75t_SL g1970 ( 
.A(n_1802),
.B(n_1799),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1808),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1739),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1787),
.B(n_1750),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1784),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1739),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1741),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1741),
.Y(n_1977)
);

INVxp67_ASAP7_75t_L g1978 ( 
.A(n_1839),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1872),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1791),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1921),
.B(n_1770),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1908),
.A2(n_1884),
.B1(n_1882),
.B2(n_1881),
.C(n_1869),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1959),
.B(n_1897),
.Y(n_1983)
);

AOI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1909),
.A2(n_1869),
.B1(n_1881),
.B2(n_1851),
.C(n_1847),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1956),
.A2(n_1855),
.B1(n_1871),
.B2(n_1856),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1956),
.A2(n_1847),
.B1(n_1851),
.B2(n_1759),
.C(n_1748),
.Y(n_1986)
);

OAI22xp33_ASAP7_75t_SL g1987 ( 
.A1(n_1905),
.A2(n_1761),
.B1(n_1788),
.B2(n_1775),
.Y(n_1987)
);

AO21x2_ASAP7_75t_L g1988 ( 
.A1(n_1964),
.A2(n_1748),
.B(n_1779),
.Y(n_1988)
);

OAI31xp33_ASAP7_75t_L g1989 ( 
.A1(n_1924),
.A2(n_1866),
.A3(n_1895),
.B(n_1885),
.Y(n_1989)
);

OR2x6_ASAP7_75t_L g1990 ( 
.A(n_1913),
.B(n_1838),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1959),
.B(n_1791),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_R g1992 ( 
.A(n_1974),
.B(n_1852),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1925),
.B(n_1742),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1907),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1905),
.A2(n_1895),
.B1(n_1861),
.B2(n_1891),
.Y(n_1995)
);

OAI33xp33_ASAP7_75t_L g1996 ( 
.A1(n_1935),
.A2(n_1779),
.A3(n_1824),
.B1(n_1822),
.B2(n_1864),
.B3(n_1837),
.Y(n_1996)
);

NAND3xp33_ASAP7_75t_L g1997 ( 
.A(n_1964),
.B(n_1867),
.C(n_1885),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1937),
.A2(n_1875),
.B1(n_1861),
.B2(n_1888),
.C(n_1850),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1937),
.A2(n_1746),
.B1(n_1858),
.B2(n_1850),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1913),
.Y(n_2000)
);

BUFx12f_ASAP7_75t_L g2001 ( 
.A(n_1945),
.Y(n_2001)
);

INVx8_ASAP7_75t_L g2002 ( 
.A(n_1950),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1959),
.B(n_1809),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1915),
.B(n_1873),
.Y(n_2004)
);

OAI31xp33_ASAP7_75t_L g2005 ( 
.A1(n_1944),
.A2(n_1858),
.A3(n_1763),
.B(n_1766),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1898),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1904),
.B(n_1913),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1944),
.A2(n_1756),
.B1(n_1754),
.B2(n_1763),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1913),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1929),
.A2(n_1756),
.B1(n_1766),
.B2(n_1760),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1897),
.B(n_1808),
.Y(n_2011)
);

OAI321xp33_ASAP7_75t_L g2012 ( 
.A1(n_1938),
.A2(n_1931),
.A3(n_1928),
.B1(n_1946),
.B2(n_1939),
.C(n_1954),
.Y(n_2012)
);

OAI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_1949),
.A2(n_1764),
.B1(n_1765),
.B2(n_1841),
.C(n_1892),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1910),
.Y(n_2014)
);

INVx3_ASAP7_75t_L g2015 ( 
.A(n_1923),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1907),
.Y(n_2016)
);

AOI33xp33_ASAP7_75t_L g2017 ( 
.A1(n_1947),
.A2(n_1744),
.A3(n_1887),
.B1(n_1757),
.B2(n_1767),
.B3(n_1797),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1925),
.B(n_1789),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1911),
.B(n_1744),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1923),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1939),
.B(n_1762),
.Y(n_2021)
);

NOR3xp33_ASAP7_75t_SL g2022 ( 
.A(n_1947),
.B(n_1886),
.C(n_1752),
.Y(n_2022)
);

NOR2x2_ASAP7_75t_L g2023 ( 
.A(n_1954),
.B(n_1823),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1896),
.B(n_1801),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1946),
.A2(n_1806),
.B1(n_1874),
.B2(n_1752),
.Y(n_2025)
);

OAI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1967),
.A2(n_1874),
.B1(n_1806),
.B2(n_1792),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_1939),
.B(n_1792),
.C(n_1954),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1927),
.Y(n_2028)
);

INVx5_ASAP7_75t_L g2029 ( 
.A(n_1916),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1927),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1930),
.B(n_1896),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1930),
.B(n_1914),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1903),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1914),
.B(n_1932),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1976),
.B(n_1977),
.Y(n_2035)
);

AOI222xp33_ASAP7_75t_L g2036 ( 
.A1(n_1938),
.A2(n_1969),
.B1(n_1962),
.B2(n_1970),
.C1(n_1971),
.C2(n_1980),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1976),
.B(n_1977),
.Y(n_2037)
);

OA222x2_ASAP7_75t_L g2038 ( 
.A1(n_1931),
.A2(n_1957),
.B1(n_1958),
.B2(n_1941),
.C1(n_1916),
.C2(n_1928),
.Y(n_2038)
);

AOI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_1941),
.A2(n_1963),
.B1(n_1936),
.B2(n_1975),
.C(n_1972),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_SL g2040 ( 
.A1(n_1970),
.A2(n_1962),
.B1(n_1969),
.B2(n_1929),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1980),
.A2(n_1967),
.B1(n_1929),
.B2(n_1926),
.Y(n_2041)
);

NAND2xp33_ASAP7_75t_R g2042 ( 
.A(n_1953),
.B(n_1929),
.Y(n_2042)
);

OAI31xp33_ASAP7_75t_SL g2043 ( 
.A1(n_1926),
.A2(n_1900),
.A3(n_1940),
.B(n_1904),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1910),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_1970),
.A2(n_1904),
.B1(n_1940),
.B2(n_1900),
.Y(n_2045)
);

NAND4xp25_ASAP7_75t_L g2046 ( 
.A(n_1934),
.B(n_1963),
.C(n_1975),
.D(n_1972),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1911),
.B(n_1933),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1918),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_R g2049 ( 
.A(n_1953),
.B(n_1973),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1903),
.Y(n_2050)
);

AOI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_1960),
.A2(n_1978),
.B1(n_1940),
.B2(n_1933),
.C(n_1942),
.Y(n_2051)
);

OAI221xp5_ASAP7_75t_SL g2052 ( 
.A1(n_1957),
.A2(n_1958),
.B1(n_1917),
.B2(n_1960),
.C(n_1916),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2033),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1983),
.B(n_1917),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_2014),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2035),
.B(n_1920),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_1985),
.B(n_1920),
.C(n_1966),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_1989),
.B(n_1982),
.C(n_1986),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2037),
.B(n_1919),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2015),
.B(n_1919),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2033),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2044),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2048),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2020),
.B(n_1942),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2020),
.B(n_1942),
.Y(n_2065)
);

CKINVDCx16_ASAP7_75t_R g2066 ( 
.A(n_2042),
.Y(n_2066)
);

NOR3xp33_ASAP7_75t_L g2067 ( 
.A(n_1997),
.B(n_1966),
.C(n_1968),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2050),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2047),
.B(n_1942),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2018),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2032),
.B(n_1901),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2020),
.B(n_1940),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2050),
.Y(n_2073)
);

OR2x6_ASAP7_75t_L g2074 ( 
.A(n_2002),
.B(n_1916),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_2007),
.B(n_1899),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2034),
.B(n_1902),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2006),
.B(n_1902),
.Y(n_2077)
);

NAND2xp67_ASAP7_75t_L g2078 ( 
.A(n_1981),
.B(n_1912),
.Y(n_2078)
);

AND2x4_ASAP7_75t_SL g2079 ( 
.A(n_1990),
.B(n_1904),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_SL g2080 ( 
.A(n_2027),
.B(n_2005),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1993),
.B(n_1922),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_2021),
.B(n_2046),
.Y(n_2082)
);

INVx4_ASAP7_75t_L g2083 ( 
.A(n_2002),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2007),
.B(n_2029),
.Y(n_2084)
);

AND2x4_ASAP7_75t_SL g2085 ( 
.A(n_1990),
.B(n_1916),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_2018),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2000),
.B(n_1948),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1994),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1994),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2000),
.B(n_1948),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2009),
.B(n_1948),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2009),
.B(n_1948),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2007),
.B(n_2028),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_1993),
.B(n_1906),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2019),
.B(n_1906),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2016),
.Y(n_2096)
);

OAI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_2080),
.A2(n_2058),
.B(n_2008),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_2066),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2082),
.B(n_2051),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2069),
.B(n_2031),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2069),
.B(n_2019),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2053),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2053),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_2055),
.Y(n_2104)
);

INVxp67_ASAP7_75t_SL g2105 ( 
.A(n_2082),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2071),
.B(n_2024),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2093),
.B(n_2066),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2068),
.Y(n_2108)
);

AOI32xp33_ASAP7_75t_L g2109 ( 
.A1(n_2080),
.A2(n_1984),
.A3(n_2012),
.B1(n_1995),
.B2(n_2041),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2071),
.B(n_2024),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_2084),
.B(n_2029),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_2083),
.B(n_2029),
.Y(n_2112)
);

NAND2xp33_ASAP7_75t_L g2113 ( 
.A(n_2058),
.B(n_2022),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2068),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_2056),
.Y(n_2115)
);

NOR2x1_ASAP7_75t_SL g2116 ( 
.A(n_2074),
.B(n_2029),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_2074),
.Y(n_2117)
);

BUFx2_ASAP7_75t_L g2118 ( 
.A(n_2074),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2093),
.B(n_2038),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2086),
.B(n_2076),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2055),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2061),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2062),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2093),
.B(n_2029),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2069),
.B(n_2016),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2094),
.B(n_2039),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2073),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2063),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2054),
.B(n_2003),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_2084),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2086),
.B(n_2003),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_2060),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2084),
.B(n_2030),
.Y(n_2133)
);

INVx4_ASAP7_75t_L g2134 ( 
.A(n_2083),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2054),
.B(n_1991),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2088),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2089),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2054),
.B(n_2075),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2075),
.B(n_1991),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2063),
.Y(n_2140)
);

AND2x4_ASAP7_75t_L g2141 ( 
.A(n_2084),
.B(n_2074),
.Y(n_2141)
);

INVx1_ASAP7_75t_SL g2142 ( 
.A(n_2062),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2089),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2096),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2075),
.B(n_2011),
.Y(n_2145)
);

INVx1_ASAP7_75t_SL g2146 ( 
.A(n_2094),
.Y(n_2146)
);

NOR2x1_ASAP7_75t_L g2147 ( 
.A(n_2083),
.B(n_2021),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2102),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2107),
.B(n_2084),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2105),
.B(n_2099),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2107),
.B(n_2084),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2098),
.B(n_2059),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_2101),
.B(n_2094),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_2097),
.B(n_2098),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2126),
.B(n_2067),
.Y(n_2155)
);

AOI31xp33_ASAP7_75t_L g2156 ( 
.A1(n_2097),
.A2(n_2057),
.A3(n_2040),
.B(n_2036),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2126),
.B(n_2067),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2129),
.B(n_2059),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_2134),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2131),
.B(n_2070),
.Y(n_2160)
);

INVxp67_ASAP7_75t_L g2161 ( 
.A(n_2104),
.Y(n_2161)
);

OR2x6_ASAP7_75t_L g2162 ( 
.A(n_2112),
.B(n_1990),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_2121),
.Y(n_2163)
);

AND2x4_ASAP7_75t_SL g2164 ( 
.A(n_2134),
.B(n_2111),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2129),
.B(n_2070),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2119),
.B(n_2059),
.Y(n_2166)
);

AND2x2_ASAP7_75t_SL g2167 ( 
.A(n_2113),
.B(n_2043),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2108),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2102),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2115),
.B(n_2087),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2106),
.B(n_2087),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2108),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_2141),
.B(n_2074),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2110),
.B(n_2004),
.Y(n_2174)
);

AOI221xp5_ASAP7_75t_L g2175 ( 
.A1(n_2109),
.A2(n_2057),
.B1(n_2052),
.B2(n_1996),
.C(n_1999),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2101),
.B(n_2095),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2146),
.B(n_2095),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2108),
.Y(n_2178)
);

NAND2x1_ASAP7_75t_L g2179 ( 
.A(n_2147),
.B(n_1955),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2146),
.B(n_2095),
.Y(n_2180)
);

BUFx2_ASAP7_75t_L g2181 ( 
.A(n_2147),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2114),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2103),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2135),
.B(n_2087),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2119),
.B(n_2072),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2135),
.B(n_2090),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2100),
.B(n_2081),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2145),
.B(n_2090),
.Y(n_2188)
);

INVxp67_ASAP7_75t_L g2189 ( 
.A(n_2123),
.Y(n_2189)
);

CKINVDCx16_ASAP7_75t_R g2190 ( 
.A(n_2134),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2100),
.B(n_2081),
.Y(n_2191)
);

INVx2_ASAP7_75t_SL g2192 ( 
.A(n_2130),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2145),
.B(n_2090),
.Y(n_2193)
);

INVxp67_ASAP7_75t_SL g2194 ( 
.A(n_2130),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2103),
.Y(n_2195)
);

CKINVDCx16_ASAP7_75t_R g2196 ( 
.A(n_2134),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2141),
.B(n_2072),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2120),
.B(n_2091),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2141),
.B(n_2072),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2109),
.B(n_2091),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2141),
.B(n_2075),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_2111),
.B(n_2026),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2139),
.B(n_2075),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2148),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2148),
.Y(n_2205)
);

OAI21xp33_ASAP7_75t_L g2206 ( 
.A1(n_2167),
.A2(n_2157),
.B(n_2155),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2169),
.Y(n_2207)
);

NOR2xp67_ASAP7_75t_L g2208 ( 
.A(n_2163),
.B(n_2130),
.Y(n_2208)
);

NOR2xp67_ASAP7_75t_L g2209 ( 
.A(n_2166),
.B(n_2130),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_2167),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_2167),
.A2(n_1990),
.B1(n_1998),
.B2(n_1988),
.Y(n_2211)
);

INVxp67_ASAP7_75t_SL g2212 ( 
.A(n_2179),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2154),
.B(n_2139),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2169),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_2164),
.B(n_2116),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_2150),
.B(n_1965),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2152),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2156),
.A2(n_1987),
.B1(n_2010),
.B2(n_2118),
.C(n_2117),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2183),
.Y(n_2219)
);

OAI31xp33_ASAP7_75t_SL g2220 ( 
.A1(n_2175),
.A2(n_2111),
.A3(n_2013),
.B(n_2142),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_2156),
.A2(n_2116),
.B(n_2111),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2183),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2195),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2200),
.B(n_2142),
.Y(n_2224)
);

OAI221xp5_ASAP7_75t_L g2225 ( 
.A1(n_2202),
.A2(n_2118),
.B1(n_2117),
.B2(n_2112),
.C(n_2045),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2166),
.B(n_2124),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2174),
.B(n_2152),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_2179),
.Y(n_2228)
);

OAI211xp5_ASAP7_75t_L g2229 ( 
.A1(n_2181),
.A2(n_2065),
.B(n_2064),
.C(n_2025),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2149),
.B(n_2124),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2195),
.Y(n_2231)
);

NAND2x1p5_ASAP7_75t_L g2232 ( 
.A(n_2181),
.B(n_2083),
.Y(n_2232)
);

OAI21xp33_ASAP7_75t_SL g2233 ( 
.A1(n_2149),
.A2(n_2132),
.B(n_2138),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2151),
.B(n_2138),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2165),
.B(n_2125),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2190),
.B(n_2112),
.Y(n_2236)
);

NOR2xp67_ASAP7_75t_L g2237 ( 
.A(n_2161),
.B(n_2132),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_2164),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2189),
.B(n_2158),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2184),
.B(n_2125),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2151),
.B(n_2133),
.Y(n_2241)
);

OAI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_2162),
.A2(n_2049),
.B1(n_2074),
.B2(n_2083),
.Y(n_2242)
);

OAI21xp5_ASAP7_75t_SL g2243 ( 
.A1(n_2164),
.A2(n_2085),
.B(n_2079),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2158),
.B(n_2133),
.Y(n_2244)
);

OAI211xp5_ASAP7_75t_L g2245 ( 
.A1(n_2159),
.A2(n_2065),
.B(n_2064),
.C(n_2092),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_2215),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_2206),
.A2(n_2162),
.B(n_2159),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2220),
.B(n_2190),
.Y(n_2248)
);

OAI32xp33_ASAP7_75t_L g2249 ( 
.A1(n_2210),
.A2(n_2196),
.A3(n_2180),
.B1(n_2177),
.B2(n_2153),
.Y(n_2249)
);

AOI21xp33_ASAP7_75t_L g2250 ( 
.A1(n_2212),
.A2(n_2162),
.B(n_2194),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2204),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2218),
.B(n_2196),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2204),
.Y(n_2253)
);

OAI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2221),
.A2(n_2211),
.B(n_2224),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2205),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2227),
.B(n_2185),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2238),
.Y(n_2257)
);

O2A1O1Ixp33_ASAP7_75t_L g2258 ( 
.A1(n_2225),
.A2(n_2162),
.B(n_2160),
.C(n_2170),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2216),
.B(n_2185),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2217),
.B(n_2186),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2213),
.A2(n_1988),
.B1(n_2162),
.B2(n_2173),
.Y(n_2261)
);

NOR3xp33_ASAP7_75t_SL g2262 ( 
.A(n_2236),
.B(n_2243),
.C(n_2242),
.Y(n_2262)
);

O2A1O1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_2229),
.A2(n_2192),
.B(n_2180),
.C(n_2177),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_2217),
.Y(n_2264)
);

OR2x2_ASAP7_75t_L g2265 ( 
.A(n_2239),
.B(n_2153),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2226),
.B(n_2188),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2237),
.A2(n_2173),
.B1(n_1988),
.B2(n_2085),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2205),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2226),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2208),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2215),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2215),
.A2(n_2173),
.B1(n_2085),
.B2(n_2197),
.Y(n_2272)
);

AOI32xp33_ASAP7_75t_L g2273 ( 
.A1(n_2230),
.A2(n_2233),
.A3(n_2228),
.B1(n_2234),
.B2(n_2241),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2207),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2230),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2234),
.B(n_2193),
.Y(n_2276)
);

CKINVDCx16_ASAP7_75t_R g2277 ( 
.A(n_2257),
.Y(n_2277)
);

INVxp67_ASAP7_75t_L g2278 ( 
.A(n_2246),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2264),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2271),
.B(n_2241),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2248),
.B(n_2228),
.Y(n_2281)
);

OAI31xp33_ASAP7_75t_L g2282 ( 
.A1(n_2252),
.A2(n_2232),
.A3(n_2245),
.B(n_2228),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2264),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2246),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2251),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2253),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2275),
.B(n_2232),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2255),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2268),
.Y(n_2289)
);

XNOR2xp5_ASAP7_75t_L g2290 ( 
.A(n_2262),
.B(n_2247),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_2254),
.A2(n_2232),
.B(n_2209),
.Y(n_2291)
);

INVxp67_ASAP7_75t_L g2292 ( 
.A(n_2259),
.Y(n_2292)
);

XNOR2xp5_ASAP7_75t_L g2293 ( 
.A(n_2272),
.B(n_1965),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2258),
.B(n_2261),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2275),
.B(n_2244),
.Y(n_2295)
);

NAND2xp33_ASAP7_75t_R g2296 ( 
.A(n_2265),
.B(n_1992),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_SL g2297 ( 
.A(n_2261),
.B(n_2017),
.Y(n_2297)
);

NAND2xp33_ASAP7_75t_R g2298 ( 
.A(n_2265),
.B(n_2173),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2249),
.A2(n_2223),
.B(n_2222),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_2269),
.Y(n_2300)
);

NAND3xp33_ASAP7_75t_L g2301 ( 
.A(n_2294),
.B(n_2250),
.C(n_2270),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2277),
.B(n_2256),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2282),
.B(n_2267),
.Y(n_2303)
);

NOR2x1_ASAP7_75t_L g2304 ( 
.A(n_2284),
.B(n_2274),
.Y(n_2304)
);

NAND4xp75_ASAP7_75t_L g2305 ( 
.A(n_2294),
.B(n_2269),
.C(n_2266),
.D(n_2276),
.Y(n_2305)
);

NAND3xp33_ASAP7_75t_L g2306 ( 
.A(n_2297),
.B(n_2273),
.C(n_2263),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2279),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2297),
.A2(n_2290),
.B(n_2281),
.Y(n_2308)
);

AOI211xp5_ASAP7_75t_L g2309 ( 
.A1(n_2290),
.A2(n_2260),
.B(n_2207),
.C(n_2214),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2284),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2281),
.A2(n_2260),
.B(n_2219),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2283),
.Y(n_2312)
);

AO21x1_ASAP7_75t_L g2313 ( 
.A1(n_2299),
.A2(n_2219),
.B(n_2214),
.Y(n_2313)
);

NAND4xp25_ASAP7_75t_L g2314 ( 
.A(n_2296),
.B(n_2231),
.C(n_2235),
.D(n_2017),
.Y(n_2314)
);

OAI211xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2292),
.A2(n_2231),
.B(n_2235),
.C(n_2240),
.Y(n_2315)
);

NOR3xp33_ASAP7_75t_L g2316 ( 
.A(n_2301),
.B(n_2278),
.C(n_2300),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_R g2317 ( 
.A(n_2308),
.B(n_2291),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_R g2318 ( 
.A(n_2302),
.B(n_2298),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2304),
.Y(n_2319)
);

AOI211xp5_ASAP7_75t_L g2320 ( 
.A1(n_2306),
.A2(n_2293),
.B(n_2280),
.C(n_2287),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2303),
.A2(n_2293),
.B1(n_2295),
.B2(n_2287),
.Y(n_2321)
);

NOR3xp33_ASAP7_75t_L g2322 ( 
.A(n_2309),
.B(n_2305),
.C(n_2314),
.Y(n_2322)
);

OAI211xp5_ASAP7_75t_L g2323 ( 
.A1(n_2309),
.A2(n_2289),
.B(n_2288),
.C(n_2286),
.Y(n_2323)
);

AOI211xp5_ASAP7_75t_L g2324 ( 
.A1(n_2313),
.A2(n_2285),
.B(n_2240),
.C(n_2192),
.Y(n_2324)
);

AOI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2311),
.A2(n_2244),
.B(n_2199),
.C(n_2197),
.Y(n_2325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2326 ( 
.A1(n_2307),
.A2(n_2198),
.B(n_2171),
.C(n_2137),
.D(n_2122),
.Y(n_2326)
);

AOI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_2312),
.A2(n_2182),
.B(n_2168),
.Y(n_2327)
);

AOI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2315),
.A2(n_2199),
.B(n_2201),
.C(n_2176),
.Y(n_2328)
);

AOI211xp5_ASAP7_75t_L g2329 ( 
.A1(n_2310),
.A2(n_2201),
.B(n_2176),
.C(n_2191),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2324),
.A2(n_2178),
.B(n_2182),
.Y(n_2330)
);

NOR3xp33_ASAP7_75t_L g2331 ( 
.A(n_2322),
.B(n_2316),
.C(n_2320),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2317),
.A2(n_2203),
.B1(n_2085),
.B2(n_2168),
.Y(n_2332)
);

OAI22xp33_ASAP7_75t_SL g2333 ( 
.A1(n_2319),
.A2(n_2326),
.B1(n_2318),
.B2(n_2323),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_R g2334 ( 
.A(n_2321),
.B(n_1979),
.Y(n_2334)
);

NOR3xp33_ASAP7_75t_L g2335 ( 
.A(n_2329),
.B(n_2172),
.C(n_2178),
.Y(n_2335)
);

INVx2_ASAP7_75t_SL g2336 ( 
.A(n_2325),
.Y(n_2336)
);

AOI22x1_ASAP7_75t_L g2337 ( 
.A1(n_2328),
.A2(n_2172),
.B1(n_2191),
.B2(n_2187),
.Y(n_2337)
);

NOR3x1_ASAP7_75t_L g2338 ( 
.A(n_2336),
.B(n_2327),
.C(n_2187),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2333),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2331),
.B(n_2203),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2332),
.B(n_2064),
.C(n_2065),
.Y(n_2341)
);

NOR3x1_ASAP7_75t_L g2342 ( 
.A(n_2334),
.B(n_2023),
.C(n_2081),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2330),
.B(n_2077),
.Y(n_2343)
);

OAI221xp5_ASAP7_75t_L g2344 ( 
.A1(n_2337),
.A2(n_2074),
.B1(n_1979),
.B2(n_1945),
.C(n_1951),
.Y(n_2344)
);

AOI221xp5_ASAP7_75t_L g2345 ( 
.A1(n_2335),
.A2(n_2133),
.B1(n_2091),
.B2(n_2092),
.C(n_2137),
.Y(n_2345)
);

NAND3xp33_ASAP7_75t_L g2346 ( 
.A(n_2339),
.B(n_2092),
.C(n_2128),
.Y(n_2346)
);

NAND5xp2_ASAP7_75t_L g2347 ( 
.A(n_2340),
.B(n_1951),
.C(n_1945),
.D(n_2023),
.E(n_1961),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2341),
.A2(n_2079),
.B1(n_2001),
.B2(n_2002),
.Y(n_2348)
);

XOR2xp5_ASAP7_75t_L g2349 ( 
.A(n_2343),
.B(n_1951),
.Y(n_2349)
);

O2A1O1Ixp5_ASAP7_75t_L g2350 ( 
.A1(n_2338),
.A2(n_2128),
.B(n_2140),
.C(n_2114),
.Y(n_2350)
);

XOR2xp5_ASAP7_75t_L g2351 ( 
.A(n_2342),
.B(n_1943),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2351),
.B(n_2345),
.Y(n_2352)
);

OAI321xp33_ASAP7_75t_L g2353 ( 
.A1(n_2346),
.A2(n_2344),
.A3(n_1952),
.B1(n_1968),
.B2(n_2056),
.C(n_2136),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2347),
.B(n_2349),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_2348),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2352),
.Y(n_2356)
);

OAI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2356),
.A2(n_2354),
.B(n_2350),
.Y(n_2357)
);

INVx1_ASAP7_75t_SL g2358 ( 
.A(n_2357),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2357),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2359),
.Y(n_2360)
);

OAI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2358),
.A2(n_2355),
.B(n_2353),
.Y(n_2361)
);

OAI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2361),
.A2(n_2128),
.B(n_2140),
.Y(n_2362)
);

AOI22xp33_ASAP7_75t_R g2363 ( 
.A1(n_2360),
.A2(n_2140),
.B1(n_2114),
.B2(n_2143),
.Y(n_2363)
);

NAND3xp33_ASAP7_75t_L g2364 ( 
.A(n_2362),
.B(n_2127),
.C(n_2143),
.Y(n_2364)
);

OAI221xp5_ASAP7_75t_R g2365 ( 
.A1(n_2364),
.A2(n_2363),
.B1(n_2002),
.B2(n_1955),
.C(n_2078),
.Y(n_2365)
);

AOI211xp5_ASAP7_75t_L g2366 ( 
.A1(n_2365),
.A2(n_2144),
.B(n_2136),
.C(n_2122),
.Y(n_2366)
);


endmodule