module fake_jpeg_16963_n_35 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_35);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_32;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_24)
);

AO21x2_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_18),
.B(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_12),
.Y(n_31)
);

OAI322xp33_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_25),
.A3(n_7),
.B1(n_10),
.B2(n_11),
.C1(n_6),
.C2(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_29),
.B(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_27),
.Y(n_34)
);

AOI21x1_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_28),
.B(n_15),
.Y(n_35)
);


endmodule