module real_jpeg_25051_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_0),
.A2(n_38),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_0),
.A2(n_47),
.B1(n_65),
.B2(n_67),
.Y(n_168)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_37),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_50),
.C(n_52),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_2),
.A2(n_38),
.B1(n_41),
.B2(n_110),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_105),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_110),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_65),
.C(n_77),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_2),
.A2(n_68),
.B(n_217),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_4),
.A2(n_27),
.B1(n_38),
.B2(n_41),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_4),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_27),
.B1(n_65),
.B2(n_67),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_65),
.B1(n_67),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_8),
.A2(n_43),
.B1(n_65),
.B2(n_67),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_11),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_65),
.B1(n_67),
.B2(n_82),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_38),
.B1(n_41),
.B2(n_82),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_14),
.A2(n_65),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_71),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_15),
.A2(n_38),
.B1(n_41),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_15),
.A2(n_56),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_15),
.A2(n_56),
.B1(n_65),
.B2(n_67),
.Y(n_187)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_142),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_20),
.B(n_118),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_93),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_25),
.B(n_44),
.C(n_60),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_37),
.B2(n_42),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_26),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_28),
.B(n_35),
.C(n_41),
.Y(n_112)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_32),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_32),
.A2(n_139),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_34),
.A2(n_38),
.B(n_109),
.C(n_112),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_36),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_36),
.B(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_38),
.B(n_183),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_42),
.Y(n_136)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_46),
.A2(n_48),
.B1(n_58),
.B2(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_48),
.A2(n_54),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_50),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_50),
.B(n_225),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_55),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_57),
.A2(n_103),
.B1(n_105),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_58),
.A2(n_104),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_61),
.B(n_73),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_63),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_69),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_67),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_67),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_70),
.B1(n_72),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_68),
.A2(n_85),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_68),
.A2(n_72),
.B1(n_116),
.B2(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_68),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_68),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_69),
.Y(n_240)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_72),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_74),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_74),
.A2(n_205),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_89),
.B1(n_90),
.B2(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_75),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_75),
.A2(n_90),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_79),
.A2(n_80),
.B(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_79),
.A2(n_155),
.B(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_79),
.B(n_110),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_83),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_90),
.B(n_156),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_93),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.C(n_106),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_101),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_109),
.B(n_110),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_106),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_110),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_114),
.A2(n_229),
.B1(n_231),
.B2(n_233),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_141),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_129),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_140),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_175),
.B(n_265),
.C(n_270),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_169),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_169),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_159),
.C(n_162),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_147),
.A2(n_148),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_153),
.C(n_157),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_162),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_170),
.B(n_173),
.C(n_174),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_258),
.B(n_264),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_206),
.B(n_257),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_195),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_180),
.B(n_195),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.C(n_192),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_196),
.B(n_202),
.C(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_251),
.B(n_256),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_226),
.B(n_250),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_220),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_236),
.B(n_249),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_234),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_242),
.B(n_248),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);


endmodule