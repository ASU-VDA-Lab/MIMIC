module fake_jpeg_12314_n_649 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_649);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_649;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_625;
wire n_312;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_3),
.B(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_SL g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_1),
.B(n_6),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_84),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_34),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_102),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_10),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_41),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_121),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_113),
.Y(n_129)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_115),
.A2(n_29),
.B1(n_33),
.B2(n_55),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_116),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_9),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_36),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_31),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_127),
.B(n_146),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_80),
.A2(n_40),
.B1(n_21),
.B2(n_54),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_130),
.A2(n_203),
.B1(n_73),
.B2(n_68),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_35),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_132),
.B(n_156),
.Y(n_243)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_20),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_81),
.A2(n_28),
.B1(n_54),
.B2(n_50),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_150),
.A2(n_50),
.B1(n_116),
.B2(n_74),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_41),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_162),
.B(n_167),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_90),
.B(n_41),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_164),
.B(n_181),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_42),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_172),
.B(n_180),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_58),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_58),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_201),
.B1(n_23),
.B2(n_32),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_90),
.B(n_56),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_184),
.B(n_186),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_110),
.B(n_33),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_61),
.A2(n_40),
.B1(n_28),
.B2(n_29),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_50),
.B1(n_117),
.B2(n_109),
.Y(n_218)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_67),
.Y(n_196)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_110),
.B(n_56),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_200),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_83),
.B(n_23),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_88),
.A2(n_21),
.B1(n_47),
.B2(n_43),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_116),
.A2(n_40),
.B1(n_21),
.B2(n_46),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_206),
.B(n_222),
.Y(n_317)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_207),
.Y(n_328)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_153),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_209),
.Y(n_288)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_211),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_96),
.C(n_118),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_212),
.B(n_193),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_214),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_228),
.Y(n_286)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_216),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_130),
.A2(n_203),
.B1(n_204),
.B2(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_219),
.A2(n_141),
.B1(n_49),
.B2(n_6),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_220),
.Y(n_325)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_223),
.A2(n_225),
.B1(n_234),
.B2(n_239),
.Y(n_332)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_224),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_155),
.A2(n_76),
.B1(n_66),
.B2(n_62),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_124),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_226),
.Y(n_290)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_151),
.A2(n_94),
.B1(n_93),
.B2(n_107),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_128),
.Y(n_230)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_231),
.B(n_255),
.Y(n_320)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_159),
.Y(n_232)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_155),
.A2(n_72),
.B1(n_64),
.B2(n_69),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_235),
.Y(n_292)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_133),
.Y(n_238)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_126),
.A2(n_68),
.B1(n_103),
.B2(n_101),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_240),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_189),
.A2(n_97),
.B1(n_98),
.B2(n_113),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_247),
.B1(n_39),
.B2(n_141),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_138),
.Y(n_244)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_147),
.B(n_55),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_245),
.B(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_161),
.A2(n_43),
.B1(n_36),
.B2(n_39),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_150),
.A2(n_120),
.B1(n_85),
.B2(n_50),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_261),
.B1(n_223),
.B2(n_225),
.Y(n_293)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_147),
.B(n_47),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_128),
.Y(n_253)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_181),
.A2(n_50),
.B(n_42),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_254),
.A2(n_49),
.B(n_2),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_184),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_131),
.Y(n_256)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_256),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_156),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_257),
.B(n_259),
.Y(n_330)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_258),
.Y(n_336)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g260 ( 
.A1(n_150),
.A2(n_178),
.B1(n_187),
.B2(n_195),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_269),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_148),
.A2(n_49),
.B1(n_26),
.B2(n_50),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_197),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_266),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_263),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_276),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_186),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_158),
.A2(n_139),
.B1(n_137),
.B2(n_170),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_270),
.B(n_272),
.Y(n_341)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_171),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_161),
.B(n_32),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_273),
.B(n_274),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_188),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_275),
.B(n_279),
.Y(n_304)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_149),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_278),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_129),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_149),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_271),
.B(n_169),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_281),
.B(n_291),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_213),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_296),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_267),
.B(n_169),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_293),
.A2(n_300),
.B1(n_302),
.B2(n_306),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_172),
.B(n_164),
.C(n_198),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_298),
.B(n_311),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_248),
.A2(n_219),
.B1(n_254),
.B2(n_249),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_233),
.B(n_157),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_316),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_260),
.A2(n_163),
.B1(n_168),
.B2(n_191),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_260),
.A2(n_191),
.B1(n_188),
.B2(n_154),
.Y(n_306)
);

FAx1_ASAP7_75t_L g308 ( 
.A(n_212),
.B(n_152),
.CI(n_176),
.CON(n_308),
.SN(n_308)
);

XOR2x2_ASAP7_75t_SL g383 ( 
.A(n_308),
.B(n_293),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_243),
.B(n_183),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_205),
.B(n_49),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_318),
.B(n_322),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_319),
.A2(n_327),
.B(n_270),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_194),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_216),
.B(n_2),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_2),
.Y(n_350)
);

NAND2x1_ASAP7_75t_SL g327 ( 
.A(n_237),
.B(n_2),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_334),
.B(n_8),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_241),
.A2(n_49),
.B1(n_5),
.B2(n_6),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_338),
.A2(n_339),
.B1(n_253),
.B2(n_230),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_260),
.A2(n_11),
.B1(n_5),
.B2(n_7),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_215),
.B(n_12),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_234),
.C(n_269),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_239),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_343)
);

AOI22x1_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_244),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_347),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_345),
.B(n_390),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_286),
.A2(n_232),
.B1(n_227),
.B2(n_258),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_346),
.A2(n_352),
.B1(n_364),
.B2(n_371),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_238),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_350),
.B(n_389),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_208),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_355),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_286),
.A2(n_342),
.B1(n_284),
.B2(n_300),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_291),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_357),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_250),
.C(n_240),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_359),
.C(n_362),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_224),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_214),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_370),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_358),
.A2(n_387),
.B(n_376),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_301),
.B(n_274),
.C(n_264),
.Y(n_359)
);

OAI21xp33_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_8),
.B(n_9),
.Y(n_361)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_386),
.B(n_388),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_226),
.C(n_229),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_299),
.B(n_259),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_298),
.A2(n_207),
.B1(n_265),
.B2(n_278),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_256),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_375),
.Y(n_419)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_327),
.B(n_9),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_376),
.B(n_381),
.Y(n_430)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_378),
.Y(n_434)
);

AOI32xp33_ASAP7_75t_L g379 ( 
.A1(n_308),
.A2(n_236),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_379),
.A2(n_383),
.B(n_329),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_332),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_380),
.A2(n_384),
.B1(n_305),
.B2(n_303),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_295),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_327),
.B(n_15),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_329),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_304),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_322),
.A2(n_15),
.B(n_308),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_280),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_292),
.Y(n_389)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_340),
.B(n_15),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_343),
.A2(n_324),
.B1(n_297),
.B2(n_336),
.Y(n_391)
);

BUFx5_ASAP7_75t_L g421 ( 
.A(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_392),
.B(n_393),
.Y(n_401)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_307),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_395),
.A2(n_399),
.B(n_413),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_348),
.A2(n_330),
.B(n_296),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_367),
.A2(n_338),
.B1(n_283),
.B2(n_303),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_400),
.A2(n_437),
.B1(n_371),
.B2(n_346),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_354),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_404),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_370),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_378),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_407),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_326),
.C(n_314),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_369),
.C(n_374),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_356),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_360),
.B(n_314),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_410),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_420),
.Y(n_443)
);

OA21x2_ASAP7_75t_SL g412 ( 
.A1(n_348),
.A2(n_326),
.B(n_305),
.Y(n_412)
);

AOI21xp33_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_372),
.B(n_388),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_387),
.A2(n_283),
.B(n_325),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_414),
.B(n_431),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_368),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_393),
.Y(n_467)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_360),
.A2(n_336),
.A3(n_297),
.B1(n_324),
.B2(n_289),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_358),
.A2(n_325),
.B(n_333),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_423),
.A2(n_432),
.B(n_435),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_352),
.A2(n_295),
.B1(n_328),
.B2(n_285),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_424),
.A2(n_425),
.B1(n_381),
.B2(n_382),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_377),
.A2(n_328),
.B1(n_285),
.B2(n_329),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_349),
.B(n_289),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_427),
.B(n_386),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_355),
.A2(n_333),
.B(n_280),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_377),
.A2(n_280),
.B(n_294),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_367),
.A2(n_290),
.B1(n_310),
.B2(n_321),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_429),
.B(n_349),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_440),
.B(n_464),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_441),
.B(n_454),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_444),
.A2(n_447),
.B1(n_425),
.B2(n_394),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g445 ( 
.A(n_415),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_445),
.B(n_419),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_350),
.Y(n_446)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_400),
.A2(n_377),
.B1(n_364),
.B2(n_345),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_383),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_464),
.C(n_472),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g511 ( 
.A(n_451),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_426),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_452),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_396),
.B(n_359),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_362),
.Y(n_456)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_458),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_415),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_469),
.Y(n_481)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_462),
.A2(n_437),
.B1(n_435),
.B2(n_432),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_396),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_463),
.A2(n_470),
.B1(n_471),
.B2(n_403),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_399),
.B(n_390),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_424),
.A2(n_379),
.B(n_385),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_465),
.A2(n_476),
.B(n_413),
.Y(n_488)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_467),
.Y(n_478)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_422),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_468),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_410),
.B(n_392),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_433),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_402),
.B(n_390),
.C(n_389),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_473),
.B(n_406),
.C(n_398),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_365),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_474),
.B(n_416),
.Y(n_490)
);

OA22x2_ASAP7_75t_L g475 ( 
.A1(n_408),
.A2(n_384),
.B1(n_366),
.B2(n_363),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_421),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_423),
.A2(n_384),
.B(n_337),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_447),
.A2(n_408),
.B1(n_404),
.B2(n_397),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_477),
.A2(n_484),
.B1(n_439),
.B2(n_449),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_480),
.B(n_451),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_394),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_504),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_488),
.A2(n_492),
.B(n_495),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_489),
.A2(n_444),
.B1(n_475),
.B2(n_431),
.Y(n_541)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_455),
.A2(n_453),
.B(n_443),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_443),
.A2(n_411),
.B(n_412),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_497),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_460),
.Y(n_497)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_498),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_463),
.A2(n_409),
.B1(n_398),
.B2(n_395),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_438),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_501),
.B(n_459),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_469),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_502),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_472),
.C(n_473),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_457),
.A2(n_409),
.B1(n_397),
.B2(n_430),
.Y(n_505)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_505),
.Y(n_532)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_506),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_440),
.B(n_414),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_430),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_495),
.A2(n_455),
.B(n_476),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_513),
.A2(n_495),
.B(n_481),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_514),
.B(n_524),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_515),
.A2(n_507),
.B1(n_509),
.B2(n_510),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_516),
.B(n_521),
.C(n_531),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_478),
.B(n_454),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_517),
.B(n_526),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_477),
.A2(n_462),
.B1(n_453),
.B2(n_456),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_518),
.A2(n_489),
.B1(n_488),
.B2(n_487),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_442),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_520),
.B(n_527),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_442),
.C(n_446),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_523),
.B(n_510),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_478),
.B(n_428),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_486),
.B(n_417),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_428),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_530),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_403),
.C(n_468),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_466),
.C(n_461),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_533),
.B(n_537),
.Y(n_550)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_535),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_508),
.B(n_504),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_538),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_493),
.B(n_470),
.C(n_458),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_492),
.B(n_420),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_482),
.B(n_471),
.C(n_465),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_542),
.Y(n_556)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_541),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_482),
.B(n_436),
.C(n_434),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_544),
.A2(n_547),
.B1(n_549),
.B2(n_552),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_528),
.A2(n_487),
.B1(n_502),
.B2(n_483),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_548),
.B(n_565),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_528),
.A2(n_483),
.B1(n_481),
.B2(n_491),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_515),
.A2(n_518),
.B1(n_532),
.B2(n_519),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_512),
.B(n_497),
.Y(n_554)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_554),
.Y(n_574)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_539),
.Y(n_558)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_558),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_522),
.B(n_496),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_563),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_540),
.A2(n_491),
.B1(n_496),
.B2(n_507),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_560),
.Y(n_579)
);

BUFx24_ASAP7_75t_SL g561 ( 
.A(n_520),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_309),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_539),
.B(n_537),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_562),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_564),
.B(n_566),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_513),
.A2(n_475),
.B(n_500),
.C(n_509),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_567),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_533),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_521),
.B(n_500),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_554),
.A2(n_543),
.B1(n_568),
.B2(n_553),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_571),
.B(n_572),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_555),
.B(n_531),
.C(n_516),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_522),
.C(n_527),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_573),
.B(n_583),
.C(n_586),
.Y(n_591)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_575),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_553),
.A2(n_529),
.B1(n_538),
.B2(n_525),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_576),
.Y(n_597)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_544),
.A2(n_525),
.B(n_479),
.Y(n_577)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_577),
.Y(n_607)
);

MAJx2_ASAP7_75t_L g578 ( 
.A(n_545),
.B(n_536),
.C(n_523),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_578),
.B(n_589),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_543),
.A2(n_475),
.B1(n_542),
.B2(n_479),
.Y(n_581)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_581),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_546),
.B(n_534),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_582),
.B(n_550),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_494),
.C(n_506),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_584),
.B(n_313),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_545),
.B(n_494),
.C(n_434),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_559),
.B(n_421),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_556),
.B(n_405),
.C(n_321),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_590),
.B(n_562),
.C(n_558),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_592),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_574),
.A2(n_585),
.B1(n_588),
.B2(n_579),
.Y(n_595)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_595),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_596),
.B(n_606),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_572),
.B(n_560),
.C(n_552),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_599),
.A2(n_600),
.B(n_601),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_586),
.B(n_551),
.C(n_563),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_575),
.A2(n_548),
.B(n_549),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_551),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_587),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_570),
.B(n_557),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_603),
.A2(n_604),
.B(n_290),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_575),
.A2(n_547),
.B(n_426),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_569),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_608),
.A2(n_590),
.B1(n_578),
.B2(n_309),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_573),
.C(n_588),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_609),
.B(n_611),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_591),
.B(n_583),
.C(n_580),
.Y(n_611)
);

FAx1_ASAP7_75t_SL g613 ( 
.A(n_597),
.B(n_577),
.CI(n_580),
.CON(n_613),
.SN(n_613)
);

NOR3x1_ASAP7_75t_SL g628 ( 
.A(n_613),
.B(n_607),
.C(n_605),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_598),
.A2(n_577),
.B1(n_576),
.B2(n_587),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_614),
.A2(n_619),
.B1(n_622),
.B2(n_610),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_615),
.A2(n_621),
.B(n_604),
.Y(n_626)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_616),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_592),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_599),
.B(n_380),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_620),
.B(n_603),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_593),
.A2(n_310),
.B(n_337),
.Y(n_621)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_624),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_613),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_626),
.A2(n_627),
.B(n_630),
.Y(n_636)
);

NOR2x1_ASAP7_75t_L g627 ( 
.A(n_614),
.B(n_605),
.Y(n_627)
);

XNOR2x2_ASAP7_75t_SL g638 ( 
.A(n_628),
.B(n_631),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_612),
.A2(n_607),
.B(n_601),
.Y(n_630)
);

OAI21xp33_ASAP7_75t_L g631 ( 
.A1(n_617),
.A2(n_594),
.B(n_602),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_610),
.B(n_594),
.Y(n_632)
);

AOI21xp33_ASAP7_75t_L g633 ( 
.A1(n_632),
.A2(n_619),
.B(n_615),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_633),
.B(n_635),
.Y(n_641)
);

AOI21x1_ASAP7_75t_L g642 ( 
.A1(n_634),
.A2(n_636),
.B(n_627),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_609),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_629),
.B(n_611),
.C(n_620),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_637),
.B(n_618),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_628),
.C(n_600),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_640),
.A2(n_643),
.B(n_638),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_642),
.A2(n_638),
.B(n_631),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_644),
.A2(n_645),
.B(n_641),
.Y(n_646)
);

AOI21x1_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_613),
.B(n_312),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_312),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_648),
.Y(n_649)
);


endmodule