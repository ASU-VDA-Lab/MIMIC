module fake_aes_1273_n_1211 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1211);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1211;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_353;
wire n_564;
wire n_1122;
wire n_779;
wire n_993;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1078;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_1204;
wire n_652;
wire n_968;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1188;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1159;
wire n_1011;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_1132;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_1160;
wire n_1184;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_1046;
wire n_460;
wire n_1183;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_1106;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_1206;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_1178;
wire n_1209;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1210;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_950;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_1199;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_1110;
wire n_327;
wire n_944;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_1208;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_582;
wire n_378;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_335;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1117;
wire n_859;
wire n_1007;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_1137;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_819;
wire n_405;
wire n_772;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
INVx2_ASAP7_75t_L g291 ( .A(n_272), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_170), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_124), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_231), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_81), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_179), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_217), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_239), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_238), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_268), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_8), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_155), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_2), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_156), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_197), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_254), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_224), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_148), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_276), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_215), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_161), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_235), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_263), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_53), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_109), .Y(n_315) );
BUFx10_ASAP7_75t_L g316 ( .A(n_194), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_36), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_283), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_91), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_265), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_216), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_122), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_38), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_165), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_101), .Y(n_326) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_267), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_25), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_198), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_28), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_38), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_85), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_74), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g335 ( .A(n_209), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_142), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_221), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_259), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_172), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_252), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_34), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_75), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_89), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_81), .Y(n_344) );
CKINVDCx11_ASAP7_75t_R g345 ( .A(n_126), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_54), .Y(n_346) );
BUFx5_ASAP7_75t_L g347 ( .A(n_176), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_66), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_162), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_24), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_159), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_18), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_187), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_182), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_140), .Y(n_355) );
CKINVDCx14_ASAP7_75t_R g356 ( .A(n_110), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_145), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_34), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_290), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_270), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_122), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_37), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_250), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_97), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_274), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_53), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_285), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_120), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_52), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_39), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_110), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_26), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_6), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_208), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_99), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_284), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_286), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_150), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_43), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_87), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_27), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_147), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_183), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_160), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_20), .B(n_173), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_185), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_61), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_200), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_226), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_257), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_152), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_188), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_78), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_178), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_211), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_94), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_220), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_73), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_202), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_99), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_42), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_229), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_149), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_78), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_207), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_23), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_255), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_225), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_249), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_280), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_234), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_251), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_132), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_223), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_143), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_46), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_3), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_109), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_236), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_50), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_82), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_32), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_279), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_46), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_62), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_210), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_196), .B(n_134), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_193), .Y(n_428) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_51), .B(n_55), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_49), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_213), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_144), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_189), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_20), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_219), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_146), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_16), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_123), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_151), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_44), .Y(n_440) );
CKINVDCx11_ASAP7_75t_R g441 ( .A(n_171), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_65), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_37), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_127), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_260), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_264), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_240), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g448 ( .A(n_247), .B(n_117), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_89), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_29), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_382), .B(n_0), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_356), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_361), .B(n_1), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_382), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_361), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_356), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_297), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_297), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_315), .A2(n_7), .B1(n_4), .B2(n_5), .Y(n_460) );
INVx4_ASAP7_75t_L g461 ( .A(n_294), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_297), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_347), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_361), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_347), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_347), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_315), .A2(n_10), .B1(n_7), .B2(n_9), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_297), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_296), .B(n_9), .Y(n_469) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_335), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_335), .B(n_10), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_345), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_347), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_295), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_347), .Y(n_475) );
OAI21x1_ASAP7_75t_L g476 ( .A1(n_291), .A2(n_138), .B(n_137), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_303), .B(n_11), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_295), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_316), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_424), .B(n_11), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_355), .B(n_12), .Y(n_481) );
BUFx8_ASAP7_75t_L g482 ( .A(n_347), .Y(n_482) );
INVx4_ASAP7_75t_L g483 ( .A(n_316), .Y(n_483) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_291), .A2(n_141), .B(n_139), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_317), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_485) );
BUFx8_ASAP7_75t_L g486 ( .A(n_347), .Y(n_486) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_326), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_487) );
OAI21x1_ASAP7_75t_L g488 ( .A1(n_311), .A2(n_395), .B(n_349), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_323), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_449), .B(n_15), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_326), .A2(n_18), .B1(n_16), .B2(n_17), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_309), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_327), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_488), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_482), .Y(n_495) );
AO22x2_ASAP7_75t_L g496 ( .A1(n_456), .A2(n_427), .B1(n_385), .B2(n_349), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_455), .B(n_325), .Y(n_497) );
BUFx6f_ASAP7_75t_SL g498 ( .A(n_483), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_482), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_488), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_483), .B(n_316), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_463), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_483), .B(n_300), .Y(n_504) );
BUFx4f_ASAP7_75t_L g505 ( .A(n_453), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_455), .B(n_394), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_461), .B(n_322), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_457), .Y(n_509) );
CKINVDCx6p67_ASAP7_75t_R g510 ( .A(n_493), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_465), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_471), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_465), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_457), .Y(n_514) );
BUFx10_ASAP7_75t_L g515 ( .A(n_453), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_466), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_466), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_482), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_473), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_457), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_457), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_475), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_479), .B(n_318), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_464), .B(n_410), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_461), .B(n_322), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_479), .B(n_318), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_458), .Y(n_529) );
NOR2x1p5_ASAP7_75t_L g530 ( .A(n_461), .B(n_317), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_493), .B(n_376), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_495), .B(n_471), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_530), .A2(n_469), .B1(n_470), .B2(n_480), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_506), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_506), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_530), .A2(n_480), .B1(n_453), .B2(n_452), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_512), .A2(n_452), .B1(n_490), .B2(n_477), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_510), .B(n_319), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_508), .B(n_482), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_512), .A2(n_481), .B1(n_456), .B2(n_308), .Y(n_540) );
INVx5_ASAP7_75t_L g541 ( .A(n_515), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_527), .B(n_486), .Y(n_542) );
NAND3xp33_ASAP7_75t_SL g543 ( .A(n_531), .B(n_472), .C(n_321), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_510), .B(n_319), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_515), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_505), .A2(n_308), .B1(n_363), .B2(n_321), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_505), .A2(n_363), .B1(n_386), .B2(n_383), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_498), .A2(n_383), .B1(n_386), .B2(n_487), .Y(n_548) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_499), .B(n_506), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_497), .B(n_492), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_497), .B(n_492), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_515), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_498), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_498), .A2(n_491), .B1(n_487), .B2(n_396), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_494), .Y(n_555) );
NOR2xp33_ASAP7_75t_SL g556 ( .A(n_499), .B(n_491), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_505), .A2(n_459), .B1(n_454), .B2(n_464), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_502), .B(n_460), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_505), .A2(n_459), .B1(n_454), .B2(n_475), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_496), .A2(n_459), .B1(n_454), .B2(n_475), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_498), .A2(n_396), .B1(n_358), .B2(n_460), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_507), .B(n_492), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_494), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_525), .B(n_451), .Y(n_564) );
AND2x6_ASAP7_75t_SL g565 ( .A(n_510), .B(n_293), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_499), .B(n_320), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_507), .B(n_320), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_496), .A2(n_478), .B1(n_489), .B2(n_474), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_519), .B(n_360), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_501), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_526), .B(n_360), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_528), .B(n_474), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_496), .A2(n_489), .B1(n_478), .B2(n_333), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_504), .B(n_407), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_496), .A2(n_358), .B1(n_467), .B2(n_485), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_500), .B(n_407), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_500), .B(n_409), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_501), .B(n_467), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_503), .A2(n_343), .B(n_344), .C(n_342), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_496), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_511), .B(n_433), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_511), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_513), .A2(n_352), .B1(n_401), .B2(n_334), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_513), .B(n_433), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_516), .A2(n_348), .B1(n_350), .B2(n_346), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_516), .B(n_345), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_517), .A2(n_373), .B1(n_375), .B2(n_362), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_517), .B(n_445), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_518), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_SL g592 ( .A1(n_518), .A2(n_395), .B(n_412), .C(n_311), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_520), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_523), .A2(n_381), .B1(n_398), .B2(n_379), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_523), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_524), .B(n_441), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_509), .A2(n_485), .B1(n_400), .B2(n_406), .C(n_404), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_521), .A2(n_476), .B(n_371), .C(n_330), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_514), .B(n_367), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_521), .B(n_292), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_522), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_514), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_572), .A2(n_476), .B(n_371), .C(n_330), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_567), .B(n_301), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_544), .B(n_334), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_588), .B(n_352), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_573), .B(n_314), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_546), .B(n_370), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_563), .A2(n_484), .B(n_299), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_580), .A2(n_441), .B1(n_417), .B2(n_418), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_580), .A2(n_420), .B1(n_421), .B2(n_416), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_596), .B(n_429), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_538), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_582), .A2(n_425), .B1(n_430), .B2(n_422), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_558), .A2(n_366), .B1(n_369), .B2(n_341), .Y(n_616) );
OAI22x1_ASAP7_75t_L g617 ( .A1(n_548), .A2(n_387), .B1(n_393), .B2(n_372), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_547), .Y(n_618) );
BUFx3_ASAP7_75t_L g619 ( .A(n_591), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_541), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_534), .Y(n_621) );
AO21x1_ASAP7_75t_L g622 ( .A1(n_600), .A2(n_302), .B(n_298), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_541), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_537), .B(n_437), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_535), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_568), .A2(n_571), .B(n_555), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_571), .A2(n_306), .B(n_305), .Y(n_627) );
BUFx12f_ASAP7_75t_L g628 ( .A(n_565), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_575), .A2(n_440), .B1(n_442), .B2(n_434), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_549), .A2(n_310), .B(n_307), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_550), .B(n_443), .Y(n_631) );
AO32x2_ASAP7_75t_L g632 ( .A1(n_592), .A2(n_448), .A3(n_462), .B1(n_468), .B2(n_458), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_551), .B(n_323), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_536), .A2(n_328), .B1(n_364), .B2(n_331), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_562), .B(n_328), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_575), .A2(n_380), .B1(n_438), .B2(n_331), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_539), .A2(n_329), .B(n_324), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_542), .A2(n_338), .B(n_332), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_569), .A2(n_450), .B1(n_413), .B2(n_444), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_559), .A2(n_340), .B(n_339), .Y(n_640) );
AO22x1_ASAP7_75t_L g641 ( .A1(n_556), .A2(n_436), .B1(n_446), .B2(n_439), .Y(n_641) );
INVx4_ASAP7_75t_L g642 ( .A(n_545), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_560), .A2(n_353), .B1(n_357), .B2(n_351), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_533), .B(n_336), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_593), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_593), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_561), .B(n_365), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_570), .B(n_377), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_585), .Y(n_649) );
CKINVDCx14_ASAP7_75t_R g650 ( .A(n_543), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_545), .B(n_378), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_564), .B(n_368), .Y(n_652) );
AO32x1_ASAP7_75t_L g653 ( .A1(n_595), .A2(n_389), .A3(n_390), .B1(n_388), .B2(n_384), .Y(n_653) );
INVx3_ASAP7_75t_SL g654 ( .A(n_583), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_553), .Y(n_655) );
OAI22xp5_ASAP7_75t_SL g656 ( .A1(n_554), .A2(n_391), .B1(n_397), .B2(n_392), .Y(n_656) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_576), .B(n_399), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_540), .A2(n_403), .B(n_402), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_559), .A2(n_411), .B(n_405), .Y(n_659) );
BUFx3_ASAP7_75t_L g660 ( .A(n_574), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_557), .A2(n_415), .B(n_414), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_532), .A2(n_423), .B(n_419), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_574), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_577), .A2(n_413), .B1(n_444), .B2(n_368), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_552), .A2(n_428), .B(n_426), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_586), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_557), .A2(n_432), .B(n_431), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_578), .B(n_435), .Y(n_668) );
OAI22xp5_ASAP7_75t_SL g669 ( .A1(n_587), .A2(n_312), .B1(n_374), .B2(n_354), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_587), .B(n_19), .Y(n_670) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_566), .B(n_312), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_597), .A2(n_447), .B1(n_374), .B2(n_408), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_579), .B(n_354), .Y(n_673) );
INVx3_ASAP7_75t_L g674 ( .A(n_602), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_601), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_590), .B(n_21), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_589), .B(n_21), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_589), .B(n_22), .Y(n_678) );
BUFx2_ASAP7_75t_SL g679 ( .A(n_599), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_581), .A2(n_529), .B(n_514), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_594), .B(n_313), .C(n_304), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_594), .B(n_23), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_600), .A2(n_26), .B(n_24), .C(n_25), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_572), .B(n_27), .Y(n_684) );
OAI21xp33_ASAP7_75t_L g685 ( .A1(n_572), .A2(n_337), .B(n_304), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_572), .Y(n_686) );
INVx4_ASAP7_75t_L g687 ( .A(n_541), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_572), .B(n_28), .Y(n_688) );
INVxp33_ASAP7_75t_L g689 ( .A(n_585), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_572), .B(n_29), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_575), .A2(n_359), .B1(n_462), .B2(n_458), .Y(n_691) );
AO22x1_ASAP7_75t_L g692 ( .A1(n_546), .A2(n_359), .B1(n_32), .B2(n_30), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_558), .A2(n_359), .B1(n_462), .B2(n_458), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_572), .Y(n_694) );
O2A1O1Ixp33_ASAP7_75t_L g695 ( .A1(n_572), .A2(n_33), .B(n_30), .C(n_31), .Y(n_695) );
NOR2xp33_ASAP7_75t_SL g696 ( .A(n_541), .B(n_359), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_584), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_572), .B(n_31), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_558), .A2(n_468), .B1(n_462), .B2(n_36), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_558), .A2(n_468), .B1(n_462), .B2(n_41), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_572), .B(n_35), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_575), .A2(n_468), .B1(n_41), .B2(n_35), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_572), .Y(n_703) );
INVx2_ASAP7_75t_SL g704 ( .A(n_596), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_541), .B(n_40), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_584), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_572), .B(n_40), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_572), .B(n_42), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_686), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_694), .B(n_44), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_603), .A2(n_154), .B(n_153), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_610), .A2(n_158), .B(n_157), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_620), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_664), .B(n_45), .C(n_47), .Y(n_714) );
AO31x2_ASAP7_75t_L g715 ( .A1(n_622), .A2(n_51), .A3(n_48), .B(n_50), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_703), .B(n_52), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_698), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_688), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_605), .B(n_54), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_658), .B(n_56), .Y(n_720) );
AO21x1_ASAP7_75t_L g721 ( .A1(n_702), .A2(n_164), .B(n_163), .Y(n_721) );
INVx3_ASAP7_75t_L g722 ( .A(n_687), .Y(n_722) );
NAND2x1p5_ASAP7_75t_L g723 ( .A(n_620), .B(n_56), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_670), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_684), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_690), .A2(n_57), .B(n_58), .C(n_59), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_687), .B(n_620), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g728 ( .A1(n_701), .A2(n_57), .B(n_58), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_707), .A2(n_59), .B(n_60), .C(n_61), .Y(n_729) );
NAND3x1_ASAP7_75t_L g730 ( .A(n_608), .B(n_60), .C(n_62), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_708), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_606), .B(n_63), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_618), .B(n_63), .Y(n_733) );
NOR2xp67_ASAP7_75t_L g734 ( .A(n_642), .B(n_166), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_619), .Y(n_735) );
AOI31xp67_ASAP7_75t_L g736 ( .A1(n_652), .A2(n_195), .A3(n_289), .B(n_288), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_689), .A2(n_64), .B(n_65), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_612), .B(n_64), .Y(n_738) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_650), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_646), .Y(n_740) );
AO31x2_ASAP7_75t_L g741 ( .A1(n_691), .A2(n_67), .A3(n_68), .B(n_69), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_677), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_651), .A2(n_168), .B(n_167), .Y(n_743) );
AO31x2_ASAP7_75t_L g744 ( .A1(n_691), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_649), .B(n_72), .Y(n_745) );
AOI31xp67_ASAP7_75t_L g746 ( .A1(n_693), .A2(n_204), .A3(n_287), .B(n_282), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_663), .B(n_73), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_678), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_614), .B(n_74), .Y(n_749) );
NAND2x1p5_ASAP7_75t_L g750 ( .A(n_623), .B(n_76), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_645), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g752 ( .A1(n_680), .A2(n_174), .B(n_169), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_637), .A2(n_177), .B(n_175), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_624), .B(n_76), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_647), .B(n_611), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_640), .A2(n_77), .B(n_79), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_640), .A2(n_77), .B(n_79), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_682), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_638), .A2(n_181), .B(n_180), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g760 ( .A1(n_629), .A2(n_80), .B(n_83), .C(n_84), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_L g761 ( .A1(n_629), .A2(n_83), .B(n_84), .C(n_85), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_675), .Y(n_762) );
INVx5_ASAP7_75t_L g763 ( .A(n_655), .Y(n_763) );
AO31x2_ASAP7_75t_L g764 ( .A1(n_643), .A2(n_86), .A3(n_87), .B(n_88), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_704), .B(n_86), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_683), .A2(n_90), .B(n_91), .C(n_92), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_668), .A2(n_186), .B(n_184), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_623), .B(n_90), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_609), .A2(n_222), .B(n_278), .Y(n_769) );
AO21x1_ASAP7_75t_L g770 ( .A1(n_702), .A2(n_218), .B(n_277), .Y(n_770) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_674), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_642), .B(n_92), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_633), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_621), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_616), .B(n_93), .Y(n_775) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_655), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_660), .B(n_93), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_697), .A2(n_214), .B(n_273), .Y(n_778) );
INVx2_ASAP7_75t_SL g779 ( .A(n_628), .Y(n_779) );
BUFx2_ASAP7_75t_L g780 ( .A(n_671), .Y(n_780) );
NOR2x1_ASAP7_75t_L g781 ( .A(n_681), .B(n_95), .Y(n_781) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_627), .A2(n_212), .B(n_271), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_705), .B(n_95), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_699), .B(n_96), .C(n_97), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_706), .A2(n_227), .B(n_269), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g786 ( .A1(n_634), .A2(n_695), .B(n_643), .C(n_615), .Y(n_786) );
AO31x2_ASAP7_75t_L g787 ( .A1(n_639), .A2(n_96), .A3(n_98), .B(n_100), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_635), .Y(n_788) );
A2O1A1Ixp33_ASAP7_75t_L g789 ( .A1(n_676), .A2(n_98), .B(n_100), .C(n_101), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_644), .B(n_102), .Y(n_790) );
AO31x2_ASAP7_75t_L g791 ( .A1(n_636), .A2(n_102), .A3(n_103), .B(n_104), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g792 ( .A1(n_665), .A2(n_103), .B(n_104), .C(n_105), .Y(n_792) );
BUFx4_ASAP7_75t_SL g793 ( .A(n_625), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_604), .B(n_105), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_673), .A2(n_206), .B(n_266), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_659), .A2(n_106), .B(n_107), .Y(n_796) );
OAI21xp33_ASAP7_75t_L g797 ( .A1(n_700), .A2(n_107), .B(n_108), .Y(n_797) );
INVxp67_ASAP7_75t_L g798 ( .A(n_669), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_659), .A2(n_108), .B1(n_111), .B2(n_112), .Y(n_799) );
BUFx2_ASAP7_75t_L g800 ( .A(n_671), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_630), .A2(n_228), .B(n_262), .Y(n_801) );
BUFx3_ASAP7_75t_L g802 ( .A(n_654), .Y(n_802) );
BUFx10_ASAP7_75t_L g803 ( .A(n_613), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_661), .A2(n_203), .B(n_261), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_631), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_607), .A2(n_201), .B(n_258), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_696), .A2(n_199), .B(n_256), .Y(n_807) );
BUFx3_ASAP7_75t_L g808 ( .A(n_613), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_648), .B(n_113), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_667), .A2(n_205), .B(n_253), .Y(n_810) );
AO31x2_ASAP7_75t_L g811 ( .A1(n_632), .A2(n_114), .A3(n_115), .B(n_116), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_666), .Y(n_812) );
AOI21xp5_ASAP7_75t_SL g813 ( .A1(n_667), .A2(n_192), .B(n_248), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_679), .Y(n_814) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_685), .A2(n_191), .B(n_246), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_672), .B(n_114), .Y(n_816) );
OR2x2_ASAP7_75t_L g817 ( .A(n_617), .B(n_115), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_692), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_657), .B(n_116), .Y(n_819) );
OAI22x1_ASAP7_75t_L g820 ( .A1(n_656), .A2(n_117), .B1(n_118), .B2(n_119), .Y(n_820) );
OAI21xp5_ASAP7_75t_L g821 ( .A1(n_662), .A2(n_118), .B(n_120), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_641), .B(n_121), .Y(n_822) );
AO31x2_ASAP7_75t_L g823 ( .A1(n_632), .A2(n_121), .A3(n_123), .B(n_125), .Y(n_823) );
AOI21x1_ASAP7_75t_L g824 ( .A1(n_632), .A2(n_232), .B(n_245), .Y(n_824) );
BUFx3_ASAP7_75t_L g825 ( .A(n_653), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_653), .A2(n_230), .B(n_244), .Y(n_826) );
BUFx24_ASAP7_75t_L g827 ( .A(n_653), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_686), .B(n_126), .Y(n_828) );
A2O1A1Ixp33_ASAP7_75t_L g829 ( .A1(n_684), .A2(n_127), .B(n_128), .C(n_129), .Y(n_829) );
OR2x6_ASAP7_75t_L g830 ( .A(n_687), .B(n_128), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g831 ( .A1(n_626), .A2(n_233), .B(n_243), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_686), .B(n_129), .Y(n_832) );
NOR4xp25_ASAP7_75t_L g833 ( .A(n_695), .B(n_130), .C(n_131), .D(n_132), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_626), .A2(n_190), .B(n_242), .Y(n_834) );
NAND3xp33_ASAP7_75t_L g835 ( .A(n_603), .B(n_130), .C(n_131), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_614), .Y(n_836) );
NAND2x1p5_ASAP7_75t_L g837 ( .A(n_620), .B(n_133), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_686), .B(n_135), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_793), .Y(n_839) );
OA21x2_ASAP7_75t_L g840 ( .A1(n_711), .A2(n_237), .B(n_241), .Y(n_840) );
AND2x4_ASAP7_75t_L g841 ( .A(n_805), .B(n_135), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_748), .A2(n_136), .B(n_758), .Y(n_842) );
NAND2x1p5_ASAP7_75t_L g843 ( .A(n_802), .B(n_136), .Y(n_843) );
AOI21xp33_ASAP7_75t_L g844 ( .A1(n_786), .A2(n_818), .B(n_766), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_718), .A2(n_712), .B(n_725), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_724), .B(n_742), .Y(n_846) );
OA21x2_ASAP7_75t_L g847 ( .A1(n_824), .A2(n_835), .B(n_815), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g848 ( .A1(n_835), .A2(n_788), .B(n_773), .Y(n_848) );
OA21x2_ASAP7_75t_L g849 ( .A1(n_804), .A2(n_810), .B(n_826), .Y(n_849) );
BUFx3_ASAP7_75t_L g850 ( .A(n_836), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_830), .Y(n_851) );
OAI21x1_ASAP7_75t_SL g852 ( .A1(n_756), .A2(n_796), .B(n_757), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_762), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_830), .A2(n_796), .B1(n_757), .B2(n_756), .Y(n_854) );
OA21x2_ASAP7_75t_L g855 ( .A1(n_797), .A2(n_770), .B(n_721), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_755), .B(n_808), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_774), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_751), .Y(n_858) );
BUFx2_ASAP7_75t_R g859 ( .A(n_822), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_727), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_710), .Y(n_861) );
OR2x6_ASAP7_75t_L g862 ( .A(n_779), .B(n_727), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_719), .B(n_732), .Y(n_863) );
AND2x4_ASAP7_75t_L g864 ( .A(n_727), .B(n_722), .Y(n_864) );
OAI21xp5_ASAP7_75t_L g865 ( .A1(n_784), .A2(n_747), .B(n_816), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_716), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_828), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_733), .B(n_717), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_745), .A2(n_775), .B1(n_738), .B2(n_754), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_749), .B(n_790), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_832), .Y(n_871) );
BUFx12f_ASAP7_75t_L g872 ( .A(n_803), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_794), .B(n_765), .Y(n_873) );
BUFx2_ASAP7_75t_L g874 ( .A(n_722), .Y(n_874) );
OR2x6_ASAP7_75t_L g875 ( .A(n_750), .B(n_814), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_838), .B(n_735), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_817), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_809), .B(n_777), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_812), .B(n_820), .Y(n_879) );
AO31x2_ASAP7_75t_L g880 ( .A1(n_799), .A2(n_827), .A3(n_729), .B(n_726), .Y(n_880) );
BUFx3_ASAP7_75t_L g881 ( .A(n_713), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_771), .B(n_833), .Y(n_882) );
BUFx2_ASAP7_75t_SL g883 ( .A(n_763), .Y(n_883) );
OA21x2_ASAP7_75t_L g884 ( .A1(n_782), .A2(n_801), .B(n_728), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_715), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_784), .A2(n_825), .B(n_806), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_715), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_833), .B(n_819), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_739), .A2(n_737), .B1(n_800), .B2(n_780), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_791), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_739), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_821), .B(n_760), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_791), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_821), .B(n_764), .Y(n_894) );
AND2x4_ASAP7_75t_L g895 ( .A(n_763), .B(n_776), .Y(n_895) );
OR2x6_ASAP7_75t_L g896 ( .A(n_723), .B(n_837), .Y(n_896) );
O2A1O1Ixp33_ASAP7_75t_L g897 ( .A1(n_829), .A2(n_789), .B(n_761), .C(n_792), .Y(n_897) );
INVx4_ASAP7_75t_L g898 ( .A(n_776), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_753), .A2(n_759), .B(n_714), .Y(n_899) );
OA21x2_ASAP7_75t_L g900 ( .A1(n_834), .A2(n_831), .B(n_767), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_720), .B(n_783), .Y(n_901) );
OR2x6_ASAP7_75t_L g902 ( .A(n_730), .B(n_813), .Y(n_902) );
OAI222xp33_ASAP7_75t_L g903 ( .A1(n_772), .A2(n_768), .B1(n_781), .B2(n_807), .C1(n_743), .C2(n_795), .Y(n_903) );
OA21x2_ASAP7_75t_L g904 ( .A1(n_769), .A2(n_778), .B(n_785), .Y(n_904) );
OA21x2_ASAP7_75t_L g905 ( .A1(n_734), .A2(n_746), .B(n_736), .Y(n_905) );
AOI21xp5_ASAP7_75t_SL g906 ( .A1(n_741), .A2(n_744), .B(n_764), .Y(n_906) );
AND2x4_ASAP7_75t_L g907 ( .A(n_787), .B(n_744), .Y(n_907) );
AND2x4_ASAP7_75t_SL g908 ( .A(n_811), .B(n_823), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_793), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_724), .B(n_742), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_L g911 ( .A1(n_786), .A2(n_766), .B(n_731), .C(n_725), .Y(n_911) );
OAI21xp5_ASAP7_75t_L g912 ( .A1(n_748), .A2(n_603), .B(n_758), .Y(n_912) );
AO31x2_ASAP7_75t_L g913 ( .A1(n_721), .A2(n_603), .A3(n_598), .B(n_770), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_836), .B(n_546), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_711), .A2(n_603), .B(n_752), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_802), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g917 ( .A1(n_786), .A2(n_766), .B(n_731), .C(n_725), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_724), .B(n_742), .Y(n_918) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_740), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_793), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_836), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_798), .B(n_689), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_802), .Y(n_923) );
INVx2_ASAP7_75t_SL g924 ( .A(n_793), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_798), .A2(n_689), .B1(n_618), .B2(n_649), .Y(n_925) );
INVx1_ASAP7_75t_SL g926 ( .A(n_836), .Y(n_926) );
AND2x6_ASAP7_75t_L g927 ( .A(n_740), .B(n_646), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_709), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_724), .B(n_742), .Y(n_929) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_748), .A2(n_603), .B(n_758), .Y(n_930) );
AND2x4_ASAP7_75t_L g931 ( .A(n_805), .B(n_686), .Y(n_931) );
BUFx8_ASAP7_75t_L g932 ( .A(n_779), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_709), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_798), .B(n_572), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_709), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g936 ( .A1(n_786), .A2(n_766), .B(n_731), .C(n_725), .Y(n_936) );
BUFx2_ASAP7_75t_L g937 ( .A(n_836), .Y(n_937) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_740), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_724), .B(n_742), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_836), .B(n_546), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_724), .B(n_742), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_709), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_724), .B(n_742), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_931), .Y(n_944) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_919), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_928), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_882), .B(n_888), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_921), .Y(n_948) );
HB1xp67_ASAP7_75t_SL g949 ( .A(n_932), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_934), .B(n_925), .Y(n_950) );
OR2x2_ASAP7_75t_L g951 ( .A(n_888), .B(n_846), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_846), .B(n_910), .Y(n_952) );
OR2x6_ASAP7_75t_L g953 ( .A(n_875), .B(n_854), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_937), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_885), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_910), .B(n_918), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_858), .B(n_853), .Y(n_957) );
AND2x4_ASAP7_75t_L g958 ( .A(n_864), .B(n_895), .Y(n_958) );
HB1xp67_ASAP7_75t_L g959 ( .A(n_926), .Y(n_959) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_926), .Y(n_960) );
OR2x6_ASAP7_75t_L g961 ( .A(n_875), .B(n_854), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_887), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_922), .B(n_914), .Y(n_963) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_850), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_857), .B(n_911), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_889), .A2(n_891), .B1(n_877), .B2(n_841), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_841), .A2(n_869), .B1(n_856), .B2(n_851), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_917), .B(n_936), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_890), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_933), .B(n_935), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_893), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_942), .B(n_894), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_929), .Y(n_973) );
OR2x2_ASAP7_75t_L g974 ( .A(n_929), .B(n_939), .Y(n_974) );
INVxp67_ASAP7_75t_SL g975 ( .A(n_938), .Y(n_975) );
INVxp67_ASAP7_75t_SL g976 ( .A(n_863), .Y(n_976) );
INVx3_ASAP7_75t_L g977 ( .A(n_898), .Y(n_977) );
NOR2x1_ASAP7_75t_L g978 ( .A(n_883), .B(n_875), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_941), .Y(n_979) );
BUFx3_ASAP7_75t_L g980 ( .A(n_923), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_842), .B(n_861), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_943), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_943), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_842), .B(n_866), .Y(n_984) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_881), .Y(n_985) );
OR2x6_ASAP7_75t_L g986 ( .A(n_896), .B(n_902), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_867), .B(n_871), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_907), .B(n_912), .Y(n_988) );
OR2x6_ASAP7_75t_L g989 ( .A(n_896), .B(n_902), .Y(n_989) );
BUFx3_ASAP7_75t_L g990 ( .A(n_872), .Y(n_990) );
OR2x6_ASAP7_75t_L g991 ( .A(n_896), .B(n_902), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_907), .Y(n_992) );
OR2x6_ASAP7_75t_L g993 ( .A(n_862), .B(n_860), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_912), .B(n_930), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_930), .Y(n_995) );
OR2x2_ASAP7_75t_L g996 ( .A(n_868), .B(n_940), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_844), .B(n_874), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_908), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_870), .B(n_876), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_906), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_927), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_844), .B(n_848), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_927), .Y(n_1003) );
AO21x2_ASAP7_75t_L g1004 ( .A1(n_886), .A2(n_852), .B(n_899), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_848), .B(n_892), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1006 ( .A(n_876), .B(n_892), .Y(n_1006) );
OR2x2_ASAP7_75t_L g1007 ( .A(n_878), .B(n_873), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_879), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_878), .B(n_869), .Y(n_1009) );
INVx5_ASAP7_75t_L g1010 ( .A(n_898), .Y(n_1010) );
OAI222xp33_ASAP7_75t_L g1011 ( .A1(n_843), .A2(n_924), .B1(n_839), .B2(n_920), .C1(n_909), .C2(n_897), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_865), .B(n_845), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_865), .B(n_880), .Y(n_1013) );
INVxp67_ASAP7_75t_SL g1014 ( .A(n_901), .Y(n_1014) );
INVx2_ASAP7_75t_L g1015 ( .A(n_905), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_880), .B(n_901), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_859), .Y(n_1017) );
INVx3_ASAP7_75t_L g1018 ( .A(n_880), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_972), .B(n_855), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_972), .B(n_855), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_988), .B(n_913), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_969), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_969), .Y(n_1023) );
AND2x4_ASAP7_75t_SL g1024 ( .A(n_986), .B(n_916), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_988), .B(n_913), .Y(n_1025) );
INVx1_ASAP7_75t_SL g1026 ( .A(n_949), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_971), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_971), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_1010), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1016), .B(n_884), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_959), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_960), .Y(n_1032) );
INVx3_ASAP7_75t_L g1033 ( .A(n_1010), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1016), .B(n_884), .Y(n_1034) );
INVx5_ASAP7_75t_SL g1035 ( .A(n_986), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_952), .B(n_932), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1013), .B(n_847), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1013), .B(n_847), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1005), .B(n_915), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1005), .B(n_849), .Y(n_1040) );
INVx5_ASAP7_75t_SL g1041 ( .A(n_986), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_947), .B(n_840), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_992), .B(n_900), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_955), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_992), .B(n_900), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_945), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_947), .B(n_904), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1002), .B(n_904), .Y(n_1048) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_980), .Y(n_1049) );
NAND2x1_ASAP7_75t_L g1050 ( .A(n_953), .B(n_903), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1002), .B(n_994), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_956), .B(n_974), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_994), .B(n_970), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_962), .B(n_953), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_951), .B(n_1009), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_961), .B(n_968), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_951), .B(n_1009), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_976), .B(n_956), .Y(n_1058) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_964), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_961), .B(n_968), .Y(n_1060) );
INVx3_ASAP7_75t_L g1061 ( .A(n_1010), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_973), .B(n_979), .Y(n_1062) );
INVxp67_ASAP7_75t_L g1063 ( .A(n_948), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_961), .B(n_957), .Y(n_1064) );
INVxp67_ASAP7_75t_L g1065 ( .A(n_954), .Y(n_1065) );
NAND2xp5_ASAP7_75t_SL g1066 ( .A(n_1010), .B(n_978), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1015), .Y(n_1067) );
INVx4_ASAP7_75t_L g1068 ( .A(n_986), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_961), .B(n_957), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1014), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1071 ( .A(n_975), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_998), .B(n_989), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1022), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1051), .B(n_1018), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1051), .B(n_1004), .Y(n_1075) );
INVx2_ASAP7_75t_L g1076 ( .A(n_1067), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1053), .B(n_987), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1053), .B(n_1004), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1021), .B(n_1000), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1025), .B(n_1012), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g1081 ( .A(n_1046), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1071), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1039), .B(n_1012), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1039), .B(n_998), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_1031), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1019), .B(n_1008), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1023), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1019), .B(n_965), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1032), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_1055), .B(n_1006), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1027), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1028), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1055), .B(n_999), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1020), .B(n_965), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1057), .B(n_999), .Y(n_1095) );
AOI21xp5_ASAP7_75t_L g1096 ( .A1(n_1050), .A2(n_989), .B(n_991), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1057), .B(n_996), .Y(n_1097) );
CKINVDCx16_ASAP7_75t_R g1098 ( .A(n_1026), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1020), .B(n_997), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1100 ( .A(n_1054), .B(n_1001), .Y(n_1100) );
NAND3xp33_ASAP7_75t_L g1101 ( .A(n_1063), .B(n_963), .C(n_966), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_1059), .Y(n_1102) );
AND2x4_ASAP7_75t_L g1103 ( .A(n_1068), .B(n_1003), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1040), .B(n_997), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1040), .B(n_981), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_1058), .B(n_996), .Y(n_1106) );
NAND2x1_ASAP7_75t_SL g1107 ( .A(n_1033), .B(n_977), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1048), .B(n_981), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1048), .B(n_984), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1064), .B(n_984), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1049), .Y(n_1111) );
INVx1_ASAP7_75t_SL g1112 ( .A(n_1049), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1064), .B(n_995), .Y(n_1113) );
NOR2xp67_ASAP7_75t_L g1114 ( .A(n_1033), .B(n_1017), .Y(n_1114) );
INVxp67_ASAP7_75t_L g1115 ( .A(n_1036), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1069), .B(n_995), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1073), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1083), .B(n_1047), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1076), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1099), .B(n_1037), .Y(n_1120) );
AND2x2_ASAP7_75t_SL g1121 ( .A(n_1111), .B(n_1068), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1076), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1080), .B(n_1065), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1099), .B(n_1037), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1104), .B(n_1038), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1083), .B(n_1047), .Y(n_1126) );
OR2x6_ASAP7_75t_L g1127 ( .A(n_1096), .B(n_1068), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1104), .B(n_1078), .Y(n_1128) );
INVxp67_ASAP7_75t_L g1129 ( .A(n_1081), .Y(n_1129) );
INVx2_ASAP7_75t_SL g1130 ( .A(n_1107), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1075), .B(n_1030), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1087), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1075), .B(n_1030), .Y(n_1133) );
NOR2x1_ASAP7_75t_L g1134 ( .A(n_1112), .B(n_1066), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1080), .B(n_1052), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1108), .B(n_1034), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1108), .B(n_1034), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1086), .B(n_1070), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1109), .B(n_1043), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1109), .B(n_1042), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1088), .B(n_1043), .Y(n_1141) );
NAND2xp67_ASAP7_75t_L g1142 ( .A(n_1084), .B(n_1024), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1082), .Y(n_1143) );
NAND2xp67_ASAP7_75t_L g1144 ( .A(n_1084), .B(n_1024), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1088), .B(n_1045), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1077), .B(n_1044), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1094), .B(n_1045), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1091), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1092), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1092), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1128), .B(n_1074), .Y(n_1151) );
OAI222xp33_ASAP7_75t_L g1152 ( .A1(n_1127), .A2(n_1095), .B1(n_1093), .B2(n_1106), .C1(n_1097), .C2(n_1098), .Y(n_1152) );
INVx2_ASAP7_75t_SL g1153 ( .A(n_1121), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1128), .B(n_1074), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_1129), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1117), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1118), .B(n_1085), .Y(n_1157) );
INVx1_ASAP7_75t_SL g1158 ( .A(n_1123), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1118), .B(n_1089), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1135), .B(n_1115), .Y(n_1160) );
NAND2xp5_ASAP7_75t_SL g1161 ( .A(n_1121), .B(n_1114), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1136), .B(n_1105), .Y(n_1162) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1119), .Y(n_1163) );
INVxp33_ASAP7_75t_L g1164 ( .A(n_1138), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1126), .Y(n_1165) );
INVxp67_ASAP7_75t_L g1166 ( .A(n_1143), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1126), .B(n_1090), .Y(n_1167) );
NAND2xp33_ASAP7_75t_L g1168 ( .A(n_1134), .B(n_1029), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1140), .B(n_1090), .Y(n_1169) );
BUFx3_ASAP7_75t_L g1170 ( .A(n_1130), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1139), .B(n_1102), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1122), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1165), .B(n_1136), .Y(n_1173) );
AOI22xp33_ASAP7_75t_SL g1174 ( .A1(n_1153), .A2(n_1035), .B1(n_1041), .B2(n_1101), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1167), .B(n_1137), .Y(n_1175) );
OAI21xp33_ASAP7_75t_SL g1176 ( .A1(n_1161), .A2(n_1107), .B(n_1137), .Y(n_1176) );
AOI32xp33_ASAP7_75t_L g1177 ( .A1(n_1168), .A2(n_1125), .A3(n_1120), .B1(n_1124), .B2(n_1147), .Y(n_1177) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1163), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1169), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1162), .B(n_1120), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_1158), .A2(n_1060), .B1(n_1056), .B2(n_1079), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1157), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1162), .B(n_1141), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1159), .Y(n_1184) );
INVxp67_ASAP7_75t_L g1185 ( .A(n_1155), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1156), .Y(n_1186) );
OAI221xp5_ASAP7_75t_SL g1187 ( .A1(n_1177), .A2(n_1171), .B1(n_967), .B2(n_1095), .C(n_1170), .Y(n_1187) );
AOI221xp5_ASAP7_75t_L g1188 ( .A1(n_1185), .A2(n_1152), .B1(n_1160), .B2(n_1164), .C(n_1166), .Y(n_1188) );
OAI21xp5_ASAP7_75t_L g1189 ( .A1(n_1176), .A2(n_1168), .B(n_1011), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_1185), .A2(n_1154), .B1(n_1151), .B2(n_1146), .Y(n_1190) );
A2O1A1Ixp33_ASAP7_75t_R g1191 ( .A1(n_1173), .A2(n_1180), .B(n_1175), .C(n_1142), .Y(n_1191) );
INVxp67_ASAP7_75t_L g1192 ( .A(n_1186), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_1181), .A2(n_1100), .B1(n_1131), .B2(n_1133), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1179), .Y(n_1194) );
OAI21xp33_ASAP7_75t_SL g1195 ( .A1(n_1183), .A2(n_1147), .B(n_1145), .Y(n_1195) );
AOI322xp5_ASAP7_75t_L g1196 ( .A1(n_1182), .A2(n_1145), .A3(n_1133), .B1(n_1131), .B2(n_1110), .C1(n_1116), .C2(n_1113), .Y(n_1196) );
O2A1O1Ixp5_ASAP7_75t_L g1197 ( .A1(n_1184), .A2(n_1061), .B(n_1172), .C(n_1149), .Y(n_1197) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_1178), .A2(n_1132), .B1(n_1150), .B2(n_1149), .C(n_1148), .Y(n_1198) );
NAND4xp25_ASAP7_75t_L g1199 ( .A(n_1174), .B(n_990), .C(n_950), .D(n_1072), .Y(n_1199) );
NAND4xp25_ASAP7_75t_L g1200 ( .A(n_1189), .B(n_1187), .C(n_1188), .D(n_1199), .Y(n_1200) );
A2O1A1Ixp33_ASAP7_75t_L g1201 ( .A1(n_1195), .A2(n_1197), .B(n_1191), .C(n_1196), .Y(n_1201) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1193), .A2(n_1190), .B(n_1192), .C(n_1194), .Y(n_1202) );
NOR4xp25_ASAP7_75t_L g1203 ( .A(n_1200), .B(n_1007), .C(n_1198), .D(n_946), .Y(n_1203) );
NAND3xp33_ASAP7_75t_SL g1204 ( .A(n_1203), .B(n_1201), .C(n_1202), .Y(n_1204) );
INVxp67_ASAP7_75t_L g1205 ( .A(n_1204), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1205), .Y(n_1206) );
AO221x2_ASAP7_75t_L g1207 ( .A1(n_1206), .A2(n_1144), .B1(n_983), .B2(n_982), .C(n_1062), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1207), .A2(n_1061), .B1(n_1103), .B2(n_944), .Y(n_1208) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1208), .B(n_985), .C(n_993), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1209), .B(n_993), .Y(n_1210) );
AOI21xp33_ASAP7_75t_L g1211 ( .A1(n_1210), .A2(n_985), .B(n_958), .Y(n_1211) );
endmodule