module fake_jpeg_2381_n_404 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_404);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_404;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_56),
.Y(n_116)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_57),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_12),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_59),
.B(n_64),
.Y(n_120)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_66),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_65),
.B(n_96),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_10),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_70),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_10),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_74),
.B(n_75),
.Y(n_159)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_77),
.B(n_82),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_80),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_84),
.B(n_88),
.Y(n_164)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_89),
.B(n_90),
.Y(n_173)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_91),
.B(n_99),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_11),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_39),
.B(n_9),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_104),
.B(n_105),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_25),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_110),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_109),
.B1(n_46),
.B2(n_50),
.Y(n_114)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_8),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_25),
.B1(n_50),
.B2(n_46),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_115),
.A2(n_121),
.B1(n_122),
.B2(n_142),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_49),
.B(n_35),
.C(n_30),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_117),
.A2(n_137),
.B(n_123),
.C(n_153),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_52),
.B1(n_36),
.B2(n_42),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_118),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_28),
.B1(n_43),
.B2(n_35),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_27),
.B1(n_43),
.B2(n_30),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_50),
.B1(n_52),
.B2(n_26),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_128),
.A2(n_130),
.B1(n_150),
.B2(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_50),
.B1(n_52),
.B2(n_26),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_54),
.B(n_42),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_117),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_63),
.A2(n_21),
.B1(n_41),
.B2(n_36),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_60),
.A2(n_21),
.B1(n_41),
.B2(n_39),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_55),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_161),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_140),
.A2(n_152),
.B1(n_162),
.B2(n_165),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_47),
.B1(n_1),
.B2(n_3),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_146),
.A2(n_155),
.B1(n_112),
.B2(n_154),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_47),
.B1(n_4),
.B2(n_5),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_69),
.A2(n_0),
.B1(n_6),
.B2(n_80),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_86),
.A2(n_6),
.B1(n_106),
.B2(n_92),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_109),
.B1(n_81),
.B2(n_93),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_76),
.A2(n_81),
.B1(n_93),
.B2(n_95),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_76),
.A2(n_44),
.B1(n_97),
.B2(n_103),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_166),
.A2(n_168),
.B1(n_175),
.B2(n_153),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_95),
.A2(n_84),
.B1(n_77),
.B2(n_105),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_170),
.B1(n_174),
.B2(n_176),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_97),
.A2(n_44),
.B1(n_103),
.B2(n_52),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_84),
.B1(n_88),
.B2(n_105),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_97),
.A2(n_44),
.B1(n_103),
.B2(n_52),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_174),
.B1(n_127),
.B2(n_141),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_182),
.A2(n_193),
.B1(n_200),
.B2(n_180),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_223),
.Y(n_251)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_120),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_186),
.B(n_190),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_187),
.B(n_188),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_189),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_116),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_133),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_224),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_158),
.CI(n_160),
.CON(n_192),
.SN(n_192)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_192),
.B(n_196),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_123),
.A2(n_141),
.B1(n_130),
.B2(n_128),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_177),
.C(n_131),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_206),
.C(n_183),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_113),
.Y(n_197)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_151),
.B1(n_167),
.B2(n_113),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

OR2x4_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_131),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_233),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_137),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_132),
.B(n_147),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_217),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_163),
.B(n_143),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_210),
.B(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_119),
.B(n_124),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_212),
.C(n_232),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_119),
.B(n_124),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_213),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_143),
.B(n_144),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_144),
.B(n_111),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_219),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_111),
.B(n_145),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_156),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_126),
.A2(n_156),
.B1(n_148),
.B2(n_149),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_148),
.A2(n_112),
.B1(n_149),
.B2(n_139),
.Y(n_229)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_127),
.B(n_139),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_237),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_159),
.Y(n_232)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_117),
.A2(n_175),
.B(n_168),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_225),
.B(n_202),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_113),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_258),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_187),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_191),
.B(n_183),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_207),
.A2(n_204),
.B1(n_197),
.B2(n_237),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_209),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_244),
.B1(n_267),
.B2(n_263),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_181),
.B1(n_229),
.B2(n_213),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_226),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_180),
.A2(n_200),
.B1(n_234),
.B2(n_220),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_227),
.B1(n_223),
.B2(n_184),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_192),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_192),
.B(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_198),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_276),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_253),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_284),
.B1(n_287),
.B2(n_294),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_214),
.B1(n_201),
.B2(n_222),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_283),
.A2(n_286),
.B1(n_251),
.B2(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_285),
.B(n_291),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_199),
.B1(n_205),
.B2(n_230),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_219),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_246),
.B(n_238),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_289),
.B(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_215),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_203),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_215),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_295),
.Y(n_325)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_215),
.B1(n_233),
.B2(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_247),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_240),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_297),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_240),
.B(n_256),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_254),
.B(n_255),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_249),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_243),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_248),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_301),
.A2(n_245),
.B(n_243),
.Y(n_323)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_281),
.A2(n_251),
.B(n_250),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_311),
.A2(n_312),
.B(n_282),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_250),
.B(n_266),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_255),
.B1(n_239),
.B2(n_251),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_239),
.B1(n_272),
.B2(n_252),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_288),
.B1(n_283),
.B2(n_292),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_325),
.Y(n_340)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_286),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_329),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_273),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_314),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_289),
.Y(n_330)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_330),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_331),
.A2(n_343),
.B(n_311),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_298),
.C(n_295),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_320),
.C(n_306),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_276),
.Y(n_333)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_294),
.B1(n_316),
.B2(n_315),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_319),
.B(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_325),
.B(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_341),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_279),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_313),
.B1(n_304),
.B2(n_312),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_344),
.A2(n_338),
.B1(n_343),
.B2(n_330),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_308),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_352),
.C(n_355),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_323),
.B(n_279),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_327),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_333),
.C(n_342),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_277),
.C(n_318),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_277),
.C(n_285),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_338),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_349),
.B(n_326),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_364),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_361),
.Y(n_376)
);

OAI21x1_ASAP7_75t_SL g371 ( 
.A1(n_362),
.A2(n_357),
.B(n_350),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_351),
.C(n_349),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_365),
.A2(n_368),
.B1(n_358),
.B2(n_344),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_366),
.Y(n_375)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_367),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_301),
.C(n_296),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_346),
.C(n_354),
.Y(n_373)
);

AOI21xp33_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_336),
.B(n_348),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_363),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_373),
.B(n_376),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_352),
.C(n_345),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_339),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_381),
.B(n_355),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_384),
.A2(n_363),
.B1(n_329),
.B2(n_371),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_366),
.B1(n_368),
.B2(n_338),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_378),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_389),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_376),
.C(n_377),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_388),
.A2(n_392),
.B(n_384),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_382),
.A2(n_372),
.B1(n_362),
.B2(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_390),
.B(n_391),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_395),
.C(n_388),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_387),
.A2(n_386),
.B(n_356),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_SL g397 ( 
.A1(n_396),
.A2(n_392),
.B(n_348),
.C(n_356),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_398),
.Y(n_401)
);

AOI322xp5_ASAP7_75t_L g398 ( 
.A1(n_394),
.A2(n_337),
.A3(n_335),
.B1(n_328),
.B2(n_307),
.C1(n_309),
.C2(n_321),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_399),
.B(n_314),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_328),
.C(n_337),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_401),
.B(n_335),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_322),
.Y(n_404)
);


endmodule