module real_aes_9110_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_653;
wire n_365;
wire n_637;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_0), .A2(n_190), .B1(n_481), .B2(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_1), .A2(n_197), .B1(n_470), .B2(n_506), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_2), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_3), .B(n_298), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_4), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_5), .B(n_296), .Y(n_623) );
AOI22xp5_ASAP7_75t_SL g513 ( .A1(n_6), .A2(n_50), .B1(n_448), .B2(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_7), .B(n_298), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_8), .A2(n_59), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_9), .A2(n_101), .B1(n_451), .B2(n_452), .Y(n_450) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_10), .B(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_11), .A2(n_147), .B1(n_393), .B2(n_530), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_12), .A2(n_96), .B1(n_347), .B2(n_426), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_13), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_14), .A2(n_114), .B1(n_499), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_15), .A2(n_109), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_16), .A2(n_86), .B1(n_105), .B2(n_376), .C1(n_586), .C2(n_619), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_17), .A2(n_154), .B1(n_407), .B2(n_628), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_18), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_19), .A2(n_28), .B1(n_290), .B2(n_416), .Y(n_475) );
INVx1_ASAP7_75t_L g309 ( .A(n_20), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_21), .A2(n_520), .B1(n_557), .B2(n_558), .Y(n_519) );
INVx1_ASAP7_75t_L g558 ( .A(n_21), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_22), .A2(n_142), .B1(n_442), .B2(n_443), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_23), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_24), .Y(n_334) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_25), .A2(n_69), .B1(n_231), .B2(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g648 ( .A(n_25), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_26), .Y(n_394) );
AOI22xp5_ASAP7_75t_SL g512 ( .A1(n_27), .A2(n_202), .B1(n_351), .B2(n_481), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_29), .A2(n_52), .B1(n_605), .B2(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_30), .B(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_31), .A2(n_32), .B1(n_290), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_33), .A2(n_65), .B1(n_439), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_34), .A2(n_130), .B1(n_271), .B2(n_630), .Y(n_662) );
AOI22xp5_ASAP7_75t_SL g508 ( .A1(n_35), .A2(n_113), .B1(n_345), .B2(n_480), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_36), .A2(n_47), .B1(n_375), .B2(n_376), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_37), .A2(n_200), .B1(n_304), .B2(n_422), .Y(n_421) );
AO22x2_ASAP7_75t_L g235 ( .A1(n_38), .A2(n_72), .B1(n_231), .B2(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g649 ( .A(n_38), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_39), .A2(n_54), .B1(n_302), .B2(n_416), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_40), .A2(n_128), .B1(n_168), .B2(n_289), .C1(n_332), .C2(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_41), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_42), .A2(n_132), .B1(n_389), .B2(n_410), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_43), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_44), .A2(n_206), .B1(n_353), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_45), .A2(n_66), .B1(n_595), .B2(n_596), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_46), .Y(n_379) );
INVxp67_ASAP7_75t_L g672 ( .A(n_48), .Y(n_672) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_48), .B(n_654), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_49), .A2(n_581), .B1(n_582), .B2(n_608), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_49), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_51), .A2(n_183), .B1(n_355), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_53), .A2(n_103), .B1(n_343), .B2(n_345), .Y(n_342) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_55), .A2(n_92), .B1(n_347), .B2(n_348), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_56), .A2(n_119), .B1(n_470), .B2(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g576 ( .A(n_57), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_58), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_60), .A2(n_191), .B1(n_306), .B2(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_61), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_62), .A2(n_129), .B1(n_408), .B2(n_436), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_63), .A2(n_194), .B1(n_291), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_64), .A2(n_70), .B1(n_419), .B2(n_573), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_67), .A2(n_165), .B1(n_307), .B2(n_506), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_68), .A2(n_102), .B1(n_226), .B2(n_353), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_71), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_73), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_74), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g214 ( .A(n_75), .B(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_76), .A2(n_126), .B1(n_351), .B2(n_447), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_77), .A2(n_90), .B1(n_437), .B2(n_530), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_78), .A2(n_111), .B1(n_284), .B2(n_290), .Y(n_330) );
INVx1_ASAP7_75t_L g211 ( .A(n_79), .Y(n_211) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_80), .A2(n_208), .B(n_216), .C(n_650), .Y(n_207) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_81), .A2(n_88), .B1(n_226), .B2(n_348), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_82), .Y(n_370) );
OA22x2_ASAP7_75t_L g316 ( .A1(n_83), .A2(n_317), .B1(n_318), .B2(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_83), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_84), .A2(n_115), .B1(n_428), .B2(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_85), .A2(n_87), .B1(n_536), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_89), .A2(n_104), .B1(n_304), .B2(n_578), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_91), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_93), .A2(n_167), .B1(n_343), .B2(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_94), .A2(n_100), .B1(n_434), .B2(n_437), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_95), .A2(n_138), .B1(n_290), .B2(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_97), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_98), .A2(n_652), .B1(n_653), .B2(n_664), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_98), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_99), .Y(n_269) );
XNOR2x2_ASAP7_75t_L g430 ( .A(n_106), .B(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_107), .A2(n_127), .B1(n_448), .B2(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_108), .Y(n_273) );
INVx2_ASAP7_75t_L g215 ( .A(n_110), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_112), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_116), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_117), .A2(n_169), .B1(n_226), .B2(n_241), .Y(n_225) );
OA22x2_ASAP7_75t_L g461 ( .A1(n_118), .A2(n_462), .B1(n_463), .B2(n_486), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_118), .Y(n_462) );
INVx1_ASAP7_75t_L g634 ( .A(n_120), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_121), .B(n_332), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_122), .A2(n_201), .B1(n_388), .B2(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_123), .B(n_419), .Y(n_418) );
AND2x6_ASAP7_75t_L g210 ( .A(n_124), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_124), .Y(n_642) );
AO22x2_ASAP7_75t_L g240 ( .A1(n_125), .A2(n_179), .B1(n_231), .B2(n_236), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_131), .A2(n_192), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI22xp5_ASAP7_75t_SL g509 ( .A1(n_133), .A2(n_177), .B1(n_348), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_134), .A2(n_182), .B1(n_351), .B2(n_353), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_135), .A2(n_189), .B1(n_302), .B2(n_306), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_136), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_137), .B(n_504), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_139), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_140), .A2(n_186), .B1(n_246), .B2(n_254), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_141), .B(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_143), .A2(n_149), .B1(n_355), .B2(n_357), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_144), .A2(n_205), .B1(n_419), .B2(n_573), .Y(n_572) );
AO22x2_ASAP7_75t_L g238 ( .A1(n_145), .A2(n_184), .B1(n_231), .B2(n_232), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_146), .A2(n_204), .B1(n_271), .B2(n_428), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_148), .Y(n_322) );
AOI22xp33_ASAP7_75t_SL g283 ( .A1(n_150), .A2(n_163), .B1(n_284), .B2(n_289), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_151), .A2(n_193), .B1(n_348), .B2(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_152), .B(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_153), .A2(n_175), .B1(n_271), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_155), .A2(n_170), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_156), .A2(n_171), .B1(n_447), .B2(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g515 ( .A(n_157), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_158), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_159), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_160), .A2(n_203), .B1(n_425), .B2(n_426), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_161), .A2(n_162), .B1(n_355), .B2(n_448), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_164), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_166), .B(n_296), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_172), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_173), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_174), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_176), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_178), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_179), .B(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_180), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_181), .Y(n_543) );
INVx1_ASAP7_75t_L g645 ( .A(n_184), .Y(n_645) );
OA22x2_ASAP7_75t_L g359 ( .A1(n_185), .A2(n_360), .B1(n_361), .B2(n_362), .Y(n_359) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_185), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_187), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_188), .Y(n_391) );
INVx1_ASAP7_75t_L g231 ( .A(n_195), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_195), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_196), .A2(n_199), .B1(n_357), .B2(n_428), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_198), .B(n_467), .Y(n_502) );
INVx1_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_211), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_212), .A2(n_640), .B(n_671), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_489), .B1(n_635), .B2(n_636), .C(n_637), .Y(n_216) );
INVx1_ASAP7_75t_L g635 ( .A(n_217), .Y(n_635) );
AOI22xp5_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_460), .B1(n_487), .B2(n_488), .Y(n_217) );
INVx1_ASAP7_75t_L g487 ( .A(n_218), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B1(n_310), .B2(n_459), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
XOR2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_309), .Y(n_221) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_223), .B(n_277), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_257), .C(n_268), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_245), .Y(n_224) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx3_ASAP7_75t_L g345 ( .A(n_227), .Y(n_345) );
BUFx3_ASAP7_75t_L g410 ( .A(n_227), .Y(n_410) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_227), .Y(n_436) );
INVx2_ASAP7_75t_L g532 ( .A(n_227), .Y(n_532) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_237), .Y(n_227) );
AND2x4_ASAP7_75t_L g242 ( .A(n_228), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g272 ( .A(n_228), .B(n_263), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_228), .B(n_251), .Y(n_276) );
AND2x2_ASAP7_75t_L g352 ( .A(n_228), .B(n_251), .Y(n_352) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
AND2x2_ASAP7_75t_L g253 ( .A(n_229), .B(n_235), .Y(n_253) );
OR2x2_ASAP7_75t_L g262 ( .A(n_229), .B(n_235), .Y(n_262) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g281 ( .A(n_230), .B(n_235), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_230), .B(n_240), .Y(n_288) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g236 ( .A(n_233), .Y(n_236) );
AND2x2_ASAP7_75t_L g286 ( .A(n_234), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g336 ( .A(n_234), .Y(n_336) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g256 ( .A(n_235), .Y(n_256) );
AND2x6_ASAP7_75t_L g296 ( .A(n_237), .B(n_253), .Y(n_296) );
AND2x4_ASAP7_75t_L g300 ( .A(n_237), .B(n_261), .Y(n_300) );
INVx1_ASAP7_75t_L g325 ( .A(n_237), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_237), .B(n_253), .Y(n_328) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_238), .B(n_240), .Y(n_244) );
INVx1_ASAP7_75t_L g252 ( .A(n_238), .Y(n_252) );
INVx1_ASAP7_75t_L g264 ( .A(n_238), .Y(n_264) );
INVx1_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
AND2x2_ASAP7_75t_L g263 ( .A(n_239), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g251 ( .A(n_240), .B(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
BUFx3_ASAP7_75t_L g353 ( .A(n_242), .Y(n_353) );
INVx1_ASAP7_75t_L g399 ( .A(n_242), .Y(n_399) );
BUFx3_ASAP7_75t_L g437 ( .A(n_242), .Y(n_437) );
BUFx2_ASAP7_75t_L g481 ( .A(n_242), .Y(n_481) );
BUFx3_ASAP7_75t_L g628 ( .A(n_242), .Y(n_628) );
AND2x2_ASAP7_75t_L g408 ( .A(n_243), .B(n_336), .Y(n_408) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x6_ASAP7_75t_L g255 ( .A(n_244), .B(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_248), .Y(n_388) );
BUFx2_ASAP7_75t_L g510 ( .A(n_248), .Y(n_510) );
INVx4_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx5_ASAP7_75t_L g347 ( .A(n_249), .Y(n_347) );
INVx3_ASAP7_75t_L g428 ( .A(n_249), .Y(n_428) );
INVx1_ASAP7_75t_L g484 ( .A(n_249), .Y(n_484) );
BUFx3_ASAP7_75t_L g537 ( .A(n_249), .Y(n_537) );
INVx2_ASAP7_75t_L g566 ( .A(n_249), .Y(n_566) );
INVx8_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g308 ( .A(n_252), .Y(n_308) );
AND2x4_ASAP7_75t_L g267 ( .A(n_253), .B(n_263), .Y(n_267) );
BUFx2_ASAP7_75t_L g348 ( .A(n_254), .Y(n_348) );
BUFx2_ASAP7_75t_L g389 ( .A(n_254), .Y(n_389) );
INVx6_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g439 ( .A(n_255), .Y(n_439) );
INVx1_ASAP7_75t_SL g602 ( .A(n_255), .Y(n_602) );
INVx1_ASAP7_75t_L g305 ( .A(n_256), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B1(n_265), .B2(n_266), .Y(n_257) );
INVx2_ASAP7_75t_L g386 ( .A(n_259), .Y(n_386) );
INVx2_ASAP7_75t_SL g425 ( .A(n_259), .Y(n_425) );
INVx4_ASAP7_75t_L g447 ( .A(n_259), .Y(n_447) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_259), .Y(n_523) );
INVx5_ASAP7_75t_SL g630 ( .A(n_259), .Y(n_630) );
INVx11_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx11_ASAP7_75t_L g356 ( .A(n_260), .Y(n_356) );
AND2x6_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g324 ( .A(n_262), .B(n_325), .Y(n_324) );
AND2x6_ASAP7_75t_L g280 ( .A(n_263), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g393 ( .A(n_266), .Y(n_393) );
INVx2_ASAP7_75t_L g448 ( .A(n_266), .Y(n_448) );
INVx6_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g357 ( .A(n_267), .Y(n_357) );
BUFx3_ASAP7_75t_L g426 ( .A(n_267), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B1(n_273), .B2(n_274), .Y(n_268) );
INVx2_ASAP7_75t_L g528 ( .A(n_270), .Y(n_528) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g442 ( .A(n_271), .Y(n_442) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_271), .Y(n_605) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
BUFx2_ASAP7_75t_SL g480 ( .A(n_272), .Y(n_480) );
BUFx2_ASAP7_75t_SL g569 ( .A(n_272), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_274), .A2(n_391), .B1(n_392), .B2(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_293), .Y(n_277) );
OAI21xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_282), .B(n_283), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_279), .A2(n_413), .B(n_414), .Y(n_412) );
BUFx2_ASAP7_75t_L g473 ( .A(n_279), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_279), .A2(n_497), .B(n_498), .Y(n_496) );
INVx4_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
INVx2_ASAP7_75t_L g547 ( .A(n_280), .Y(n_547) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_280), .Y(n_586) );
AND2x4_ASAP7_75t_L g307 ( .A(n_281), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g339 ( .A(n_281), .Y(n_339) );
BUFx2_ASAP7_75t_L g375 ( .A(n_284), .Y(n_375) );
INVx4_ASAP7_75t_L g500 ( .A(n_284), .Y(n_500) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx4f_ASAP7_75t_SL g422 ( .A(n_285), .Y(n_422) );
BUFx2_ASAP7_75t_L g456 ( .A(n_285), .Y(n_456) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_285), .Y(n_470) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_285), .Y(n_578) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g292 ( .A(n_287), .Y(n_292) );
AND2x4_ASAP7_75t_L g291 ( .A(n_288), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g304 ( .A(n_288), .B(n_305), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_288), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g554 ( .A(n_289), .Y(n_554) );
BUFx4f_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g377 ( .A(n_290), .Y(n_377) );
BUFx12f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_291), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .C(n_301), .Y(n_293) );
BUFx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g453 ( .A(n_296), .Y(n_453) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_296), .Y(n_573) );
BUFx2_ASAP7_75t_L g592 ( .A(n_296), .Y(n_592) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g419 ( .A(n_299), .Y(n_419) );
INVx5_ASAP7_75t_L g451 ( .A(n_299), .Y(n_451) );
INVx2_ASAP7_75t_L g622 ( .A(n_299), .Y(n_622) );
INVx4_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g595 ( .A(n_303), .Y(n_595) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g471 ( .A(n_304), .Y(n_471) );
BUFx3_ASAP7_75t_L g506 ( .A(n_304), .Y(n_506) );
BUFx2_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_307), .Y(n_416) );
BUFx3_ASAP7_75t_L g619 ( .A(n_307), .Y(n_619) );
INVx1_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
INVx1_ASAP7_75t_L g459 ( .A(n_310), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_400), .B2(n_458), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_358), .B2(n_359), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND3x1_ASAP7_75t_L g319 ( .A(n_320), .B(n_341), .C(n_349), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_329), .C(n_333), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_326), .B2(n_327), .Y(n_321) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_324), .Y(n_367) );
INVx2_ASAP7_75t_L g542 ( .A(n_324), .Y(n_542) );
BUFx3_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_327), .A2(n_540), .B1(n_541), .B2(n_543), .Y(n_539) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx3_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_337), .B2(n_338), .Y(n_333) );
OAI22xp33_ASAP7_75t_SL g378 ( .A1(n_335), .A2(n_379), .B1(n_380), .B2(n_382), .Y(n_378) );
INVx4_ASAP7_75t_L g550 ( .A(n_335), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g381 ( .A(n_338), .Y(n_381) );
BUFx2_ASAP7_75t_L g556 ( .A(n_338), .Y(n_556) );
OR2x6_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_346), .Y(n_341) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g397 ( .A(n_345), .Y(n_397) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .Y(n_349) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g407 ( .A(n_352), .Y(n_407) );
BUFx3_ASAP7_75t_L g445 ( .A(n_352), .Y(n_445) );
BUFx3_ASAP7_75t_L g530 ( .A(n_352), .Y(n_530) );
INVx4_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g514 ( .A(n_356), .Y(n_514) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_383), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_371), .C(n_378), .Y(n_363) );
OAI22xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_368), .B1(n_369), .B2(n_370), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_373), .B(n_374), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_372), .A2(n_576), .B(n_577), .Y(n_575) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_390), .C(n_395), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g531 ( .A1(n_399), .A2(n_532), .B1(n_533), .B2(n_534), .C(n_535), .Y(n_531) );
INVx1_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_430), .B2(n_457), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
XOR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_429), .Y(n_403) );
NAND3x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_411), .C(n_423), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
NOR2x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_417), .Y(n_411) );
BUFx4f_ASAP7_75t_L g589 ( .A(n_415), .Y(n_589) );
INVx1_ASAP7_75t_SL g597 ( .A(n_416), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g545 ( .A(n_422), .Y(n_545) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
INVx3_ASAP7_75t_L g525 ( .A(n_426), .Y(n_525) );
INVx2_ASAP7_75t_L g457 ( .A(n_430), .Y(n_457) );
NAND4xp75_ASAP7_75t_L g431 ( .A(n_432), .B(n_440), .C(n_449), .D(n_455), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_438), .Y(n_432) );
INVx4_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g600 ( .A(n_435), .Y(n_600) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx4f_ASAP7_75t_SL g606 ( .A(n_445), .Y(n_606) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_450), .B(n_454), .Y(n_449) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_451), .Y(n_504) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g467 ( .A(n_453), .Y(n_467) );
INVx1_ASAP7_75t_L g488 ( .A(n_460), .Y(n_488) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g486 ( .A(n_463), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_464), .B(n_476), .Y(n_463) );
NOR2xp67_ASAP7_75t_SL g464 ( .A(n_465), .B(n_472), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .C(n_469), .Y(n_465) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_474), .B(n_475), .Y(n_472) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_482), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g636 ( .A(n_489), .Y(n_636) );
XNOR2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_611), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B1(n_516), .B2(n_610), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
XOR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_515), .Y(n_493) );
NAND3x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .C(n_511), .Y(n_494) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_501), .Y(n_495) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .C(n_505), .Y(n_501) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g610 ( .A(n_516), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_559), .B2(n_560), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g557 ( .A(n_520), .Y(n_557) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_521), .B(n_538), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
OAI221xp5_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_524), .B1(n_525), .B2(n_526), .C(n_527), .Y(n_522) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .C(n_552), .Y(n_538) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
OAI222xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_547), .B2(n_548), .C1(n_549), .C2(n_551), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_547), .A2(n_617), .B(n_618), .Y(n_616) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_552) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AO22x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_579), .B1(n_580), .B2(n_609), .Y(n_560) );
INVx1_ASAP7_75t_SL g609 ( .A(n_561), .Y(n_609) );
NOR4xp75_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .C(n_571), .D(n_575), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g608 ( .A(n_582), .Y(n_608) );
NAND3x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_598), .C(n_603), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_590), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B(n_588), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .C(n_594), .Y(n_590) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
XOR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_634), .Y(n_613) );
NAND2x1p5_ASAP7_75t_L g614 ( .A(n_615), .B(n_625), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .C(n_624), .Y(n_620) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_631), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_643), .Y(n_638) );
OR2x2_ASAP7_75t_SL g678 ( .A(n_639), .B(n_644), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_641), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_641), .B(n_668), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g668 ( .A(n_642), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OAI322xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_665), .A3(n_666), .B1(n_669), .B2(n_672), .C1(n_673), .C2(n_676), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND5xp2_ASAP7_75t_SL g654 ( .A(n_655), .B(n_656), .C(n_657), .D(n_660), .E(n_663), .Y(n_654) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
CKINVDCx16_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_677), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
endmodule