module fake_jpeg_29804_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_30),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_22),
.C(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_25),
.B1(n_12),
.B2(n_22),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_34),
.B(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_13),
.B1(n_28),
.B2(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_17),
.Y(n_46)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_13),
.B(n_16),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_32),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_33),
.C(n_29),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_54),
.Y(n_65)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_12),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_33),
.B(n_29),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_59),
.B(n_3),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_7),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_44),
.C(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_7),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_73),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_38),
.B1(n_35),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_55),
.B1(n_58),
.B2(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_38),
.C(n_23),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_89),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_38),
.B1(n_47),
.B2(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_45),
.C(n_57),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_75),
.C(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_45),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_78),
.B(n_67),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_65),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.C(n_92),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_45),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_107),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_97),
.B1(n_87),
.B2(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_88),
.C(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_86),
.C(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_98),
.C(n_104),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_90),
.B(n_47),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_90),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_113),
.B(n_64),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_3),
.B(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_4),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_53),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_4),
.A3(n_5),
.B1(n_108),
.B2(n_121),
.C(n_123),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_127),
.Y(n_129)
);


endmodule