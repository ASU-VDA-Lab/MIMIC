module fake_jpeg_5160_n_31 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_31);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_9),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_14),
.B1(n_15),
.B2(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.C(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_24),
.B(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_1),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_1),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_21),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_28),
.B(n_22),
.Y(n_30)
);

AOI321xp33_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_2),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.C(n_20),
.Y(n_31)
);


endmodule