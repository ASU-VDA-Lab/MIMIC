module fake_jpeg_6202_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_7),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_45),
.B(n_60),
.C(n_24),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_53),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_58),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_23),
.C(n_2),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_30),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_35),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_40),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_67),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_25),
.B1(n_49),
.B2(n_36),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_25),
.B1(n_36),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_25),
.B1(n_38),
.B2(n_36),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_38),
.B1(n_20),
.B2(n_33),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_74),
.B(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_20),
.B1(n_33),
.B2(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_20),
.B1(n_47),
.B2(n_28),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_40),
.B(n_39),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_29),
.B(n_55),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_89),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_24),
.B1(n_22),
.B2(n_27),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_95),
.B1(n_98),
.B2(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_16),
.B1(n_37),
.B2(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_31),
.B(n_39),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_37),
.B1(n_18),
.B2(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_107),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_39),
.B1(n_37),
.B2(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_37),
.B1(n_18),
.B2(n_32),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_43),
.A2(n_39),
.B1(n_40),
.B2(n_32),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_39),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_29),
.B1(n_32),
.B2(n_3),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_110),
.B(n_115),
.Y(n_160)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_2),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_123),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_94),
.B(n_55),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NOR4xp25_ASAP7_75t_SL g125 ( 
.A(n_77),
.B(n_10),
.C(n_4),
.D(n_6),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_91),
.B(n_68),
.C(n_96),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_137),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_4),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_99),
.B1(n_105),
.B2(n_104),
.Y(n_147)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_150),
.Y(n_184)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_80),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_113),
.C(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_89),
.B1(n_92),
.B2(n_70),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_159),
.B1(n_179),
.B2(n_128),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_100),
.B1(n_67),
.B2(n_64),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_162),
.Y(n_182)
);

INVx6_ASAP7_75t_SL g162 ( 
.A(n_123),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_118),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_173),
.Y(n_195)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_119),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_80),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_121),
.A2(n_107),
.B1(n_99),
.B2(n_90),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_170),
.B1(n_11),
.B2(n_13),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_83),
.B1(n_8),
.B2(n_9),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_29),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx6_ASAP7_75t_SL g173 ( 
.A(n_142),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_14),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_71),
.B(n_103),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_178),
.B(n_134),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_103),
.B(n_86),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_86),
.B1(n_8),
.B2(n_10),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_192),
.B1(n_198),
.B2(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_202),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_187),
.A2(n_189),
.B1(n_165),
.B2(n_177),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_139),
.B1(n_120),
.B2(n_133),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_133),
.C(n_120),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_190),
.B(n_208),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_143),
.B1(n_137),
.B2(n_124),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_117),
.C(n_124),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_213),
.C(n_179),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_119),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_193),
.B(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_138),
.B1(n_141),
.B2(n_135),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_151),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_13),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_14),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_172),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_160),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_153),
.B1(n_159),
.B2(n_154),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_161),
.C(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_231),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_239),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_171),
.B(n_149),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_230),
.B(n_234),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_186),
.B(n_195),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_191),
.C(n_182),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_168),
.B1(n_180),
.B2(n_148),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_225),
.A2(n_200),
.B1(n_212),
.B2(n_174),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_157),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_235),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_151),
.B(n_152),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_207),
.C(n_199),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_196),
.B(n_163),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_172),
.C(n_177),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_192),
.Y(n_247)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_200),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_172),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_187),
.B1(n_197),
.B2(n_198),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_250),
.B1(n_251),
.B2(n_261),
.Y(n_270)
);

CKINVDCx6p67_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_224),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_249),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_239),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_252),
.C(n_259),
.Y(n_262)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_197),
.B1(n_182),
.B2(n_203),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_191),
.B1(n_186),
.B2(n_214),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_195),
.C(n_188),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_215),
.B(n_221),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_204),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_275),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_274),
.B(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_230),
.C(n_236),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_235),
.C(n_226),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_278),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_244),
.A2(n_228),
.B1(n_223),
.B2(n_219),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_228),
.B1(n_240),
.B2(n_227),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_258),
.B1(n_253),
.B2(n_255),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_181),
.B1(n_271),
.B2(n_267),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_260),
.A2(n_218),
.B(n_216),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_254),
.B(n_174),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_174),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_248),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_278),
.Y(n_293)
);

OAI211xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_253),
.B(n_246),
.C(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_246),
.B(n_252),
.C(n_261),
.D(n_256),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_287),
.C(n_288),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_285),
.A2(n_266),
.B(n_262),
.Y(n_299)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_254),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_289),
.B(n_292),
.CI(n_181),
.CON(n_300),
.SN(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_262),
.C(n_270),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_301),
.C(n_303),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_290),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_181),
.B1(n_291),
.B2(n_292),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_287),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_294),
.B1(n_289),
.B2(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_281),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_281),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_283),
.C(n_282),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_298),
.B(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_310),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_319),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_305),
.A3(n_306),
.B1(n_309),
.B2(n_313),
.C1(n_300),
.C2(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_300),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_316),
.Y(n_326)
);


endmodule