module fake_jpeg_19776_n_9 (n_3, n_2, n_1, n_0, n_4, n_9);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_9;

wire n_8;
wire n_6;
wire n_5;
wire n_7;

OAI22xp5_ASAP7_75t_SL g5 ( 
.A1(n_2),
.A2(n_3),
.B1(n_0),
.B2(n_4),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

FAx1_ASAP7_75t_SL g7 ( 
.A(n_3),
.B(n_1),
.CI(n_0),
.CON(n_7),
.SN(n_7)
);

MAJIxp5_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_1),
.C(n_7),
.Y(n_8)
);

NAND4xp25_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_7),
.C(n_6),
.D(n_5),
.Y(n_9)
);


endmodule