module fake_jpeg_14167_n_490 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_490);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_490;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_62),
.Y(n_101)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_33),
.B1(n_36),
.B2(n_25),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_71),
.Y(n_107)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_37),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_78),
.Y(n_111)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_2),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_31),
.B(n_2),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_79),
.Y(n_116)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_86),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_3),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_92),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_95),
.Y(n_139)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_94),
.Y(n_140)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_31),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_41),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_98),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_100),
.B(n_123),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_102),
.A2(n_89),
.B1(n_91),
.B2(n_72),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_32),
.B1(n_36),
.B2(n_33),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_105),
.A2(n_137),
.B1(n_143),
.B2(n_155),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_36),
.B(n_40),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_101),
.C(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_87),
.B1(n_57),
.B2(n_77),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_117),
.B1(n_132),
.B2(n_147),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_50),
.B(n_47),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_41),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_125),
.B(n_153),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_48),
.B1(n_39),
.B2(n_30),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_32),
.B1(n_30),
.B2(n_40),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_58),
.B(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_151),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_51),
.A2(n_32),
.B1(n_48),
.B2(n_19),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_52),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_81),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_56),
.A2(n_48),
.B1(n_49),
.B2(n_19),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_60),
.A2(n_47),
.B1(n_45),
.B2(n_42),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_148),
.A2(n_49),
.B1(n_19),
.B2(n_81),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_45),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_42),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_74),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_8),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_49),
.B1(n_19),
.B2(n_21),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_102),
.A2(n_84),
.B1(n_82),
.B2(n_54),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_179),
.A3(n_204),
.B1(n_112),
.B2(n_144),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_63),
.B1(n_86),
.B2(n_85),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_158),
.A2(n_180),
.B1(n_185),
.B2(n_193),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_161),
.B(n_190),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_100),
.A2(n_98),
.B1(n_61),
.B2(n_76),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_162),
.A2(n_170),
.B1(n_178),
.B2(n_181),
.Y(n_229)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_74),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_138),
.C(n_145),
.Y(n_217)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_21),
.B1(n_24),
.B2(n_80),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_101),
.B(n_109),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_175),
.A2(n_119),
.B(n_15),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_73),
.B1(n_75),
.B2(n_69),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_101),
.A2(n_107),
.B(n_111),
.C(n_139),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_104),
.A2(n_92),
.B1(n_62),
.B2(n_49),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_64),
.B1(n_67),
.B2(n_79),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_49),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_122),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_121),
.A2(n_19),
.B1(n_79),
.B2(n_64),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_103),
.B1(n_144),
.B2(n_127),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_120),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_134),
.A2(n_152),
.B1(n_150),
.B2(n_128),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_196),
.Y(n_254)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

AO22x2_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_206),
.Y(n_225)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g199 ( 
.A(n_122),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_134),
.A2(n_16),
.B1(n_10),
.B2(n_12),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_200),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_253)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_112),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_209),
.B(n_208),
.Y(n_234)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_139),
.A2(n_9),
.B(n_10),
.C(n_13),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_9),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_207),
.Y(n_213)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_110),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_119),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_138),
.A2(n_9),
.B1(n_14),
.B2(n_15),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_138),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_211),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_219),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_217),
.B(n_215),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_152),
.B1(n_150),
.B2(n_135),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_236),
.B1(n_249),
.B2(n_162),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_234),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_159),
.B(n_104),
.C(n_103),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_242),
.C(n_157),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_207),
.A2(n_103),
.B1(n_127),
.B2(n_124),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_187),
.A2(n_118),
.B1(n_135),
.B2(n_128),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_166),
.A2(n_136),
.B(n_104),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_238),
.A2(n_201),
.B(n_185),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_251),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_124),
.C(n_118),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_167),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_231),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_202),
.A2(n_120),
.B1(n_129),
.B2(n_130),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_129),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_196),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_253),
.A2(n_209),
.B1(n_201),
.B2(n_198),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_119),
.B(n_130),
.C(n_14),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_240),
.B(n_238),
.C(n_254),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_266),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_261),
.A2(n_293),
.B(n_257),
.Y(n_334)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_265),
.A2(n_267),
.B1(n_282),
.B2(n_258),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_216),
.B(n_183),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_164),
.B1(n_210),
.B2(n_200),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_213),
.B(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_268),
.B(n_272),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_269),
.A2(n_302),
.B1(n_255),
.B2(n_290),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_188),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_270),
.B(n_275),
.Y(n_312)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_196),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_196),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_215),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_176),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_179),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_277),
.B(n_279),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_211),
.A2(n_157),
.A3(n_156),
.B1(n_160),
.B2(n_173),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_285),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_191),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_296),
.Y(n_308)
);

INVx2_ASAP7_75t_R g281 ( 
.A(n_223),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_281),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_157),
.B1(n_168),
.B2(n_184),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_234),
.A2(n_190),
.B(n_195),
.C(n_174),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_283),
.B(n_288),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_230),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_287),
.Y(n_321)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_182),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_290),
.A2(n_292),
.B(n_244),
.Y(n_315)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_295),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_240),
.A2(n_163),
.B(n_165),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_206),
.B(n_203),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx6_ASAP7_75t_SL g297 ( 
.A(n_244),
.Y(n_297)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

INVx13_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_229),
.A2(n_217),
.B1(n_254),
.B2(n_252),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_229),
.B1(n_254),
.B2(n_232),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_303),
.A2(n_304),
.B1(n_309),
.B2(n_323),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_265),
.A2(n_249),
.B1(n_233),
.B2(n_215),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_310),
.B(n_308),
.Y(n_350)
);

HAxp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_256),
.CON(n_311),
.SN(n_311)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_239),
.C(n_231),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_322),
.C(n_330),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_298),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_335),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_294),
.A2(n_246),
.B(n_239),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_318),
.A2(n_325),
.B(n_340),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_221),
.C(n_224),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_289),
.A2(n_246),
.B1(n_247),
.B2(n_214),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_294),
.A2(n_248),
.B(n_218),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_260),
.A2(n_267),
.B1(n_293),
.B2(n_274),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_328),
.A2(n_337),
.B1(n_304),
.B2(n_309),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_221),
.C(n_224),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_329),
.B(n_327),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_281),
.B(n_277),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_272),
.A2(n_214),
.B1(n_257),
.B2(n_218),
.Y(n_337)
);

INVx13_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_338),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_339),
.A2(n_318),
.B1(n_334),
.B2(n_340),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_292),
.A2(n_255),
.B(n_283),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_266),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_313),
.C(n_322),
.Y(n_372)
);

OAI32xp33_ASAP7_75t_L g342 ( 
.A1(n_305),
.A2(n_273),
.A3(n_278),
.B1(n_276),
.B2(n_263),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_343),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_339),
.A2(n_293),
.B1(n_282),
.B2(n_273),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_285),
.Y(n_344)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_344),
.Y(n_375)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_261),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_352),
.C(n_359),
.Y(n_389)
);

OAI22x1_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_259),
.B1(n_299),
.B2(n_281),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_355),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_310),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_262),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_354),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_305),
.A2(n_299),
.B1(n_276),
.B2(n_269),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_361),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_291),
.B1(n_286),
.B2(n_287),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_358),
.A2(n_326),
.B(n_314),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_295),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_367),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_316),
.A2(n_300),
.B1(n_301),
.B2(n_284),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_319),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_364),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_284),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_271),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_372),
.C(n_353),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_313),
.B1(n_330),
.B2(n_332),
.Y(n_380)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_320),
.A2(n_329),
.B1(n_312),
.B2(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_369),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_328),
.A2(n_303),
.B1(n_331),
.B2(n_327),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_366),
.A2(n_331),
.B1(n_322),
.B2(n_320),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_374),
.B(n_382),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_359),
.Y(n_404)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_312),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_381),
.B(n_387),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_344),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_330),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_390),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_325),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_337),
.Y(n_388)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_323),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_351),
.A2(n_326),
.B1(n_336),
.B2(n_324),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_363),
.B1(n_371),
.B2(n_362),
.Y(n_419)
);

NAND2x1p5_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_358),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_364),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_361),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_395),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_314),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_363),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_352),
.C(n_347),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_412),
.C(n_420),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_413),
.Y(n_433)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_365),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_409),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_351),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_376),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_422),
.Y(n_424)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_390),
.C(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_377),
.Y(n_415)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_342),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_397),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_417),
.A2(n_348),
.B(n_394),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_419),
.A2(n_391),
.B1(n_393),
.B2(n_392),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_371),
.C(n_355),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_370),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_349),
.C(n_343),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_385),
.C(n_378),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_429),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_421),
.A2(n_400),
.B1(n_378),
.B2(n_393),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_374),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_375),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_430),
.A2(n_435),
.B1(n_442),
.B2(n_437),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_402),
.A2(n_385),
.B(n_348),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_431),
.A2(n_417),
.B(n_423),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_405),
.A2(n_400),
.B1(n_382),
.B2(n_388),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_421),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_413),
.B(n_384),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_420),
.A2(n_397),
.B1(n_377),
.B2(n_386),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_402),
.B1(n_417),
.B2(n_386),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_440),
.B(n_441),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_384),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_439),
.B1(n_435),
.B2(n_438),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_442),
.B(n_415),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_445),
.B(n_451),
.Y(n_467)
);

BUFx24_ASAP7_75t_SL g446 ( 
.A(n_432),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_446),
.B(n_447),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_414),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_455),
.B(n_436),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_456),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_406),
.C(n_409),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_430),
.C(n_427),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_425),
.C(n_441),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_425),
.C(n_429),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_404),
.Y(n_456)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_451),
.C(n_448),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_440),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_463),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_426),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_462),
.B(n_452),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_468),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_455),
.A2(n_416),
.B(n_403),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_465),
.A2(n_412),
.B(n_443),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_433),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_306),
.C(n_338),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_475),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_470),
.B(n_474),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g478 ( 
.A1(n_471),
.A2(n_461),
.B(n_457),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_456),
.C(n_336),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_467),
.A2(n_314),
.B(n_306),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_476),
.B(n_466),
.C(n_338),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_478),
.B(n_479),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_472),
.A2(n_458),
.B1(n_460),
.B2(n_457),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_481),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_SL g485 ( 
.A1(n_482),
.A2(n_477),
.B(n_473),
.C(n_333),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_482),
.C(n_473),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_487),
.B(n_484),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_483),
.A2(n_480),
.B(n_306),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_333),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_333),
.Y(n_490)
);


endmodule