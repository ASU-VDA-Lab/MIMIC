module fake_jpeg_31311_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_13),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_18),
.Y(n_80)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_18),
.B1(n_17),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_28),
.B1(n_34),
.B2(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_68),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_75),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_31),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_19),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_34),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_49),
.B1(n_48),
.B2(n_38),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_87),
.B1(n_91),
.B2(n_58),
.Y(n_121)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_87)
);

AO22x2_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_54),
.B(n_79),
.C(n_60),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_77),
.B1(n_53),
.B2(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_94),
.B1(n_101),
.B2(n_102),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_5),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_82),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_57),
.C(n_58),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_56),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_85),
.B(n_108),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_5),
.B(n_6),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_122),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_79),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_84),
.B1(n_100),
.B2(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_54),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_129),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_107),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_134),
.B1(n_143),
.B2(n_123),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_97),
.B(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_129),
.B(n_109),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_81),
.B1(n_96),
.B2(n_92),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_81),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_122),
.B(n_109),
.Y(n_150)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_134),
.A3(n_139),
.B1(n_113),
.B2(n_117),
.C1(n_120),
.C2(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_112),
.C(n_130),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_161),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_162),
.B1(n_164),
.B2(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_110),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_126),
.B1(n_123),
.B2(n_116),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_120),
.B1(n_124),
.B2(n_117),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_142),
.B(n_135),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_135),
.B(n_149),
.C(n_132),
.D(n_137),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_153),
.C(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

AO221x1_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_124),
.B1(n_141),
.B2(n_138),
.C(n_133),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_134),
.B1(n_163),
.B2(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_158),
.B1(n_159),
.B2(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_159),
.B1(n_153),
.B2(n_105),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_167),
.B(n_166),
.C(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_178),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_168),
.B(n_159),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_181),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_194),
.B(n_10),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_190),
.B1(n_183),
.B2(n_177),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_86),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_199),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_200),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_10),
.C(n_7),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.C(n_193),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_197),
.C(n_196),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_7),
.Y(n_206)
);


endmodule