module fake_jpeg_4104_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_67),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_69),
.B1(n_59),
.B2(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_61),
.B1(n_56),
.B2(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_76),
.B1(n_50),
.B2(n_55),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_79),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_46),
.B1(n_44),
.B2(n_71),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_53),
.C(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_76),
.B1(n_71),
.B2(n_58),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_58),
.A3(n_17),
.B1(n_19),
.B2(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_13),
.B1(n_42),
.B2(n_32),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_85),
.Y(n_88)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_0),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_11),
.C(n_28),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_90),
.B(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_93),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_88),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_7),
.C2(n_8),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_15),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_12),
.C(n_26),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_10),
.A3(n_24),
.B1(n_21),
.B2(n_20),
.C1(n_9),
.C2(n_43),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_1),
.Y(n_102)
);


endmodule