module fake_jpeg_20370_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_24),
.Y(n_27)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_24),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_10),
.B1(n_12),
.B2(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_19),
.B(n_18),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_20),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_9),
.B(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_20),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_13),
.B(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_36),
.C(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.C(n_41),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.C(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_51),
.B1(n_21),
.B2(n_23),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_39),
.C(n_34),
.Y(n_57)
);

OA21x2_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_50),
.B(n_49),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_60),
.B(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_61),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_1),
.B(n_2),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_62),
.C(n_20),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.C(n_23),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_20),
.C(n_12),
.Y(n_68)
);

A2O1A1O1Ixp25_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B(n_7),
.C(n_3),
.D(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_1),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);


endmodule