module fake_jpeg_9893_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_17),
.B1(n_33),
.B2(n_20),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_17),
.B1(n_33),
.B2(n_28),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_56),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_17),
.B1(n_20),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_67),
.B1(n_32),
.B2(n_18),
.Y(n_74)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_28),
.B1(n_33),
.B2(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_42),
.B1(n_45),
.B2(n_40),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_78),
.B1(n_97),
.B2(n_50),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_44),
.B1(n_32),
.B2(n_47),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_81),
.B1(n_95),
.B2(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_93),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_40),
.B1(n_45),
.B2(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_32),
.B1(n_30),
.B2(n_25),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_47),
.B1(n_46),
.B2(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_46),
.B1(n_36),
.B2(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_25),
.B1(n_30),
.B2(n_35),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_37),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_64),
.C(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_36),
.B1(n_30),
.B2(n_21),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_115),
.C(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_65),
.B1(n_68),
.B2(n_62),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_77),
.B1(n_71),
.B2(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_22),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_108),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_62),
.B1(n_64),
.B2(n_59),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_114),
.B1(n_121),
.B2(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_125),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_116),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_59),
.B(n_50),
.C(n_64),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_74),
.B(n_77),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_70),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_121),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_123),
.B1(n_126),
.B2(n_87),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_48),
.B1(n_11),
.B2(n_16),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_75),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_149),
.B(n_114),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_134),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_130),
.B(n_138),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_92),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_14),
.C(n_15),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_143),
.B1(n_144),
.B2(n_152),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_71),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_71),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_140),
.C(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_107),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_38),
.C(n_84),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_19),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_145),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_83),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_58),
.B1(n_29),
.B2(n_26),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_29),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_23),
.C(n_26),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_29),
.B(n_26),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_105),
.Y(n_177)
);

NOR2x1_ASAP7_75t_R g157 ( 
.A(n_139),
.B(n_115),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_175),
.B(n_149),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_115),
.B(n_125),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_158),
.A2(n_167),
.B(n_168),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_165),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_115),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_107),
.B1(n_118),
.B2(n_110),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_178),
.B1(n_180),
.B2(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_172),
.C(n_181),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_111),
.B(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_104),
.B1(n_123),
.B2(n_109),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_140),
.B1(n_145),
.B2(n_141),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_120),
.C(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_112),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_136),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_136),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_185),
.B(n_176),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_146),
.B1(n_151),
.B2(n_119),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_194),
.B1(n_200),
.B2(n_160),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_167),
.B(n_156),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_130),
.B(n_146),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_161),
.B(n_167),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_146),
.B1(n_119),
.B2(n_109),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_130),
.B1(n_109),
.B2(n_116),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_198),
.B1(n_201),
.B2(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_157),
.A2(n_116),
.B1(n_120),
.B2(n_119),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_162),
.A2(n_116),
.B1(n_26),
.B2(n_19),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_206),
.Y(n_219)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_212),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_156),
.B1(n_178),
.B2(n_169),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_166),
.C(n_172),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_234),
.C(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_221),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_231),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_198),
.B1(n_207),
.B2(n_206),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_236),
.C(n_240),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_171),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_239),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_166),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_193),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_180),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_0),
.C(n_1),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_1),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_15),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_209),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_3),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_196),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_249),
.B1(n_256),
.B2(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_211),
.C(n_200),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_254),
.C(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_194),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_210),
.B1(n_195),
.B2(n_191),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_234),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_216),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_211),
.C(n_197),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_189),
.B1(n_192),
.B2(n_186),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_186),
.B1(n_12),
.B2(n_9),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_8),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_219),
.B(n_230),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_264),
.A2(n_267),
.B(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_219),
.B(n_217),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_276),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_225),
.C(n_226),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_254),
.C(n_245),
.Y(n_288)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_287)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_248),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_228),
.B1(n_215),
.B2(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_224),
.B1(n_236),
.B2(n_237),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_246),
.A2(n_239),
.B(n_235),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_266),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_282),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_295),
.C(n_273),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_277),
.B1(n_268),
.B2(n_274),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_253),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_253),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_255),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_293),
.A2(n_284),
.B(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_279),
.B1(n_266),
.B2(n_276),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_305),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_302),
.B(n_294),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_281),
.A2(n_269),
.B(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_271),
.C(n_280),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_265),
.B1(n_263),
.B2(n_5),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_4),
.Y(n_311)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_9),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_9),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_316),
.B(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_317),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_4),
.B(n_5),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_4),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_310),
.B(n_297),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_301),
.C(n_6),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_6),
.C(n_7),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_301),
.Y(n_332)
);

NAND4xp25_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_330),
.C(n_326),
.D(n_325),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_331),
.B(n_323),
.Y(n_334)
);

OAI211xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_327),
.B(n_324),
.C(n_7),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_6),
.B(n_7),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_7),
.Y(n_337)
);


endmodule