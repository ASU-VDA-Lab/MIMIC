module fake_netlist_1_12348_n_668 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_668, n_669);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_668;
output n_669;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g88 ( .A(n_70), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_31), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_2), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_73), .Y(n_92) );
INVx2_ASAP7_75t_SL g93 ( .A(n_7), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_28), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_7), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_34), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_64), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_2), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_10), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_67), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_25), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_48), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_23), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_29), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_21), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_78), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_61), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_84), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_47), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_43), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_38), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_76), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_27), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_10), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_77), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_45), .Y(n_125) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_69), .B(n_58), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_52), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_32), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_74), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_85), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_35), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_132), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_132), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_112), .B(n_0), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_112), .B(n_0), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
OR2x2_ASAP7_75t_L g141 ( .A(n_90), .B(n_98), .Y(n_141) );
BUFx8_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_91), .A2(n_50), .B(n_83), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_132), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_132), .Y(n_147) );
AOI22xp5_ASAP7_75t_SL g148 ( .A1(n_100), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_148) );
INVx2_ASAP7_75t_SL g149 ( .A(n_129), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
XOR2xp5_ASAP7_75t_L g151 ( .A(n_104), .B(n_1), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx2_ASAP7_75t_SL g153 ( .A(n_142), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_142), .B(n_107), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_134), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
OR2x2_ASAP7_75t_L g162 ( .A(n_149), .B(n_95), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_149), .B(n_125), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_137), .A2(n_113), .B1(n_119), .B2(n_106), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_149), .B(n_102), .Y(n_169) );
BUFx8_ASAP7_75t_SL g170 ( .A(n_137), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_136), .B(n_110), .Y(n_171) );
INVx1_ASAP7_75t_SL g172 ( .A(n_141), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_142), .B(n_93), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_141), .B(n_98), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_172), .A2(n_137), .B1(n_142), .B2(n_139), .Y(n_178) );
OR2x6_ASAP7_75t_L g179 ( .A(n_153), .B(n_139), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_172), .B(n_136), .Y(n_180) );
INVxp67_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_158), .A2(n_150), .B1(n_143), .B2(n_144), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_158), .A2(n_150), .B1(n_143), .B2(n_144), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_169), .B(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_157), .B(n_138), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_157), .B(n_138), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_157), .B(n_138), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_157), .B(n_94), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_155), .B(n_97), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_173), .B(n_92), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_93), .B1(n_99), .B2(n_108), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_165), .B(n_96), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_162), .B(n_105), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_174), .B(n_111), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_174), .B(n_117), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_155), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_154), .B(n_128), .Y(n_200) );
BUFx12f_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_156), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_156), .A2(n_99), .B1(n_122), .B2(n_115), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_171), .B(n_130), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_161), .B(n_101), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_171), .B(n_101), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_167), .B(n_103), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_161), .B(n_103), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_166), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_166), .B(n_109), .Y(n_211) );
AND2x6_ASAP7_75t_SL g212 ( .A(n_175), .B(n_151), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_181), .B(n_151), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_187), .A2(n_189), .B(n_188), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_187), .A2(n_177), .B(n_176), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_191), .B(n_175), .Y(n_216) );
AOI21x1_ASAP7_75t_L g217 ( .A1(n_211), .A2(n_177), .B(n_176), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_186), .B(n_151), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_188), .A2(n_145), .B(n_164), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_189), .Y(n_221) );
OAI21x1_ASAP7_75t_SL g222 ( .A1(n_178), .A2(n_145), .B(n_109), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_208), .B(n_148), .Y(n_223) );
OR2x6_ASAP7_75t_SL g224 ( .A(n_201), .B(n_148), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_205), .B(n_108), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_180), .B(n_115), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_190), .A2(n_145), .B(n_164), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_197), .B(n_122), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_196), .B(n_114), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_191), .B(n_114), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_198), .B(n_118), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_178), .A2(n_124), .B1(n_121), .B2(n_118), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_179), .A2(n_124), .B1(n_121), .B2(n_120), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_190), .A2(n_145), .B(n_164), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_184), .A2(n_120), .B1(n_110), .B2(n_123), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_185), .B(n_116), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_183), .A2(n_145), .B(n_163), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_204), .B(n_116), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_183), .A2(n_168), .B(n_163), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_210), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_199), .A2(n_168), .B(n_163), .Y(n_241) );
OAI22x1_ASAP7_75t_L g242 ( .A1(n_212), .A2(n_123), .B1(n_131), .B2(n_6), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_210), .B(n_131), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_200), .B(n_4), .Y(n_244) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_232), .A2(n_211), .B(n_147), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_237), .A2(n_192), .B(n_209), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
BUFx4f_ASAP7_75t_SL g248 ( .A(n_213), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_240), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_216), .A2(n_199), .B(n_179), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_192), .B(n_202), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_220), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_240), .B(n_210), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_230), .A2(n_179), .B(n_182), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_222), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_229), .A2(n_207), .B(n_206), .C(n_202), .Y(n_261) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_227), .A2(n_126), .B(n_133), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_234), .A2(n_179), .B(n_182), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_239), .A2(n_179), .B(n_182), .Y(n_264) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_146), .A3(n_133), .B(n_147), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_220), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_223), .B(n_194), .Y(n_267) );
NAND3xp33_ASAP7_75t_L g268 ( .A(n_233), .B(n_203), .C(n_135), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_202), .B(n_193), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_260), .B(n_225), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_260), .B(n_226), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_249), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_249), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_252), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_248), .Y(n_275) );
OAI21x1_ASAP7_75t_SL g276 ( .A1(n_247), .A2(n_235), .B(n_238), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_252), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_256), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_267), .B(n_218), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_247), .Y(n_280) );
BUFx8_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_253), .B(n_231), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_263), .A2(n_243), .B(n_235), .Y(n_283) );
INVx4_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_244), .B(n_228), .C(n_236), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_246), .A2(n_202), .B(n_133), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_246), .A2(n_147), .B(n_146), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_259), .A2(n_146), .B(n_160), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_253), .B(n_242), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_254), .A2(n_195), .B(n_159), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_245), .B(n_224), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_276), .A2(n_262), .B(n_245), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_247), .Y(n_293) );
AOI21x1_ASAP7_75t_L g294 ( .A1(n_276), .A2(n_259), .B(n_264), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_286), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_289), .A2(n_262), .B(n_259), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_285), .A2(n_268), .B(n_258), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_274), .B(n_262), .Y(n_301) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_289), .A2(n_268), .B(n_251), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_274), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_272), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_272), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_287), .A2(n_269), .B(n_250), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_287), .A2(n_269), .B(n_250), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_273), .B(n_271), .Y(n_310) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_286), .A2(n_250), .B(n_257), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_284), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_273), .B(n_265), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_291), .B(n_265), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_290), .A2(n_265), .B(n_160), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_299), .B(n_284), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_305), .B(n_265), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_305), .B(n_288), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_305), .B(n_265), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_316), .B(n_291), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_319), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_316), .B(n_282), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_301), .B(n_265), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_316), .B(n_271), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_299), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_301), .B(n_283), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_319), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_303), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_306), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_306), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_298), .Y(n_347) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_300), .A2(n_290), .B(n_288), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_301), .B(n_293), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_301), .B(n_283), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_293), .B(n_278), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_312), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_293), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_293), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_319), .A2(n_279), .B1(n_270), .B2(n_278), .Y(n_361) );
OR2x2_ASAP7_75t_SL g362 ( .A(n_312), .B(n_275), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_315), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_294), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_349), .B(n_315), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_349), .B(n_315), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_349), .B(n_315), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_362), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_332), .B(n_317), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_363), .B(n_297), .Y(n_371) );
INVx5_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
NOR2xp67_ASAP7_75t_L g373 ( .A(n_355), .B(n_312), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_332), .B(n_317), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_331), .B(n_297), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_331), .B(n_297), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_327), .B(n_310), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_338), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_324), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_297), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_360), .B(n_310), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_341), .B(n_297), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_341), .B(n_292), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_341), .B(n_351), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_333), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_333), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_360), .B(n_279), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_351), .B(n_292), .Y(n_388) );
NAND2x1p5_ASAP7_75t_L g389 ( .A(n_355), .B(n_313), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_340), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_340), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_345), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_355), .A2(n_314), .B1(n_313), .B2(n_201), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_327), .B(n_314), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_358), .B(n_314), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_355), .B(n_314), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_351), .B(n_292), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_345), .B(n_302), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_338), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_329), .B(n_302), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_292), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_329), .B(n_302), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_329), .B(n_302), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_328), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_358), .B(n_292), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_350), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_354), .B(n_270), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_326), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_354), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_359), .B(n_318), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_353), .B(n_318), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_328), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_359), .B(n_318), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_353), .B(n_318), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_353), .B(n_318), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_336), .B(n_256), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_362), .B(n_5), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_321), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_343), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_321), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_334), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_352), .B(n_294), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_365), .B(n_321), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_365), .B(n_321), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_371), .B(n_334), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_422), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_367), .B(n_321), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_367), .B(n_344), .Y(n_433) );
AND2x4_ASAP7_75t_SL g434 ( .A(n_421), .B(n_352), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_368), .B(n_384), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_369), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_372), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_368), .B(n_336), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_373), .B(n_352), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_371), .B(n_337), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_414), .B(n_357), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_411), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_414), .B(n_352), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_395), .B(n_337), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_425), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_417), .B(n_356), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_372), .B(n_356), .Y(n_448) );
NOR2x1_ASAP7_75t_SL g449 ( .A(n_372), .B(n_339), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_370), .B(n_356), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_375), .B(n_322), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_420), .B(n_361), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_417), .B(n_356), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_378), .B(n_326), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_375), .B(n_322), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_425), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_376), .B(n_322), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_385), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_386), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_390), .Y(n_461) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_421), .B(n_423), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_380), .B(n_325), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_392), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_372), .B(n_326), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_380), .B(n_325), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_393), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_383), .B(n_330), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_382), .B(n_330), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_383), .B(n_335), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_388), .B(n_335), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_401), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_421), .B(n_364), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_407), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_409), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_412), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_400), .B(n_335), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_374), .B(n_342), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_388), .B(n_342), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_398), .B(n_342), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_391), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_391), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_424), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_398), .B(n_347), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_420), .B(n_361), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_381), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_377), .B(n_347), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_415), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_415), .B(n_347), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_377), .B(n_323), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_396), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_410), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_389), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_389), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_387), .B(n_5), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_418), .B(n_323), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_406), .B(n_323), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_405), .B(n_323), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_397), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_435), .B(n_402), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_493), .B(n_403), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_429), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_437), .B(n_394), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_433), .B(n_404), .Y(n_507) );
NOR2xp33_ASAP7_75t_SL g508 ( .A(n_437), .B(n_397), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_487), .B(n_408), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_451), .B(n_413), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_451), .B(n_416), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_455), .B(n_408), .Y(n_513) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_465), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_431), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_452), .B(n_201), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_426), .B(n_399), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_455), .B(n_364), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g520 ( .A1(n_496), .A2(n_348), .B(n_300), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_458), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_461), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_464), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_467), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_496), .B(n_281), .C(n_152), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_457), .B(n_419), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_452), .A2(n_419), .B1(n_296), .B2(n_294), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_446), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_436), .B(n_281), .C(n_140), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_430), .B(n_348), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_427), .B(n_348), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_432), .B(n_296), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_476), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_430), .B(n_308), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_484), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_446), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_459), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_459), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_486), .B(n_6), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_448), .B(n_296), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_436), .B(n_8), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_472), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_489), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_440), .B(n_308), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_472), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_438), .B(n_296), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_444), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_483), .B(n_281), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_478), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_488), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g556 ( .A1(n_494), .A2(n_127), .A3(n_266), .B1(n_256), .B2(n_13), .Y(n_556) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_465), .B(n_311), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_448), .B(n_296), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_440), .B(n_488), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_456), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_491), .A2(n_311), .B1(n_296), .B2(n_308), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_463), .B(n_308), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_441), .B(n_308), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_448), .B(n_311), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_456), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_450), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_463), .B(n_309), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_466), .B(n_309), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_555), .B(n_466), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_520), .A2(n_468), .B1(n_443), .B2(n_447), .C(n_453), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_501), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_516), .B(n_500), .C(n_495), .Y(n_572) );
AOI21xp33_ASAP7_75t_L g573 ( .A1(n_543), .A2(n_483), .B(n_462), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_559), .B(n_469), .Y(n_574) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_531), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_526), .A2(n_498), .B1(n_480), .B2(n_470), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_547), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_553), .B(n_551), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_513), .B(n_468), .Y(n_579) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_515), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_526), .A2(n_439), .B(n_473), .Y(n_581) );
AOI322xp5_ASAP7_75t_L g582 ( .A1(n_506), .A2(n_485), .A3(n_471), .B1(n_479), .B2(n_439), .C1(n_482), .C2(n_492), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_508), .A2(n_499), .B1(n_497), .B2(n_492), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_531), .A2(n_482), .B1(n_473), .B2(n_434), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_521), .Y(n_585) );
O2A1O1Ixp33_ASAP7_75t_SL g586 ( .A1(n_539), .A2(n_434), .B(n_445), .C(n_442), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_554), .B(n_442), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_517), .B(n_445), .Y(n_588) );
NOR4xp25_ASAP7_75t_SL g589 ( .A(n_514), .B(n_9), .C(n_11), .D(n_12), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_545), .A2(n_9), .B(n_11), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_505), .A2(n_309), .B1(n_255), .B2(n_152), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_540), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_520), .A2(n_140), .B1(n_152), .B2(n_14), .C(n_15), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_547), .B(n_12), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_511), .B(n_309), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_512), .B(n_309), .Y(n_598) );
XOR2x2_ASAP7_75t_L g599 ( .A(n_552), .B(n_13), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_508), .B(n_140), .C(n_152), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_527), .Y(n_601) );
NOR2xp33_ASAP7_75t_SL g602 ( .A(n_504), .B(n_255), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_524), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_556), .B(n_14), .C(n_15), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_564), .B(n_311), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_564), .B(n_16), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_558), .A2(n_255), .B1(n_152), .B2(n_140), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_557), .B(n_140), .C(n_255), .Y(n_609) );
OAI211xp5_ASAP7_75t_L g610 ( .A1(n_561), .A2(n_18), .B(n_19), .C(n_20), .Y(n_610) );
AOI321xp33_ASAP7_75t_L g611 ( .A1(n_572), .A2(n_529), .A3(n_561), .B1(n_533), .B2(n_532), .C(n_568), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_570), .B(n_503), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_575), .A2(n_529), .B(n_558), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_582), .A2(n_510), .B1(n_536), .B2(n_534), .C(n_538), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_582), .B(n_605), .C(n_595), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_583), .A2(n_528), .B1(n_525), .B2(n_566), .C(n_560), .Y(n_616) );
NAND4xp75_ASAP7_75t_L g617 ( .A(n_573), .B(n_567), .C(n_563), .D(n_537), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_581), .A2(n_518), .B1(n_562), .B2(n_507), .C(n_502), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_591), .A2(n_548), .B(n_541), .C(n_549), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g620 ( .A1(n_576), .A2(n_535), .B1(n_550), .B2(n_519), .C(n_509), .Y(n_620) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_584), .B(n_565), .C(n_546), .D(n_542), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_577), .A2(n_544), .B1(n_19), .B2(n_20), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_569), .B(n_544), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_578), .A2(n_18), .B1(n_21), .B2(n_168), .C(n_160), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_580), .B(n_22), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_601), .B(n_24), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g627 ( .A1(n_600), .A2(n_26), .B(n_30), .Y(n_627) );
NAND2xp33_ASAP7_75t_SL g628 ( .A(n_607), .B(n_33), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_599), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_607), .A2(n_36), .B1(n_37), .B2(n_41), .C1(n_42), .C2(n_44), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_594), .B(n_46), .C(n_49), .D(n_51), .Y(n_631) );
AOI322xp5_ASAP7_75t_L g632 ( .A1(n_574), .A2(n_53), .A3(n_55), .B1(n_56), .B2(n_57), .C1(n_59), .C2(n_60), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_587), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_586), .A2(n_63), .B1(n_65), .B2(n_66), .C(n_68), .Y(n_635) );
NOR2xp67_ASAP7_75t_L g636 ( .A(n_600), .B(n_72), .Y(n_636) );
OAI31xp33_ASAP7_75t_L g637 ( .A1(n_610), .A2(n_79), .A3(n_80), .B(n_82), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_596), .A2(n_86), .B1(n_598), .B2(n_585), .C(n_597), .Y(n_638) );
NAND4xp25_ASAP7_75t_SL g639 ( .A(n_609), .B(n_608), .C(n_579), .D(n_588), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_603), .A2(n_604), .B(n_592), .C(n_606), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_589), .B(n_606), .C(n_602), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_590), .A2(n_575), .B(n_573), .C(n_586), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_593), .A2(n_570), .B1(n_572), .B2(n_583), .C(n_543), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_586), .A2(n_575), .B(n_506), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_633), .Y(n_645) );
NAND4xp75_ASAP7_75t_L g646 ( .A(n_644), .B(n_625), .C(n_622), .D(n_613), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_612), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_615), .A2(n_629), .B1(n_614), .B2(n_643), .C(n_613), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_642), .B(n_616), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g650 ( .A(n_620), .B(n_619), .C(n_611), .D(n_639), .Y(n_650) );
NOR2xp33_ASAP7_75t_SL g651 ( .A(n_635), .B(n_636), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_641), .B(n_637), .C(n_628), .D(n_631), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_649), .B(n_634), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_650), .B(n_640), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g655 ( .A(n_648), .B(n_627), .C(n_619), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_648), .B(n_630), .C(n_624), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_653), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_654), .B(n_647), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_656), .B(n_646), .Y(n_659) );
NAND2xp33_ASAP7_75t_R g660 ( .A(n_659), .B(n_655), .Y(n_660) );
INVx3_ASAP7_75t_SL g661 ( .A(n_658), .Y(n_661) );
OAI22x1_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_658), .B1(n_657), .B2(n_645), .Y(n_662) );
AND2x2_ASAP7_75t_SL g663 ( .A(n_660), .B(n_657), .Y(n_663) );
XOR2xp5_ASAP7_75t_L g664 ( .A(n_662), .B(n_652), .Y(n_664) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_663), .B(n_621), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_664), .A2(n_651), .B1(n_626), .B2(n_618), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_665), .B(n_632), .Y(n_667) );
UNKNOWN g668 ( );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_617), .B1(n_638), .B2(n_623), .Y(n_669) );
endmodule