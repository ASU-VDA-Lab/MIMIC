module fake_ibex_1590_n_988 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_988);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_988;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_510;
wire n_418;
wire n_193;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_899;
wire n_843;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_597;
wire n_415;
wire n_285;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_955;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_912;
wire n_874;
wire n_921;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_99),
.B(n_2),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_105),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_31),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_41),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_31),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_33),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_87),
.B(n_126),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_76),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_119),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_72),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_25),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_60),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_149),
.B(n_122),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_153),
.B(n_46),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_8),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_35),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_38),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_117),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_93),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_84),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_68),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_4),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_163),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_106),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_120),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_63),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_184),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_132),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_186),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_90),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_61),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_168),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_75),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_56),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_139),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_1),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_94),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_28),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_136),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_152),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_32),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_112),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_155),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_66),
.B(n_24),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_171),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_10),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_57),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_160),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_52),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_103),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_162),
.B(n_174),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_140),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_64),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_28),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_109),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_154),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_91),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_39),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_176),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_111),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_49),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_80),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_150),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_125),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_133),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_29),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_32),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_67),
.B(n_145),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_71),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_44),
.B(n_86),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_11),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_24),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_185),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_121),
.B(n_147),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_108),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_3),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_96),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_45),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_161),
.B(n_124),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_227),
.B(n_0),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_227),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_264),
.B1(n_272),
.B2(n_197),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_227),
.B(n_0),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_211),
.A2(n_89),
.B(n_182),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_2),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_228),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_229),
.B(n_303),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_4),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_197),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_245),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_213),
.B(n_5),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_221),
.B(n_6),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_221),
.B(n_7),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_211),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_240),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_212),
.B(n_10),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_258),
.B(n_12),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_258),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_243),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_252),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_217),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g350 ( 
.A1(n_252),
.A2(n_92),
.B(n_181),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

BUFx12f_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_264),
.B(n_12),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_272),
.B(n_14),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_265),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_260),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_269),
.B(n_62),
.Y(n_361)
);

CKINVDCx6p67_ASAP7_75t_R g362 ( 
.A(n_193),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_191),
.B(n_16),
.Y(n_367)
);

BUFx8_ASAP7_75t_SL g368 ( 
.A(n_188),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_274),
.B(n_18),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_280),
.B(n_18),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_280),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_255),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_291),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_198),
.B(n_19),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_203),
.B(n_20),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_205),
.B(n_21),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_255),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_190),
.Y(n_380)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_192),
.B(n_65),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_195),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_206),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_255),
.Y(n_384)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_255),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_200),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_209),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_218),
.B(n_21),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_201),
.A2(n_98),
.B(n_178),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_219),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_202),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_215),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_216),
.A2(n_97),
.B(n_175),
.Y(n_393)
);

OAI22x1_ASAP7_75t_L g394 ( 
.A1(n_271),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_279),
.Y(n_395)
);

CKINVDCx8_ASAP7_75t_R g396 ( 
.A(n_194),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_285),
.B(n_22),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_222),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_316),
.B(n_224),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_329),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_321),
.B(n_380),
.Y(n_403)
);

NOR2x1p5_ASAP7_75t_L g404 ( 
.A(n_325),
.B(n_286),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_321),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_355),
.Y(n_409)
);

CKINVDCx11_ASAP7_75t_R g410 ( 
.A(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_226),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_355),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_328),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_318),
.B(n_196),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_330),
.B(n_204),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_318),
.B(n_312),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_322),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_339),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_339),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

CKINVDCx6p67_ASAP7_75t_R g435 ( 
.A(n_362),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_235),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g437 ( 
.A(n_341),
.B(n_193),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_329),
.A2(n_225),
.B1(n_232),
.B2(n_249),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_333),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_349),
.B(n_283),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_385),
.B(n_241),
.C(n_234),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_334),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_331),
.B(n_289),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_341),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_342),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_334),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_331),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_331),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_331),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_343),
.B(n_189),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_381),
.B(n_208),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_343),
.Y(n_459)
);

AND3x2_ASAP7_75t_L g460 ( 
.A(n_376),
.B(n_259),
.C(n_223),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_348),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_348),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_348),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_336),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_336),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_320),
.B(n_242),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_336),
.B(n_236),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_394),
.B(n_210),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_336),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_336),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

BUFx6f_ASAP7_75t_SL g474 ( 
.A(n_376),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_363),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_388),
.A2(n_397),
.B1(n_377),
.B2(n_387),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_319),
.B(n_387),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_359),
.B(n_210),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

BUFx4f_ASAP7_75t_L g482 ( 
.A(n_397),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_SL g483 ( 
.A(n_394),
.B(n_225),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_363),
.A2(n_244),
.B1(n_249),
.B2(n_232),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_351),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_363),
.B(n_302),
.C(n_256),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_398),
.B(n_263),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_346),
.B(n_358),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_345),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_356),
.B(n_267),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_398),
.B(n_277),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_345),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_357),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_353),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_364),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_364),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_396),
.B(n_261),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_383),
.B(n_395),
.C(n_390),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_367),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_353),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_L g501 ( 
.A(n_378),
.B(n_306),
.C(n_304),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_382),
.B(n_282),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_372),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_398),
.B(n_287),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_372),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_364),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_366),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_365),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_366),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_386),
.B(n_261),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_350),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_366),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_369),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_360),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_482),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_386),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_499),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_391),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_423),
.B(n_375),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_426),
.B(n_270),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_423),
.B(n_270),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_244),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_429),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_427),
.B(n_188),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_426),
.B(n_273),
.Y(n_527)
);

BUFx5_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_476),
.B(n_199),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_434),
.B(n_275),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_482),
.B(n_278),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_410),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_508),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_375),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_448),
.B(n_421),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_375),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_436),
.B(n_443),
.Y(n_538)
);

O2A1O1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_425),
.A2(n_327),
.B(n_324),
.C(n_340),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_436),
.B(n_324),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_513),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_477),
.B(n_340),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_417),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_419),
.A2(n_361),
.B1(n_315),
.B2(n_314),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_404),
.B(n_310),
.Y(n_546)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_444),
.B(n_373),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_462),
.B(n_373),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_473),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_475),
.B(n_230),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_233),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_474),
.A2(n_199),
.B1(n_214),
.B2(n_361),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_400),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_481),
.B(n_238),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_451),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_501),
.B(n_288),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_490),
.B(n_301),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_420),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_497),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_422),
.A2(n_361),
.B1(n_314),
.B2(n_315),
.Y(n_561)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_399),
.B(n_290),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_478),
.B(n_239),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_452),
.B(n_361),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_424),
.B(n_326),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_402),
.B(n_247),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_430),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_489),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_457),
.B(n_250),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_432),
.A2(n_344),
.B1(n_335),
.B2(n_366),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_407),
.B(n_403),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_494),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_L g576 ( 
.A(n_470),
.B(n_295),
.C(n_311),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_500),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_403),
.B(n_253),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_457),
.B(n_254),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_446),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_440),
.B(n_257),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_505),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_442),
.B(n_281),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_450),
.A2(n_354),
.B1(n_352),
.B2(n_317),
.Y(n_586)
);

O2A1O1Ixp33_ASAP7_75t_L g587 ( 
.A1(n_468),
.A2(n_231),
.B(n_246),
.C(n_262),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_459),
.B(n_293),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_437),
.Y(n_589)
);

BUFx5_ASAP7_75t_L g590 ( 
.A(n_452),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_437),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_305),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_488),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_460),
.B(n_307),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_439),
.A2(n_352),
.B1(n_354),
.B2(n_309),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_502),
.A2(n_207),
.B(n_220),
.C(n_308),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_411),
.B(n_447),
.Y(n_597)
);

AND2x6_ASAP7_75t_SL g598 ( 
.A(n_410),
.B(n_298),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_447),
.B(n_317),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_490),
.A2(n_313),
.B1(n_393),
.B2(n_389),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_458),
.B(n_389),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_467),
.B(n_23),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_469),
.B(n_393),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_466),
.B(n_453),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_454),
.B(n_455),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_412),
.B(n_26),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_R g607 ( 
.A(n_476),
.B(n_69),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_524),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_601),
.A2(n_511),
.B(n_428),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_524),
.A2(n_470),
.B1(n_483),
.B2(n_484),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_569),
.A2(n_435),
.B1(n_479),
.B2(n_511),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_526),
.B(n_483),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_601),
.A2(n_511),
.B(n_471),
.Y(n_613)
);

BUFx2_ASAP7_75t_SL g614 ( 
.A(n_565),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_465),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_552),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_516),
.B(n_472),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_552),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_516),
.B(n_487),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_566),
.A2(n_597),
.B(n_538),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_529),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_573),
.A2(n_491),
.B(n_504),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_518),
.B(n_491),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_526),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_552),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_536),
.B(n_27),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_552),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_591),
.A2(n_512),
.B1(n_509),
.B2(n_507),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_517),
.A2(n_509),
.B1(n_507),
.B2(n_506),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_549),
.B(n_27),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_528),
.B(n_405),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_567),
.B(n_29),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_600),
.B(n_496),
.C(n_495),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_562),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_540),
.B(n_30),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_554),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_549),
.B(n_30),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_540),
.A2(n_519),
.B(n_539),
.C(n_543),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_585),
.B(n_519),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_544),
.B(n_34),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_559),
.B(n_533),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_591),
.A2(n_464),
.B1(n_463),
.B2(n_461),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_526),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_563),
.B(n_36),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_562),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_607),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_563),
.B(n_36),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_542),
.A2(n_416),
.B1(n_449),
.B2(n_441),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_576),
.B(n_441),
.C(n_438),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_562),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_560),
.B(n_37),
.Y(n_652)
);

AO21x2_ASAP7_75t_L g653 ( 
.A1(n_599),
.A2(n_433),
.B(n_431),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_589),
.A2(n_576),
.B1(n_571),
.B2(n_580),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_522),
.B(n_39),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_546),
.B(n_40),
.Y(n_657)
);

BUFx12f_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_598),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_606),
.B(n_42),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_553),
.A2(n_415),
.B1(n_413),
.B2(n_408),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_575),
.B(n_602),
.Y(n_662)
);

NOR2x1_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_406),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_557),
.A2(n_384),
.B(n_379),
.C(n_374),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_557),
.B(n_43),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_534),
.A2(n_379),
.B1(n_45),
.B2(n_48),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_R g668 ( 
.A(n_515),
.B(n_44),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_556),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_581),
.B(n_115),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_545),
.A2(n_118),
.B(n_172),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_570),
.B(n_49),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_604),
.A2(n_568),
.B(n_550),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_574),
.B(n_50),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_551),
.A2(n_114),
.B(n_170),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_523),
.B(n_50),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_595),
.B(n_51),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_577),
.B(n_583),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_537),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_555),
.A2(n_123),
.B(n_169),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_594),
.B(n_52),
.Y(n_683)
);

O2A1O1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_587),
.A2(n_548),
.B(n_596),
.C(n_582),
.Y(n_684)
);

BUFx4f_ASAP7_75t_L g685 ( 
.A(n_558),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_588),
.A2(n_128),
.B(n_167),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_558),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_564),
.A2(n_110),
.B(n_165),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_579),
.A2(n_104),
.B(n_164),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_545),
.B(n_54),
.C(n_55),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_541),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_521),
.B(n_59),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_520),
.A2(n_73),
.B(n_78),
.C(n_79),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_527),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_561),
.A2(n_81),
.B(n_85),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_547),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_584),
.A2(n_95),
.B(n_100),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_592),
.A2(n_131),
.B(n_134),
.C(n_135),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_530),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_531),
.A2(n_151),
.B(n_142),
.C(n_143),
.Y(n_700)
);

OAI22x1_ASAP7_75t_L g701 ( 
.A1(n_643),
.A2(n_605),
.B1(n_144),
.B2(n_146),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_639),
.A2(n_561),
.B1(n_572),
.B2(n_605),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_SL g703 ( 
.A1(n_610),
.A2(n_586),
.B(n_590),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_624),
.B(n_590),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_614),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_662),
.B(n_621),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_626),
.B(n_657),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_668),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_665),
.A2(n_644),
.B(n_648),
.C(n_656),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_634),
.B(n_646),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_654),
.B(n_680),
.Y(n_711)
);

AO31x2_ASAP7_75t_L g712 ( 
.A1(n_664),
.A2(n_698),
.A3(n_649),
.B(n_688),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_640),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_692),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_666),
.B(n_681),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_611),
.B(n_678),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_677),
.A2(n_686),
.A3(n_682),
.B(n_689),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_630),
.B(n_637),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_658),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_615),
.A2(n_617),
.B1(n_660),
.B2(n_623),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_622),
.A2(n_650),
.B(n_619),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_612),
.B(n_647),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_663),
.B(n_652),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_694),
.B(n_699),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_SL g726 ( 
.A(n_616),
.B(n_618),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_696),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_674),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_679),
.B(n_655),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_690),
.A2(n_691),
.B1(n_676),
.B2(n_667),
.Y(n_730)
);

CKINVDCx8_ASAP7_75t_R g731 ( 
.A(n_659),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_631),
.A2(n_629),
.B(n_642),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_685),
.B(n_683),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_685),
.B(n_670),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_687),
.B(n_636),
.Y(n_735)
);

AO31x2_ASAP7_75t_L g736 ( 
.A1(n_697),
.A2(n_653),
.A3(n_671),
.B(n_700),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_645),
.A2(n_628),
.B(n_627),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_671),
.A2(n_693),
.A3(n_627),
.B(n_625),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_661),
.A2(n_620),
.B(n_633),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_669),
.B(n_593),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_658),
.Y(n_741)
);

AO31x2_ASAP7_75t_L g742 ( 
.A1(n_609),
.A2(n_601),
.A3(n_603),
.B(n_613),
.Y(n_742)
);

OAI21x1_ASAP7_75t_SL g743 ( 
.A1(n_695),
.A2(n_672),
.B(n_673),
.Y(n_743)
);

OAI22x1_ASAP7_75t_L g744 ( 
.A1(n_643),
.A2(n_439),
.B1(n_529),
.B2(n_484),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_608),
.B(n_593),
.Y(n_745)
);

AO31x2_ASAP7_75t_L g746 ( 
.A1(n_609),
.A2(n_601),
.A3(n_603),
.B(n_613),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_608),
.B(n_593),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_684),
.A2(n_638),
.B(n_675),
.C(n_620),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_608),
.B(n_593),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_658),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_639),
.A2(n_477),
.B1(n_632),
.B2(n_635),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_673),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_608),
.B(n_593),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_608),
.B(n_524),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_679),
.A2(n_626),
.B1(n_611),
.B2(n_630),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_608),
.B(n_524),
.Y(n_756)
);

OAI21x1_ASAP7_75t_SL g757 ( 
.A1(n_695),
.A2(n_672),
.B(n_673),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_SL g758 ( 
.A(n_610),
.B(n_401),
.C(n_476),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_651),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_673),
.Y(n_760)
);

NOR4xp25_ASAP7_75t_L g761 ( 
.A(n_684),
.B(n_596),
.C(n_638),
.D(n_691),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_658),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_SL g763 ( 
.A(n_610),
.B(n_401),
.C(n_476),
.Y(n_763)
);

AO31x2_ASAP7_75t_L g764 ( 
.A1(n_609),
.A2(n_601),
.A3(n_603),
.B(n_613),
.Y(n_764)
);

AOI21xp33_ASAP7_75t_L g765 ( 
.A1(n_611),
.A2(n_524),
.B(n_401),
.Y(n_765)
);

AO31x2_ASAP7_75t_L g766 ( 
.A1(n_609),
.A2(n_601),
.A3(n_603),
.B(n_613),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_608),
.B(n_593),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_593),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_R g769 ( 
.A(n_659),
.B(n_532),
.Y(n_769)
);

AOI21xp33_ASAP7_75t_L g770 ( 
.A1(n_611),
.A2(n_524),
.B(n_401),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_608),
.B(n_524),
.Y(n_771)
);

AO31x2_ASAP7_75t_L g772 ( 
.A1(n_609),
.A2(n_601),
.A3(n_603),
.B(n_613),
.Y(n_772)
);

AO31x2_ASAP7_75t_L g773 ( 
.A1(n_609),
.A2(n_601),
.A3(n_603),
.B(n_613),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_684),
.A2(n_638),
.B(n_675),
.C(n_620),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_608),
.B(n_524),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_608),
.B(n_593),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_684),
.A2(n_638),
.B(n_675),
.C(n_620),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_611),
.B(n_524),
.C(n_401),
.Y(n_778)
);

NAND3x1_ASAP7_75t_L g779 ( 
.A(n_610),
.B(n_439),
.C(n_484),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_608),
.B(n_593),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_634),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_709),
.A2(n_751),
.B(n_748),
.C(n_777),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_745),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

BUFx2_ASAP7_75t_R g785 ( 
.A(n_731),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_714),
.B(n_716),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_749),
.Y(n_787)
);

OAI21x1_ASAP7_75t_SL g788 ( 
.A1(n_743),
.A2(n_757),
.B(n_721),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_755),
.A2(n_707),
.B1(n_711),
.B2(n_717),
.Y(n_789)
);

NOR2x1_ASAP7_75t_R g790 ( 
.A(n_741),
.B(n_750),
.Y(n_790)
);

OAI221xp5_ASAP7_75t_L g791 ( 
.A1(n_755),
.A2(n_729),
.B1(n_776),
.B2(n_768),
.C(n_780),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_739),
.A2(n_722),
.B(n_761),
.Y(n_792)
);

BUFx12f_ASAP7_75t_L g793 ( 
.A(n_762),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_761),
.B(n_713),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_753),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_715),
.B(n_728),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_720),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_740),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_779),
.A2(n_778),
.B1(n_758),
.B2(n_763),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_767),
.Y(n_800)
);

NAND2x1p5_ASAP7_75t_L g801 ( 
.A(n_705),
.B(n_752),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_765),
.B(n_770),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_744),
.A2(n_706),
.B1(n_719),
.B2(n_733),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_735),
.A2(n_756),
.B1(n_754),
.B2(n_771),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_710),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_703),
.A2(n_775),
.B(n_724),
.C(n_702),
.Y(n_806)
);

INVx8_ASAP7_75t_L g807 ( 
.A(n_781),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_708),
.A2(n_734),
.B1(n_704),
.B2(n_725),
.Y(n_808)
);

AO21x2_ASAP7_75t_L g809 ( 
.A1(n_732),
.A2(n_703),
.B(n_737),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_723),
.A2(n_701),
.B1(n_727),
.B2(n_730),
.Y(n_810)
);

BUFx12f_ASAP7_75t_L g811 ( 
.A(n_769),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_760),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_742),
.Y(n_813)
);

AO21x2_ASAP7_75t_L g814 ( 
.A1(n_738),
.A2(n_746),
.B(n_772),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_773),
.A2(n_766),
.A3(n_764),
.B(n_746),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_746),
.B(n_773),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_764),
.B(n_773),
.Y(n_817)
);

INVx11_ASAP7_75t_L g818 ( 
.A(n_726),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_766),
.B(n_738),
.Y(n_819)
);

AO31x2_ASAP7_75t_L g820 ( 
.A1(n_712),
.A2(n_774),
.A3(n_777),
.B(n_748),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_736),
.A2(n_758),
.B1(n_763),
.B2(n_717),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_718),
.A2(n_774),
.B(n_748),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_714),
.B(n_716),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_741),
.Y(n_824)
);

OAI21x1_ASAP7_75t_SL g825 ( 
.A1(n_743),
.A2(n_695),
.B(n_757),
.Y(n_825)
);

NAND2x1p5_ASAP7_75t_L g826 ( 
.A(n_759),
.B(n_651),
.Y(n_826)
);

CKINVDCx11_ASAP7_75t_R g827 ( 
.A(n_731),
.Y(n_827)
);

AO21x2_ASAP7_75t_L g828 ( 
.A1(n_743),
.A2(n_757),
.B(n_739),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_758),
.A2(n_763),
.B1(n_717),
.B2(n_778),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_759),
.B(n_651),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_758),
.A2(n_763),
.B1(n_778),
.B2(n_526),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_755),
.A2(n_721),
.B1(n_714),
.B2(n_751),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_759),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_748),
.A2(n_777),
.B(n_774),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_720),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_794),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_823),
.B(n_786),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_813),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_794),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_832),
.B(n_789),
.Y(n_840)
);

HB1xp67_ASAP7_75t_SL g841 ( 
.A(n_785),
.Y(n_841)
);

BUFx4f_ASAP7_75t_L g842 ( 
.A(n_807),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_827),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_832),
.B(n_789),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_791),
.A2(n_803),
.B1(n_829),
.B2(n_802),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_798),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_788),
.B(n_825),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_793),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_818),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_782),
.A2(n_791),
.B(n_834),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_829),
.A2(n_831),
.B1(n_799),
.B2(n_783),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_816),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_824),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_817),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_782),
.B(n_792),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_815),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_815),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_797),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_785),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_784),
.Y(n_860)
);

NOR2x1p5_ASAP7_75t_L g861 ( 
.A(n_811),
.B(n_796),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_819),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_SL g863 ( 
.A1(n_807),
.A2(n_800),
.B1(n_787),
.B2(n_795),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_807),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_792),
.B(n_806),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_821),
.A2(n_810),
.B1(n_804),
.B2(n_805),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_812),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_814),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_867),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_852),
.B(n_856),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_853),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_SL g872 ( 
.A1(n_863),
.A2(n_821),
.B(n_801),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_837),
.B(n_808),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_847),
.B(n_822),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_846),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_840),
.B(n_834),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_846),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_856),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_838),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_857),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_836),
.B(n_820),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_854),
.B(n_820),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_836),
.B(n_828),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_839),
.B(n_828),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_839),
.B(n_809),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_840),
.B(n_844),
.Y(n_886)
);

BUFx4f_ASAP7_75t_SL g887 ( 
.A(n_853),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_872),
.B(n_863),
.C(n_860),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_879),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_887),
.B(n_835),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_870),
.B(n_862),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_886),
.B(n_844),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_870),
.B(n_862),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_878),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_870),
.B(n_868),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_875),
.B(n_855),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_886),
.B(n_855),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_876),
.B(n_865),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_875),
.B(n_865),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_877),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_882),
.B(n_868),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_880),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_876),
.B(n_850),
.Y(n_903)
);

NAND2x1p5_ASAP7_75t_SL g904 ( 
.A(n_885),
.B(n_849),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_901),
.B(n_885),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_892),
.B(n_869),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_901),
.B(n_885),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_898),
.B(n_883),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_895),
.B(n_883),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_894),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_899),
.B(n_896),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_899),
.B(n_877),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_896),
.B(n_881),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_891),
.B(n_884),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_902),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_907),
.B(n_905),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_911),
.B(n_893),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_907),
.B(n_893),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_911),
.B(n_900),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_912),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_912),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_906),
.B(n_897),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_910),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_913),
.B(n_889),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_913),
.B(n_904),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_910),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_907),
.B(n_874),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_915),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_906),
.B(n_903),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_908),
.B(n_903),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_915),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_929),
.B(n_905),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_916),
.B(n_909),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_919),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_923),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_930),
.B(n_914),
.Y(n_936)
);

NAND4xp25_ASAP7_75t_L g937 ( 
.A(n_922),
.B(n_888),
.C(n_845),
.D(n_851),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_919),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_924),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_916),
.B(n_909),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_924),
.Y(n_941)
);

NAND4xp25_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_888),
.C(n_866),
.D(n_873),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_926),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_928),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_931),
.Y(n_945)
);

NOR2x1p5_ASAP7_75t_L g946 ( 
.A(n_917),
.B(n_871),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_935),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_933),
.B(n_927),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_938),
.B(n_871),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_942),
.A2(n_920),
.B1(n_921),
.B2(n_927),
.C(n_918),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_935),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_943),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_949),
.B(n_871),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_950),
.A2(n_934),
.B(n_937),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_L g955 ( 
.A1(n_947),
.A2(n_941),
.B(n_939),
.C(n_944),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_948),
.B(n_887),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_948),
.A2(n_946),
.B1(n_951),
.B2(n_932),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_952),
.A2(n_933),
.B1(n_940),
.B2(n_936),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_952),
.A2(n_890),
.B(n_842),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_955),
.Y(n_960)
);

BUFx24_ASAP7_75t_SL g961 ( 
.A(n_957),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_SL g962 ( 
.A(n_956),
.B(n_853),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_954),
.B(n_940),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_L g964 ( 
.A1(n_958),
.A2(n_945),
.B1(n_944),
.B2(n_943),
.C(n_873),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_953),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_960),
.B(n_959),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_965),
.Y(n_967)
);

NOR2x1p5_ASAP7_75t_L g968 ( 
.A(n_963),
.B(n_843),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_962),
.B(n_853),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_961),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_967),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_790),
.C(n_848),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_966),
.B(n_945),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_970),
.B(n_964),
.C(n_859),
.Y(n_974)
);

NOR2x1_ASAP7_75t_L g975 ( 
.A(n_968),
.B(n_858),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_971),
.A2(n_969),
.B(n_861),
.Y(n_976)
);

NOR2x1_ASAP7_75t_L g977 ( 
.A(n_975),
.B(n_864),
.Y(n_977)
);

XNOR2x1_ASAP7_75t_L g978 ( 
.A(n_977),
.B(n_973),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_976),
.Y(n_979)
);

OAI22x1_ASAP7_75t_L g980 ( 
.A1(n_979),
.A2(n_972),
.B1(n_978),
.B2(n_861),
.Y(n_980)
);

XNOR2xp5_ASAP7_75t_L g981 ( 
.A(n_978),
.B(n_841),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_981),
.A2(n_830),
.B(n_826),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_982),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_982),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_SL g985 ( 
.A1(n_984),
.A2(n_980),
.B1(n_842),
.B2(n_974),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_985),
.A2(n_983),
.B(n_842),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_986),
.B(n_833),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_987),
.A2(n_849),
.B1(n_864),
.B2(n_842),
.Y(n_988)
);


endmodule