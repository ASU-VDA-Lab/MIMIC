module real_jpeg_31241_n_21 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_121, n_11, n_14, n_7, n_18, n_3, n_119, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_120, n_21);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_119;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;
input n_120;

output n_21;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_15),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_1),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_17),
.C(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_97),
.Y(n_96)
);

NAND2x1p5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_4),
.A2(n_15),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_4),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_7),
.A2(n_61),
.B(n_119),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.C(n_121),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_8),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_9),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_9),
.B(n_105),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_10),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_20),
.B(n_71),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_20),
.C(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_12),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_89),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_14),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_19),
.Y(n_102)
);

HAxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.CON(n_21),
.SN(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_29),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_25),
.A2(n_42),
.B(n_44),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_25),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_41),
.B(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI31xp33_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_38),
.A3(n_39),
.B(n_111),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_43),
.C(n_45),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_104),
.B(n_110),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_95),
.B(n_103),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_88),
.B(n_94),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_78),
.B(n_84),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_70),
.B(n_74),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_59),
.B(n_68),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_58),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_58),
.C(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_66),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.C(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_120),
.Y(n_65)
);


endmodule