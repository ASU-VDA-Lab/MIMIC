module fake_jpeg_9360_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_36),
.B1(n_28),
.B2(n_16),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_25),
.B1(n_36),
.B2(n_38),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_17),
.B(n_23),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_20),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_66),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_46),
.B1(n_22),
.B2(n_20),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_78),
.B1(n_81),
.B2(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_69),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_35),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_65),
.B(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_24),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_79),
.B1(n_62),
.B2(n_64),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_34),
.C(n_39),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_54),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_0),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_26),
.B(n_31),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_39),
.B1(n_42),
.B2(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_34),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_100),
.B(n_101),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_44),
.B1(n_80),
.B2(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_42),
.B(n_33),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_75),
.B1(n_74),
.B2(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_71),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_110),
.C(n_112),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_119),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_114),
.B1(n_117),
.B2(n_122),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_80),
.Y(n_110)
);

XNOR2x2_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_80),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_44),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_89),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_54),
.B1(n_51),
.B2(n_8),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_8),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_85),
.B(n_86),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_51),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_1),
.C(n_5),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_102),
.B1(n_100),
.B2(n_88),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_122),
.B1(n_117),
.B2(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_103),
.B1(n_91),
.B2(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_122),
.B1(n_112),
.B2(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_94),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_94),
.B(n_2),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_141),
.B1(n_135),
.B2(n_125),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_108),
.B(n_122),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_144),
.B(n_136),
.Y(n_153)
);

AOI321xp33_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_15),
.A3(n_7),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_99),
.B(n_2),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_128),
.C(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_142),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_147),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_137),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_127),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_149),
.C(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_157),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_155),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_126),
.B1(n_123),
.B2(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_156),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_123),
.B1(n_129),
.B2(n_125),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_125),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_164),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_156),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_138),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_7),
.B(n_14),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_6),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_170),
.B(n_152),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_155),
.B(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_173),
.C(n_174),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_162),
.B1(n_143),
.B2(n_168),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_173),
.B1(n_15),
.B2(n_6),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);


endmodule